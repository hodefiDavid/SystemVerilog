    Mac OS X            	   2  �     
                                      ATTR      
  �   v                 �     )user.drive.can_manage_team_drive_members   �     user.drive.email   �   !  user.drive.id      �      user.drive.md5     �     user.drive.mime_type        $user.drive.shortcut.target.stableid         user.drive.stableid            user.drive.team_drive_id 1medina.dorit@gmail.com1HreDOCQ7BA2TPnOP0NoSvWXdgf-2nDQc3279e52d537970fc58cf2bdc5d4caa31application/octet-stream067496