    Mac OS X            	   2  �     
                                      ATTR      
  �   v                 �     )user.drive.can_manage_team_drive_members   �     user.drive.email   �   !  user.drive.id      �      user.drive.md5     �     user.drive.mime_type        $user.drive.shortcut.target.stableid         user.drive.stableid            user.drive.team_drive_id 1medina.dorit@gmail.com1IXbgibdQaFmQJMkjvqPPRe0D66uVX0Iib183fbbaeb028670f7896d8668753237application/octet-stream067500