package fpu_txn_pkg;

  import uvm_pkg::*;

  `include "uvm_macros.svh";

  `include "fpu_sv_utils.svh";
  `include "fp_operand.svh";
  `include "fp_transaction.svh";
  `include "fpu_request.svh";
  `include "fpu_response.svh";

endpackage // fpu_txn_pkg

