    Mac OS X            	   2  �     
                                      ATTR      
  �   v                 �     )user.drive.can_manage_team_drive_members   �     user.drive.email   �   !  user.drive.id      �      user.drive.md5     �     user.drive.mime_type        $user.drive.shortcut.target.stableid         user.drive.stableid            user.drive.team_drive_id 1medina.dorit@gmail.com1IJZ1gz0_aQ3Joiyau5HQWVAbWTmfmk_Wd346bce8c7131d4dceeb1c2da52722b6application/octet-stream067501