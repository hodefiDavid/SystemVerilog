    Mac OS X            	   2  �     
                                      ATTR      
  �   v                 �     )user.drive.can_manage_team_drive_members   �     user.drive.email   �   !  user.drive.id      �      user.drive.md5     �     user.drive.mime_type        $user.drive.shortcut.target.stableid         user.drive.stableid            user.drive.team_drive_id 1medina.dorit@gmail.com1Ilkd6QOgUZCQtZyELQlgR55MaEVRjjj33062abfa3683e64ae7f9fc53e3b8d5aaapplication/octet-stream067503