
module pre_norm_addsub_DW01_cmp2_8_1 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [7:0] A;
  input [7:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43;

  inv01 U6 ( .Y(n15), .A(n26) );
  inv01 U7 ( .Y(n32), .A(n16) );
  nor02 U8 ( .Y(n17), .A0(B[4]), .A1(n34) );
  nor02 U9 ( .Y(n18), .A0(B[3]), .A1(n35) );
  inv01 U10 ( .Y(n19), .A(n36) );
  nor02 U11 ( .Y(n16), .A0(n19), .A1(n20) );
  nor02 U12 ( .Y(n21), .A0(n17), .A1(n18) );
  inv01 U13 ( .Y(n20), .A(n21) );
  inv02 U14 ( .Y(n35), .A(A[3]) );
  inv02 U15 ( .Y(n34), .A(A[4]) );
  nand02 U16 ( .Y(n39), .A0(n42), .A1(n22) );
  inv01 U17 ( .Y(n23), .A(n37) );
  inv01 U18 ( .Y(n24), .A(B[2]) );
  inv01 U19 ( .Y(n25), .A(n41) );
  inv01 U20 ( .Y(n26), .A(n40) );
  nand02 U21 ( .Y(n27), .A0(n23), .A1(n24) );
  nand02 U22 ( .Y(n28), .A0(n25), .A1(n26) );
  nand02 U23 ( .Y(n29), .A0(n27), .A1(n28) );
  inv01 U24 ( .Y(n22), .A(n29) );
  inv01 U25 ( .Y(n38), .A(n39) );
  inv02 U26 ( .Y(n41), .A(A[1]) );
  inv02 U27 ( .Y(n37), .A(A[2]) );
  or02 U28 ( .Y(n30), .A0(n31), .A1(B[5]) );
  nand02 U29 ( .Y(n31), .A0(n32), .A1(n33) );
  inv04 U30 ( .Y(n43), .A(B[0]) );
  or03 U31 ( .Y(LT_LE), .A0(B[7]), .A1(B[6]), .A2(n30) );
  nand02 U32 ( .Y(n33), .A0(B[4]), .A1(n34) );
  ao221 U33 ( .Y(n36), .A0(n37), .A1(B[2]), .B0(n35), .B1(B[3]), .C0(n38) );
  ao21 U34 ( .Y(n42), .A0(n15), .A1(n41), .B0(B[1]) );
  nor02 U35 ( .Y(n40), .A0(n43), .A1(A[0]) );
endmodule


module pre_norm_addsub_DW01_sub_8_0 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   carry_7_, carry_6_, carry_5_, carry_4_, carry_3_, carry_2_, carry_1_,
         n165, n6, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164;
  wire   [7:0] B_not;

  buf02 U6 ( .Y(DIFF[7]), .A(n165) );
  inv02 U7 ( .Y(B_not[7]), .A(B[7]) );
  xor2 U8 ( .Y(n6), .A0(B_not[0]), .A1(A[0]) );
  inv01 U9 ( .Y(DIFF[0]), .A(n6) );
  or02 U10 ( .Y(n8), .A0(B_not[0]), .A1(A[0]) );
  inv02 U11 ( .Y(B_not[0]), .A(B[0]) );
  inv01 U12 ( .Y(DIFF[6]), .A(n9) );
  inv02 U13 ( .Y(carry_7_), .A(n10) );
  inv02 U14 ( .Y(n11), .A(B_not[6]) );
  inv02 U15 ( .Y(n12), .A(A[6]) );
  inv02 U16 ( .Y(n13), .A(carry_6_) );
  nor02 U17 ( .Y(n14), .A0(n11), .A1(n15) );
  nor02 U18 ( .Y(n16), .A0(n12), .A1(n17) );
  nor02 U19 ( .Y(n18), .A0(n13), .A1(n19) );
  nor02 U20 ( .Y(n20), .A0(n13), .A1(n21) );
  nor02 U21 ( .Y(n9), .A0(n22), .A1(n23) );
  nor02 U22 ( .Y(n24), .A0(n12), .A1(n13) );
  nor02 U23 ( .Y(n25), .A0(n11), .A1(n13) );
  nor02 U24 ( .Y(n26), .A0(n11), .A1(n12) );
  nor02 U25 ( .Y(n10), .A0(n26), .A1(n27) );
  nor02 U26 ( .Y(n28), .A0(A[6]), .A1(carry_6_) );
  inv01 U27 ( .Y(n15), .A(n28) );
  nor02 U28 ( .Y(n29), .A0(B_not[6]), .A1(carry_6_) );
  inv01 U29 ( .Y(n17), .A(n29) );
  nor02 U30 ( .Y(n30), .A0(B_not[6]), .A1(A[6]) );
  inv01 U31 ( .Y(n19), .A(n30) );
  nor02 U32 ( .Y(n31), .A0(n11), .A1(n12) );
  inv01 U33 ( .Y(n21), .A(n31) );
  nor02 U34 ( .Y(n32), .A0(n14), .A1(n16) );
  inv01 U35 ( .Y(n22), .A(n32) );
  nor02 U36 ( .Y(n33), .A0(n18), .A1(n20) );
  inv01 U37 ( .Y(n23), .A(n33) );
  nor02 U38 ( .Y(n34), .A0(n24), .A1(n25) );
  inv01 U39 ( .Y(n27), .A(n34) );
  inv02 U40 ( .Y(B_not[6]), .A(B[6]) );
  inv01 U41 ( .Y(DIFF[5]), .A(n35) );
  inv02 U42 ( .Y(carry_6_), .A(n36) );
  inv02 U43 ( .Y(n37), .A(B_not[5]) );
  inv02 U44 ( .Y(n38), .A(A[5]) );
  inv02 U45 ( .Y(n39), .A(carry_5_) );
  nor02 U46 ( .Y(n40), .A0(n37), .A1(n41) );
  nor02 U47 ( .Y(n42), .A0(n38), .A1(n43) );
  nor02 U48 ( .Y(n44), .A0(n39), .A1(n45) );
  nor02 U49 ( .Y(n46), .A0(n39), .A1(n47) );
  nor02 U50 ( .Y(n35), .A0(n48), .A1(n49) );
  nor02 U51 ( .Y(n50), .A0(n38), .A1(n39) );
  nor02 U52 ( .Y(n51), .A0(n37), .A1(n39) );
  nor02 U53 ( .Y(n52), .A0(n37), .A1(n38) );
  nor02 U54 ( .Y(n36), .A0(n52), .A1(n53) );
  nor02 U55 ( .Y(n54), .A0(A[5]), .A1(carry_5_) );
  inv01 U56 ( .Y(n41), .A(n54) );
  nor02 U57 ( .Y(n55), .A0(B_not[5]), .A1(carry_5_) );
  inv01 U58 ( .Y(n43), .A(n55) );
  nor02 U59 ( .Y(n56), .A0(B_not[5]), .A1(A[5]) );
  inv01 U60 ( .Y(n45), .A(n56) );
  nor02 U61 ( .Y(n57), .A0(n37), .A1(n38) );
  inv01 U62 ( .Y(n47), .A(n57) );
  nor02 U63 ( .Y(n58), .A0(n40), .A1(n42) );
  inv01 U64 ( .Y(n48), .A(n58) );
  nor02 U65 ( .Y(n59), .A0(n44), .A1(n46) );
  inv01 U66 ( .Y(n49), .A(n59) );
  nor02 U67 ( .Y(n60), .A0(n50), .A1(n51) );
  inv01 U68 ( .Y(n53), .A(n60) );
  inv02 U69 ( .Y(B_not[5]), .A(B[5]) );
  inv01 U70 ( .Y(DIFF[4]), .A(n61) );
  inv02 U71 ( .Y(carry_5_), .A(n62) );
  inv02 U72 ( .Y(n63), .A(B_not[4]) );
  inv02 U73 ( .Y(n64), .A(A[4]) );
  inv02 U74 ( .Y(n65), .A(carry_4_) );
  nor02 U75 ( .Y(n66), .A0(n63), .A1(n67) );
  nor02 U76 ( .Y(n68), .A0(n64), .A1(n69) );
  nor02 U77 ( .Y(n70), .A0(n65), .A1(n71) );
  nor02 U78 ( .Y(n72), .A0(n65), .A1(n73) );
  nor02 U79 ( .Y(n61), .A0(n74), .A1(n75) );
  nor02 U80 ( .Y(n76), .A0(n64), .A1(n65) );
  nor02 U81 ( .Y(n77), .A0(n63), .A1(n65) );
  nor02 U82 ( .Y(n78), .A0(n63), .A1(n64) );
  nor02 U83 ( .Y(n62), .A0(n78), .A1(n79) );
  nor02 U84 ( .Y(n80), .A0(A[4]), .A1(carry_4_) );
  inv01 U85 ( .Y(n67), .A(n80) );
  nor02 U86 ( .Y(n81), .A0(B_not[4]), .A1(carry_4_) );
  inv01 U87 ( .Y(n69), .A(n81) );
  nor02 U88 ( .Y(n82), .A0(B_not[4]), .A1(A[4]) );
  inv01 U89 ( .Y(n71), .A(n82) );
  nor02 U90 ( .Y(n83), .A0(n63), .A1(n64) );
  inv01 U91 ( .Y(n73), .A(n83) );
  nor02 U92 ( .Y(n84), .A0(n66), .A1(n68) );
  inv01 U93 ( .Y(n74), .A(n84) );
  nor02 U94 ( .Y(n85), .A0(n70), .A1(n72) );
  inv01 U95 ( .Y(n75), .A(n85) );
  nor02 U96 ( .Y(n86), .A0(n76), .A1(n77) );
  inv01 U97 ( .Y(n79), .A(n86) );
  inv02 U98 ( .Y(B_not[4]), .A(B[4]) );
  inv01 U99 ( .Y(DIFF[3]), .A(n87) );
  inv02 U100 ( .Y(carry_4_), .A(n88) );
  inv02 U101 ( .Y(n89), .A(B_not[3]) );
  inv02 U102 ( .Y(n90), .A(A[3]) );
  inv02 U103 ( .Y(n91), .A(carry_3_) );
  nor02 U104 ( .Y(n92), .A0(n89), .A1(n93) );
  nor02 U105 ( .Y(n94), .A0(n90), .A1(n95) );
  nor02 U106 ( .Y(n96), .A0(n91), .A1(n97) );
  nor02 U107 ( .Y(n98), .A0(n91), .A1(n99) );
  nor02 U108 ( .Y(n87), .A0(n100), .A1(n101) );
  nor02 U109 ( .Y(n102), .A0(n90), .A1(n91) );
  nor02 U110 ( .Y(n103), .A0(n89), .A1(n91) );
  nor02 U111 ( .Y(n104), .A0(n89), .A1(n90) );
  nor02 U112 ( .Y(n88), .A0(n104), .A1(n105) );
  nor02 U113 ( .Y(n106), .A0(A[3]), .A1(carry_3_) );
  inv01 U114 ( .Y(n93), .A(n106) );
  nor02 U115 ( .Y(n107), .A0(B_not[3]), .A1(carry_3_) );
  inv01 U116 ( .Y(n95), .A(n107) );
  nor02 U117 ( .Y(n108), .A0(B_not[3]), .A1(A[3]) );
  inv01 U118 ( .Y(n97), .A(n108) );
  nor02 U119 ( .Y(n109), .A0(n89), .A1(n90) );
  inv01 U120 ( .Y(n99), .A(n109) );
  nor02 U121 ( .Y(n110), .A0(n92), .A1(n94) );
  inv01 U122 ( .Y(n100), .A(n110) );
  nor02 U123 ( .Y(n111), .A0(n96), .A1(n98) );
  inv01 U124 ( .Y(n101), .A(n111) );
  nor02 U125 ( .Y(n112), .A0(n102), .A1(n103) );
  inv01 U126 ( .Y(n105), .A(n112) );
  inv02 U127 ( .Y(B_not[3]), .A(B[3]) );
  inv01 U128 ( .Y(DIFF[2]), .A(n113) );
  inv02 U129 ( .Y(carry_3_), .A(n114) );
  inv02 U130 ( .Y(n115), .A(B_not[2]) );
  inv02 U131 ( .Y(n116), .A(A[2]) );
  inv02 U132 ( .Y(n117), .A(carry_2_) );
  nor02 U133 ( .Y(n118), .A0(n115), .A1(n119) );
  nor02 U134 ( .Y(n120), .A0(n116), .A1(n121) );
  nor02 U135 ( .Y(n122), .A0(n117), .A1(n123) );
  nor02 U136 ( .Y(n124), .A0(n117), .A1(n125) );
  nor02 U137 ( .Y(n113), .A0(n126), .A1(n127) );
  nor02 U138 ( .Y(n128), .A0(n116), .A1(n117) );
  nor02 U139 ( .Y(n129), .A0(n115), .A1(n117) );
  nor02 U140 ( .Y(n130), .A0(n115), .A1(n116) );
  nor02 U141 ( .Y(n114), .A0(n130), .A1(n131) );
  nor02 U142 ( .Y(n132), .A0(A[2]), .A1(carry_2_) );
  inv01 U143 ( .Y(n119), .A(n132) );
  nor02 U144 ( .Y(n133), .A0(B_not[2]), .A1(carry_2_) );
  inv01 U145 ( .Y(n121), .A(n133) );
  nor02 U146 ( .Y(n134), .A0(B_not[2]), .A1(A[2]) );
  inv01 U147 ( .Y(n123), .A(n134) );
  nor02 U148 ( .Y(n135), .A0(n115), .A1(n116) );
  inv01 U149 ( .Y(n125), .A(n135) );
  nor02 U150 ( .Y(n136), .A0(n118), .A1(n120) );
  inv01 U151 ( .Y(n126), .A(n136) );
  nor02 U152 ( .Y(n137), .A0(n122), .A1(n124) );
  inv01 U153 ( .Y(n127), .A(n137) );
  nor02 U154 ( .Y(n138), .A0(n128), .A1(n129) );
  inv01 U155 ( .Y(n131), .A(n138) );
  inv02 U156 ( .Y(B_not[2]), .A(B[2]) );
  inv01 U157 ( .Y(DIFF[1]), .A(n139) );
  inv02 U158 ( .Y(carry_2_), .A(n140) );
  inv02 U159 ( .Y(n141), .A(B_not[1]) );
  inv02 U160 ( .Y(n142), .A(A[1]) );
  inv02 U161 ( .Y(n143), .A(carry_1_) );
  nor02 U162 ( .Y(n144), .A0(n141), .A1(n145) );
  nor02 U163 ( .Y(n146), .A0(n142), .A1(n147) );
  nor02 U164 ( .Y(n148), .A0(n143), .A1(n149) );
  nor02 U165 ( .Y(n150), .A0(n143), .A1(n151) );
  nor02 U166 ( .Y(n139), .A0(n152), .A1(n153) );
  nor02 U167 ( .Y(n154), .A0(n142), .A1(n143) );
  nor02 U168 ( .Y(n155), .A0(n141), .A1(n143) );
  nor02 U169 ( .Y(n156), .A0(n141), .A1(n142) );
  nor02 U170 ( .Y(n140), .A0(n156), .A1(n157) );
  nor02 U171 ( .Y(n158), .A0(A[1]), .A1(n8) );
  inv01 U172 ( .Y(n145), .A(n158) );
  nor02 U173 ( .Y(n159), .A0(B_not[1]), .A1(n8) );
  inv01 U174 ( .Y(n147), .A(n159) );
  nor02 U175 ( .Y(n160), .A0(B_not[1]), .A1(A[1]) );
  inv01 U176 ( .Y(n149), .A(n160) );
  nor02 U177 ( .Y(n161), .A0(n141), .A1(n142) );
  inv01 U178 ( .Y(n151), .A(n161) );
  nor02 U179 ( .Y(n162), .A0(n144), .A1(n146) );
  inv01 U180 ( .Y(n152), .A(n162) );
  nor02 U181 ( .Y(n163), .A0(n148), .A1(n150) );
  inv01 U182 ( .Y(n153), .A(n163) );
  nor02 U183 ( .Y(n164), .A0(n154), .A1(n155) );
  inv01 U184 ( .Y(n157), .A(n164) );
  inv02 U185 ( .Y(B_not[1]), .A(B[1]) );
  or02 U186 ( .Y(carry_1_), .A0(B_not[0]), .A1(A[0]) );
  fadd1 U2_7 ( .S(n165), .A(A[7]), .B(B_not[7]), .CI(carry_7_) );
endmodule


module pre_norm_addsub_DW01_inc_8_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;
  wire   carry_7_, carry_6_, carry_5_, carry_4_, carry_3_, carry_2_, n1;

  inv02 U5 ( .Y(n1), .A(SUM[0]) );
  inv02 U6 ( .Y(SUM[0]), .A(A[0]) );
  xor2 U7 ( .Y(SUM[7]), .A0(carry_7_), .A1(A[7]) );
  hadd1 U1_1_1 ( .S(SUM[1]), .CO(carry_2_), .A(A[1]), .B(n1) );
  hadd1 U1_1_2 ( .S(SUM[2]), .CO(carry_3_), .A(A[2]), .B(carry_2_) );
  hadd1 U1_1_3 ( .S(SUM[3]), .CO(carry_4_), .A(A[3]), .B(carry_3_) );
  hadd1 U1_1_4 ( .S(SUM[4]), .CO(carry_5_), .A(A[4]), .B(carry_4_) );
  hadd1 U1_1_5 ( .S(SUM[5]), .CO(carry_6_), .A(A[5]), .B(carry_5_) );
  hadd1 U1_1_6 ( .S(SUM[6]), .CO(carry_7_), .A(A[6]), .B(carry_6_) );
endmodule


module pre_norm_addsub_DW01_cmp2_8_0 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [7:0] A;
  input [7:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n85, n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84;

  inv16 U6 ( .Y(n15), .A(n62) );
  inv16 U7 ( .Y(LT_LE), .A(n15) );
  buf02 U8 ( .Y(n17), .A(A[4]) );
  inv01 U9 ( .Y(n18), .A(n17) );
  nand02 U10 ( .Y(n68), .A0(n19), .A1(n20) );
  inv01 U11 ( .Y(n21), .A(n71) );
  inv01 U12 ( .Y(n22), .A(n69) );
  inv01 U13 ( .Y(n23), .A(A[7]) );
  inv01 U14 ( .Y(n24), .A(n70) );
  nand02 U15 ( .Y(n25), .A0(n21), .A1(n22) );
  nand02 U16 ( .Y(n26), .A0(n21), .A1(n23) );
  nand02 U17 ( .Y(n27), .A0(n22), .A1(n24) );
  nand02 U18 ( .Y(n28), .A0(n23), .A1(n24) );
  nand02 U19 ( .Y(n29), .A0(n25), .A1(n26) );
  inv01 U20 ( .Y(n19), .A(n29) );
  nand02 U21 ( .Y(n30), .A0(n27), .A1(n28) );
  inv01 U22 ( .Y(n20), .A(n30) );
  inv01 U23 ( .Y(n69), .A(B[7]) );
  or02 U24 ( .Y(n31), .A0(n84), .A1(A[0]) );
  inv01 U25 ( .Y(n32), .A(n31) );
  nand02 U26 ( .Y(n70), .A0(n74), .A1(n33) );
  inv01 U27 ( .Y(n34), .A(n72) );
  inv01 U28 ( .Y(n35), .A(B[6]) );
  inv01 U29 ( .Y(n36), .A(n73) );
  inv01 U30 ( .Y(n37), .A(B[5]) );
  nand02 U31 ( .Y(n38), .A0(n34), .A1(n35) );
  nand02 U32 ( .Y(n39), .A0(n36), .A1(n37) );
  nand02 U33 ( .Y(n40), .A0(n38), .A1(n39) );
  inv01 U34 ( .Y(n33), .A(n40) );
  inv01 U35 ( .Y(n73), .A(A[5]) );
  inv01 U36 ( .Y(n72), .A(A[6]) );
  nand02 U37 ( .Y(n81), .A0(n83), .A1(n41) );
  inv01 U38 ( .Y(n42), .A(n79) );
  inv01 U39 ( .Y(n43), .A(B[2]) );
  inv01 U40 ( .Y(n44), .A(n82) );
  inv01 U41 ( .Y(n45), .A(n32) );
  nand02 U42 ( .Y(n46), .A0(n42), .A1(n43) );
  nand02 U43 ( .Y(n47), .A0(n44), .A1(n45) );
  nand02 U44 ( .Y(n48), .A0(n46), .A1(n47) );
  inv01 U45 ( .Y(n41), .A(n48) );
  inv01 U46 ( .Y(n80), .A(n81) );
  inv01 U47 ( .Y(n82), .A(A[1]) );
  inv01 U48 ( .Y(n79), .A(A[2]) );
  inv02 U49 ( .Y(n85), .A(n49) );
  inv01 U50 ( .Y(n50), .A(n67) );
  inv01 U51 ( .Y(n51), .A(B[7]) );
  nor02 U52 ( .Y(n52), .A0(n50), .A1(n51) );
  nor02 U53 ( .Y(n49), .A0(n52), .A1(n68) );
  inv04 U54 ( .Y(n65), .A(n85) );
  inv01 U55 ( .Y(n67), .A(A[7]) );
  inv01 U56 ( .Y(n84), .A(B[0]) );
  nand02 U57 ( .Y(n76), .A0(n78), .A1(n53) );
  inv01 U58 ( .Y(n54), .A(n18) );
  inv01 U59 ( .Y(n55), .A(B[4]) );
  inv01 U60 ( .Y(n56), .A(n77) );
  inv01 U61 ( .Y(n57), .A(B[3]) );
  nand02 U62 ( .Y(n58), .A0(n54), .A1(n55) );
  nand02 U63 ( .Y(n59), .A0(n56), .A1(n57) );
  nand02 U64 ( .Y(n60), .A0(n58), .A1(n59) );
  inv01 U65 ( .Y(n53), .A(n60) );
  inv01 U66 ( .Y(n75), .A(n76) );
  inv01 U67 ( .Y(n77), .A(A[3]) );
  inv16 U68 ( .Y(n61), .A(n64) );
  inv16 U69 ( .Y(n62), .A(n61) );
  inv16 U70 ( .Y(n63), .A(n66) );
  inv16 U71 ( .Y(n64), .A(n63) );
  inv16 U72 ( .Y(n66), .A(n65) );
  nand02 U73 ( .Y(n71), .A0(B[6]), .A1(n72) );
  ao221 U74 ( .Y(n74), .A0(n18), .A1(B[4]), .B0(n73), .B1(B[5]), .C0(n75) );
  ao221 U75 ( .Y(n78), .A0(n79), .A1(B[2]), .B0(n77), .B1(B[3]), .C0(n80) );
  ao21 U76 ( .Y(n83), .A0(n32), .A1(n82), .B0(B[1]) );
endmodule


module pre_norm_addsub ( clk_i, opa_i, opb_i, fracta_28_o, fractb_28_o, exp_o
 );
  input [31:0] opa_i;
  input [31:0] opb_i;
  output [27:0] fracta_28_o;
  output [27:0] fractb_28_o;
  output [7:0] exp_o;
  input clk_i;
  wire   s_fracta_28_o_26_, s_fracta_28_o_25_, s_fracta_28_o_24_,
         s_fracta_28_o_23_, s_fracta_28_o_22_, s_fracta_28_o_21_,
         s_fracta_28_o_20_, s_fracta_28_o_19_, s_fracta_28_o_18_,
         s_fracta_28_o_17_, s_fracta_28_o_16_, s_fracta_28_o_15_,
         s_fracta_28_o_14_, s_fracta_28_o_13_, s_fracta_28_o_12_,
         s_fracta_28_o_11_, s_fracta_28_o_10_, s_fracta_28_o_9_,
         s_fracta_28_o_8_, s_fracta_28_o_7_, s_fracta_28_o_6_,
         s_fracta_28_o_5_, s_fracta_28_o_4_, s_fracta_28_o_3_,
         s_fractb_28_o_26_, s_fractb_28_o_25_, s_fractb_28_o_24_,
         s_fractb_28_o_23_, s_fractb_28_o_22_, s_fractb_28_o_21_,
         s_fractb_28_o_20_, s_fractb_28_o_19_, s_fractb_28_o_18_,
         s_fractb_28_o_17_, s_fractb_28_o_16_, s_fractb_28_o_15_,
         s_fractb_28_o_14_, s_fractb_28_o_13_, s_fractb_28_o_12_,
         s_fractb_28_o_11_, s_fractb_28_o_10_, s_fractb_28_o_9_,
         s_fractb_28_o_8_, s_fractb_28_o_7_, s_fractb_28_o_6_,
         s_fractb_28_o_5_, s_fractb_28_o_4_, s_fractb_28_o_3_, n5488, n5489,
         n____return128, s_exp_o389_7_, s_exp_o389_6_, s_exp_o389_5_,
         s_exp_o389_4_, s_exp_o389_3_, s_exp_o389_2_, s_exp_o389_1_,
         s_exp_o389_0_, s_exp_diff436_7_, s_exp_diff436_6_, s_exp_diff436_5_,
         s_exp_diff436_4_, s_exp_diff436_3_, s_exp_diff436_2_,
         s_exp_diff436_1_, s_exp_diff436_0_, s_exp_diff_7_, s_exp_diff_6_,
         s_exp_diff_5_, s_exp_diff_4_, s_exp_diff_3_, s_exp_diff_2_,
         s_exp_diff_1_, s_exp_diff_0_, n____return498_7_, n____return498_6_,
         n____return498_5_, n____return498_4_, n____return498_3_,
         n____return498_2_, n____return498_1_, n____return498_0_, s_rzeros_4_,
         s_rzeros_3_, s_rzeros_2_, s_rzeros_1_, s_rzeros_0_, n____return2686,
         U403_U6_Z_7, U403_U6_Z_6, U403_U6_Z_5, U403_U6_Z_4, U403_U6_Z_3,
         U403_U6_Z_2, U403_U6_Z_1, U403_U6_Z_0, U403_U5_Z_7, U403_U5_Z_6,
         U403_U5_Z_5, U403_U5_Z_4, U403_U5_Z_3, U403_U5_Z_2, U403_U5_Z_1,
         U403_U5_Z_0, U403_U4_Z_7, U403_U4_Z_6, U403_U4_Z_5, U403_U4_Z_4,
         U403_U4_Z_3, U403_U4_Z_2, U403_U4_Z_1, U403_U4_Z_0, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487;
  wire   [7:0] s_exp_o;

  dff fracta_28_o_reg_27_ ( .Q(fracta_28_o[27]), .D(1'b0), .CLK(clk_i) );
  dff fractb_28_o_reg_27_ ( .Q(fractb_28_o[27]), .D(1'b0), .CLK(clk_i) );
  dff exp_o_reg_7_ ( .Q(exp_o[7]), .D(s_exp_o[7]), .CLK(clk_i) );
  dff exp_o_reg_6_ ( .Q(exp_o[6]), .D(s_exp_o[6]), .CLK(clk_i) );
  dff exp_o_reg_5_ ( .Q(exp_o[5]), .D(s_exp_o[5]), .CLK(clk_i) );
  dff exp_o_reg_4_ ( .Q(n5488), .D(s_exp_o[4]), .CLK(clk_i) );
  dff exp_o_reg_3_ ( .Q(exp_o[3]), .D(s_exp_o[3]), .CLK(clk_i) );
  dff exp_o_reg_2_ ( .Q(exp_o[2]), .D(s_exp_o[2]), .CLK(clk_i) );
  dff exp_o_reg_1_ ( .Q(exp_o[1]), .D(s_exp_o[1]), .CLK(clk_i) );
  dff exp_o_reg_0_ ( .Q(n5489), .D(s_exp_o[0]), .CLK(clk_i) );
  dff fracta_28_o_reg_26_ ( .Q(fracta_28_o[26]), .D(s_fracta_28_o_26_), .CLK(
        clk_i) );
  dff fracta_28_o_reg_25_ ( .Q(fracta_28_o[25]), .D(s_fracta_28_o_25_), .CLK(
        clk_i) );
  dff fracta_28_o_reg_24_ ( .Q(fracta_28_o[24]), .D(s_fracta_28_o_24_), .CLK(
        clk_i) );
  dff fracta_28_o_reg_23_ ( .Q(fracta_28_o[23]), .D(s_fracta_28_o_23_), .CLK(
        clk_i) );
  dff fracta_28_o_reg_22_ ( .Q(fracta_28_o[22]), .D(s_fracta_28_o_22_), .CLK(
        clk_i) );
  dff fracta_28_o_reg_21_ ( .Q(fracta_28_o[21]), .D(s_fracta_28_o_21_), .CLK(
        clk_i) );
  dff fracta_28_o_reg_20_ ( .Q(fracta_28_o[20]), .D(s_fracta_28_o_20_), .CLK(
        clk_i) );
  dff fracta_28_o_reg_19_ ( .Q(fracta_28_o[19]), .D(s_fracta_28_o_19_), .CLK(
        clk_i) );
  dff fracta_28_o_reg_18_ ( .Q(fracta_28_o[18]), .D(s_fracta_28_o_18_), .CLK(
        clk_i) );
  dff fracta_28_o_reg_17_ ( .Q(fracta_28_o[17]), .D(s_fracta_28_o_17_), .CLK(
        clk_i) );
  dff fracta_28_o_reg_16_ ( .Q(fracta_28_o[16]), .D(s_fracta_28_o_16_), .CLK(
        clk_i) );
  dff fracta_28_o_reg_15_ ( .Q(fracta_28_o[15]), .D(s_fracta_28_o_15_), .CLK(
        clk_i) );
  dff fracta_28_o_reg_14_ ( .Q(fracta_28_o[14]), .D(s_fracta_28_o_14_), .CLK(
        clk_i) );
  dff fracta_28_o_reg_13_ ( .Q(fracta_28_o[13]), .D(s_fracta_28_o_13_), .CLK(
        clk_i) );
  dff fracta_28_o_reg_12_ ( .Q(fracta_28_o[12]), .D(s_fracta_28_o_12_), .CLK(
        clk_i) );
  dff fracta_28_o_reg_11_ ( .Q(fracta_28_o[11]), .D(s_fracta_28_o_11_), .CLK(
        clk_i) );
  dff fracta_28_o_reg_10_ ( .Q(fracta_28_o[10]), .D(s_fracta_28_o_10_), .CLK(
        clk_i) );
  dff fracta_28_o_reg_9_ ( .Q(fracta_28_o[9]), .D(s_fracta_28_o_9_), .CLK(
        clk_i) );
  dff fracta_28_o_reg_8_ ( .Q(fracta_28_o[8]), .D(s_fracta_28_o_8_), .CLK(
        clk_i) );
  dff fracta_28_o_reg_7_ ( .Q(fracta_28_o[7]), .D(s_fracta_28_o_7_), .CLK(
        clk_i) );
  dff fracta_28_o_reg_6_ ( .Q(fracta_28_o[6]), .D(s_fracta_28_o_6_), .CLK(
        clk_i) );
  dff fracta_28_o_reg_5_ ( .Q(fracta_28_o[5]), .D(s_fracta_28_o_5_), .CLK(
        clk_i) );
  dff fracta_28_o_reg_4_ ( .Q(fracta_28_o[4]), .D(s_fracta_28_o_4_), .CLK(
        clk_i) );
  dff fracta_28_o_reg_3_ ( .Q(fracta_28_o[3]), .D(s_fracta_28_o_3_), .CLK(
        clk_i) );
  dff fracta_28_o_reg_2_ ( .Q(fracta_28_o[2]), .D(n3413), .CLK(clk_i) );
  dff fracta_28_o_reg_1_ ( .Q(fracta_28_o[1]), .D(n3417), .CLK(clk_i) );
  dff fracta_28_o_reg_0_ ( .Q(fracta_28_o[0]), .D(n3415), .CLK(clk_i) );
  dff fractb_28_o_reg_26_ ( .Q(fractb_28_o[26]), .D(s_fractb_28_o_26_), .CLK(
        clk_i) );
  dff fractb_28_o_reg_25_ ( .Q(fractb_28_o[25]), .D(s_fractb_28_o_25_), .CLK(
        clk_i) );
  dff fractb_28_o_reg_24_ ( .Q(fractb_28_o[24]), .D(s_fractb_28_o_24_), .CLK(
        clk_i) );
  dff fractb_28_o_reg_23_ ( .Q(fractb_28_o[23]), .D(s_fractb_28_o_23_), .CLK(
        clk_i) );
  dff fractb_28_o_reg_22_ ( .Q(fractb_28_o[22]), .D(s_fractb_28_o_22_), .CLK(
        clk_i) );
  dff fractb_28_o_reg_21_ ( .Q(fractb_28_o[21]), .D(s_fractb_28_o_21_), .CLK(
        clk_i) );
  dff fractb_28_o_reg_20_ ( .Q(fractb_28_o[20]), .D(s_fractb_28_o_20_), .CLK(
        clk_i) );
  dff fractb_28_o_reg_19_ ( .Q(fractb_28_o[19]), .D(s_fractb_28_o_19_), .CLK(
        clk_i) );
  dff fractb_28_o_reg_18_ ( .Q(fractb_28_o[18]), .D(s_fractb_28_o_18_), .CLK(
        clk_i) );
  dff fractb_28_o_reg_17_ ( .Q(fractb_28_o[17]), .D(s_fractb_28_o_17_), .CLK(
        clk_i) );
  dff fractb_28_o_reg_16_ ( .Q(fractb_28_o[16]), .D(s_fractb_28_o_16_), .CLK(
        clk_i) );
  dff fractb_28_o_reg_15_ ( .Q(fractb_28_o[15]), .D(s_fractb_28_o_15_), .CLK(
        clk_i) );
  dff fractb_28_o_reg_14_ ( .Q(fractb_28_o[14]), .D(s_fractb_28_o_14_), .CLK(
        clk_i) );
  dff fractb_28_o_reg_13_ ( .Q(fractb_28_o[13]), .D(s_fractb_28_o_13_), .CLK(
        clk_i) );
  dff fractb_28_o_reg_12_ ( .Q(fractb_28_o[12]), .D(s_fractb_28_o_12_), .CLK(
        clk_i) );
  dff fractb_28_o_reg_11_ ( .Q(fractb_28_o[11]), .D(s_fractb_28_o_11_), .CLK(
        clk_i) );
  dff fractb_28_o_reg_10_ ( .Q(fractb_28_o[10]), .D(s_fractb_28_o_10_), .CLK(
        clk_i) );
  dff fractb_28_o_reg_9_ ( .Q(fractb_28_o[9]), .D(s_fractb_28_o_9_), .CLK(
        clk_i) );
  dff fractb_28_o_reg_8_ ( .Q(fractb_28_o[8]), .D(s_fractb_28_o_8_), .CLK(
        clk_i) );
  dff fractb_28_o_reg_7_ ( .Q(fractb_28_o[7]), .D(s_fractb_28_o_7_), .CLK(
        clk_i) );
  dff fractb_28_o_reg_6_ ( .Q(fractb_28_o[6]), .D(s_fractb_28_o_6_), .CLK(
        clk_i) );
  dff fractb_28_o_reg_5_ ( .Q(fractb_28_o[5]), .D(s_fractb_28_o_5_), .CLK(
        clk_i) );
  dff fractb_28_o_reg_4_ ( .Q(fractb_28_o[4]), .D(s_fractb_28_o_4_), .CLK(
        clk_i) );
  dff fractb_28_o_reg_3_ ( .Q(fractb_28_o[3]), .D(s_fractb_28_o_3_), .CLK(
        clk_i) );
  dff fractb_28_o_reg_2_ ( .Q(fractb_28_o[2]), .D(n3402), .CLK(clk_i) );
  dff fractb_28_o_reg_1_ ( .Q(fractb_28_o[1]), .D(n3400), .CLK(clk_i) );
  dff fractb_28_o_reg_0_ ( .Q(fractb_28_o[0]), .D(n3398), .CLK(clk_i) );
  dff s_exp_o_reg_7_ ( .Q(s_exp_o[7]), .D(s_exp_o389_7_), .CLK(clk_i) );
  dff s_exp_o_reg_6_ ( .Q(s_exp_o[6]), .D(s_exp_o389_6_), .CLK(clk_i) );
  dff s_exp_o_reg_5_ ( .Q(s_exp_o[5]), .D(s_exp_o389_5_), .CLK(clk_i) );
  dff s_exp_o_reg_4_ ( .Q(s_exp_o[4]), .D(s_exp_o389_4_), .CLK(clk_i) );
  dff s_exp_o_reg_3_ ( .Q(s_exp_o[3]), .D(s_exp_o389_3_), .CLK(clk_i) );
  dff s_exp_o_reg_2_ ( .Q(s_exp_o[2]), .D(s_exp_o389_2_), .CLK(clk_i) );
  dff s_exp_o_reg_1_ ( .Q(s_exp_o[1]), .D(s_exp_o389_1_), .CLK(clk_i) );
  dff s_exp_o_reg_0_ ( .Q(s_exp_o[0]), .D(s_exp_o389_0_), .CLK(clk_i) );
  dff s_exp_diff_reg_7_ ( .Q(s_exp_diff_7_), .QB(n5487), .D(s_exp_diff436_7_), 
        .CLK(clk_i) );
  dff s_exp_diff_reg_6_ ( .Q(s_exp_diff_6_), .QB(n5486), .D(s_exp_diff436_6_), 
        .CLK(clk_i) );
  dff s_exp_diff_reg_5_ ( .Q(s_exp_diff_5_), .QB(n5485), .D(s_exp_diff436_5_), 
        .CLK(clk_i) );
  dff s_exp_diff_reg_4_ ( .Q(s_exp_diff_4_), .D(s_exp_diff436_4_), .CLK(clk_i)
         );
  dff s_exp_diff_reg_3_ ( .Q(s_exp_diff_3_), .D(s_exp_diff436_3_), .CLK(clk_i)
         );
  dff s_exp_diff_reg_2_ ( .Q(s_exp_diff_2_), .D(s_exp_diff436_2_), .CLK(clk_i)
         );
  dff s_exp_diff_reg_1_ ( .Q(s_exp_diff_1_), .D(s_exp_diff436_1_), .CLK(clk_i)
         );
  dff s_exp_diff_reg_0_ ( .Q(s_exp_diff_0_), .D(s_exp_diff436_0_), .CLK(clk_i)
         );
  inv08 U978 ( .Y(n3327), .A(n4006) );
  inv02 U979 ( .Y(n4006), .A(n____return128) );
  ao22 U980 ( .Y(n3328), .A0(n5418), .A1(n5283), .B0(n5419), .B1(n5309) );
  inv01 U981 ( .Y(n3329), .A(n3328) );
  ao22 U982 ( .Y(n3330), .A0(n5418), .A1(n5286), .B0(n5419), .B1(n5311) );
  inv01 U983 ( .Y(n3331), .A(n3330) );
  ao22 U984 ( .Y(n3332), .A0(n5418), .A1(n5306), .B0(n5419), .B1(n5294) );
  inv01 U985 ( .Y(n3333), .A(n3332) );
  ao22 U986 ( .Y(n3334), .A0(n5418), .A1(n5292), .B0(n5419), .B1(n5312) );
  inv01 U987 ( .Y(n3335), .A(n3334) );
  ao22 U988 ( .Y(n3336), .A0(n5418), .A1(n5311), .B0(n5419), .B1(n5292) );
  inv01 U989 ( .Y(n3337), .A(n3336) );
  nand02 U990 ( .Y(n5459), .A0(n3338), .A1(n3339) );
  inv01 U991 ( .Y(n3340), .A(n5305) );
  inv01 U992 ( .Y(n3341), .A(n5294) );
  inv01 U993 ( .Y(n3342), .A(n5418) );
  inv01 U994 ( .Y(n3343), .A(n5419) );
  nand02 U995 ( .Y(n3344), .A0(n3340), .A1(n3341) );
  nand02 U996 ( .Y(n3345), .A0(n3340), .A1(n3342) );
  nand02 U997 ( .Y(n3346), .A0(n3341), .A1(n3343) );
  nand02 U998 ( .Y(n3347), .A0(n3342), .A1(n3343) );
  nand02 U999 ( .Y(n3348), .A0(n3344), .A1(n3345) );
  inv01 U1000 ( .Y(n3338), .A(n3348) );
  nand02 U1001 ( .Y(n3349), .A0(n3346), .A1(n3347) );
  inv01 U1002 ( .Y(n3339), .A(n3349) );
  ao22 U1003 ( .Y(n3350), .A0(n5418), .A1(n5305), .B0(n5419), .B1(n5286) );
  inv01 U1004 ( .Y(n3351), .A(n3350) );
  ao22 U1005 ( .Y(n3352), .A0(n5418), .A1(n5295), .B0(n5419), .B1(n5303) );
  inv01 U1006 ( .Y(n3353), .A(n3352) );
  ao22 U1007 ( .Y(n3354), .A0(n5418), .A1(n5307), .B0(n5419), .B1(n5288) );
  inv01 U1008 ( .Y(n3355), .A(n3354) );
  nand02 U1009 ( .Y(n5455), .A0(n3356), .A1(n3357) );
  inv01 U1010 ( .Y(n3358), .A(n5299) );
  inv01 U1011 ( .Y(n3359), .A(n5303) );
  inv01 U1012 ( .Y(n3360), .A(n5418) );
  inv01 U1013 ( .Y(n3361), .A(n5419) );
  nand02 U1014 ( .Y(n3362), .A0(n3358), .A1(n3359) );
  nand02 U1015 ( .Y(n3363), .A0(n3358), .A1(n3360) );
  nand02 U1016 ( .Y(n3364), .A0(n3359), .A1(n3361) );
  nand02 U1017 ( .Y(n3365), .A0(n3360), .A1(n3361) );
  nand02 U1018 ( .Y(n3366), .A0(n3362), .A1(n3363) );
  inv01 U1019 ( .Y(n3356), .A(n3366) );
  nand02 U1020 ( .Y(n3367), .A0(n3364), .A1(n3365) );
  inv01 U1021 ( .Y(n3357), .A(n3367) );
  ao22 U1022 ( .Y(n3368), .A0(n5418), .A1(n5299), .B0(n5419), .B1(n5313) );
  inv01 U1023 ( .Y(n3369), .A(n3368) );
  ao22 U1024 ( .Y(n3370), .A0(n5418), .A1(n5315), .B0(n5419), .B1(n5297) );
  inv01 U1025 ( .Y(n3371), .A(n3370) );
  ao22 U1026 ( .Y(n3372), .A0(n5418), .A1(n5308), .B0(n5419), .B1(n5287) );
  inv01 U1027 ( .Y(n3373), .A(n3372) );
  ao22 U1028 ( .Y(n3374), .A0(n5418), .A1(n5313), .B0(n5419), .B1(n5290) );
  inv01 U1029 ( .Y(n3375), .A(n3374) );
  ao22 U1030 ( .Y(n3376), .A0(n5418), .A1(n5309), .B0(n5419), .B1(n5296) );
  inv01 U1031 ( .Y(n3377), .A(n3376) );
  ao22 U1032 ( .Y(n3378), .A0(n5418), .A1(n5287), .B0(n5419), .B1(n5315) );
  inv01 U1033 ( .Y(n3379), .A(n3378) );
  ao22 U1034 ( .Y(n3380), .A0(n5418), .A1(n5290), .B0(n5419), .B1(n5307) );
  inv01 U1035 ( .Y(n3381), .A(n3380) );
  ao22 U1036 ( .Y(n3382), .A0(n5418), .A1(n5296), .B0(n5419), .B1(n5308) );
  inv01 U1037 ( .Y(n3383), .A(n3382) );
  buf02 U1038 ( .Y(n3384), .A(n5477) );
  buf02 U1039 ( .Y(n3385), .A(n5474) );
  buf02 U1040 ( .Y(n3386), .A(n5479) );
  buf02 U1041 ( .Y(n3387), .A(n5476) );
  buf02 U1042 ( .Y(n3388), .A(n5471) );
  buf02 U1043 ( .Y(n3389), .A(n5478) );
  buf02 U1044 ( .Y(n3390), .A(n5475) );
  ao22 U1045 ( .Y(n3391), .A0(n5418), .A1(n5462), .B0(n5419), .B1(n5306) );
  inv01 U1046 ( .Y(n3392), .A(n3391) );
  ao22 U1047 ( .Y(n3393), .A0(n5418), .A1(n5278), .B0(n5419), .B1(n5283) );
  inv01 U1048 ( .Y(n3394), .A(n3393) );
  or02 U1049 ( .Y(n3395), .A0(n5268), .A1(n5278) );
  inv01 U1050 ( .Y(n3396), .A(n3395) );
  or02 U1051 ( .Y(n3397), .A0(n5360), .A1(n5222) );
  inv01 U1052 ( .Y(n3398), .A(n3397) );
  or02 U1053 ( .Y(n3399), .A0(n5344), .A1(n5223) );
  inv01 U1054 ( .Y(n3400), .A(n3399) );
  or02 U1055 ( .Y(n3401), .A0(n5328), .A1(n5222) );
  inv01 U1056 ( .Y(n3402), .A(n3401) );
  ao22 U1057 ( .Y(n3403), .A0(n5418), .A1(n5314), .B0(n5419), .B1(n5295) );
  inv01 U1058 ( .Y(n3404), .A(n3403) );
  ao22 U1059 ( .Y(n3405), .A0(n5432), .A1(n5433), .B0(n5434), .B1(
        s_exp_diff_2_) );
  inv01 U1060 ( .Y(n3406), .A(n3405) );
  and02 U1061 ( .Y(n3408), .A0(n5212), .A1(n5197) );
  and02 U1062 ( .Y(n3407), .A0(n5212), .A1(n5197) );
  inv01 U1063 ( .Y(n5480), .A(n3409) );
  nor02 U1064 ( .Y(n3410), .A0(n4957), .A1(n5207) );
  nor02 U1065 ( .Y(n3411), .A0(n5469), .A1(n5206) );
  nor02 U1066 ( .Y(n3409), .A0(n3410), .A1(n3411) );
  inv02 U1067 ( .Y(n5232), .A(n5277) );
  or02 U1068 ( .Y(n3412), .A0(n____return128), .A1(n5328) );
  inv01 U1069 ( .Y(n3413), .A(n3412) );
  or02 U1070 ( .Y(n3414), .A0(n____return128), .A1(n5360) );
  inv01 U1071 ( .Y(n3415), .A(n3414) );
  or02 U1072 ( .Y(n3416), .A0(n____return128), .A1(n5344) );
  inv01 U1073 ( .Y(n3417), .A(n3416) );
  ao21 U1074 ( .Y(n3418), .A0(n5284), .A1(n5314), .B0(n3424) );
  inv01 U1075 ( .Y(n3419), .A(n3418) );
  inv01 U1076 ( .Y(n5440), .A(n3420) );
  nor02 U1077 ( .Y(n3421), .A0(n5180), .A1(n5219) );
  nor02 U1078 ( .Y(n3422), .A0(n5284), .A1(n4929) );
  nor02 U1079 ( .Y(n3420), .A0(n3421), .A1(n3422) );
  buf02 U1080 ( .Y(n4929), .A(n5424) );
  buf04 U1081 ( .Y(exp_o[0]), .A(n5489) );
  nand03 U1082 ( .Y(n3423), .A0(n3943), .A1(n5315), .A2(n5194) );
  inv02 U1083 ( .Y(n3424), .A(n3423) );
  inv02 U1084 ( .Y(n5433), .A(s_exp_diff_2_) );
  inv01 U1085 ( .Y(s_fracta_28_o_25_), .A(n3425) );
  nor02 U1086 ( .Y(n3426), .A0(n5333), .A1(n4861) );
  nor02 U1087 ( .Y(n3427), .A0(n5222), .A1(n5427) );
  nor02 U1088 ( .Y(n3425), .A0(n3426), .A1(n3427) );
  inv01 U1089 ( .Y(s_fracta_28_o_23_), .A(n3428) );
  nor02 U1090 ( .Y(n3429), .A0(n5337), .A1(n4861) );
  nor02 U1091 ( .Y(n3430), .A0(n5222), .A1(n5429) );
  nor02 U1092 ( .Y(n3428), .A0(n3429), .A1(n3430) );
  inv01 U1093 ( .Y(s_fracta_28_o_21_), .A(n3431) );
  nor02 U1094 ( .Y(n3432), .A0(n4860), .A1(n5202) );
  nor02 U1095 ( .Y(n3433), .A0(n5223), .A1(n5435) );
  nor02 U1096 ( .Y(n3431), .A0(n3432), .A1(n3433) );
  inv01 U1097 ( .Y(s_fracta_28_o_24_), .A(n3434) );
  nor02 U1098 ( .Y(n3435), .A0(n5335), .A1(n5426) );
  nor02 U1099 ( .Y(n3436), .A0(n5222), .A1(n5428) );
  nor02 U1100 ( .Y(n3434), .A0(n3435), .A1(n3436) );
  inv01 U1101 ( .Y(s_fracta_28_o_18_), .A(n3437) );
  nor02 U1102 ( .Y(n3438), .A0(n5347), .A1(n5202) );
  nor02 U1103 ( .Y(n3439), .A0(n5223), .A1(n5442) );
  nor02 U1104 ( .Y(n3437), .A0(n3438), .A1(n3439) );
  inv01 U1105 ( .Y(s_fracta_28_o_22_), .A(n3440) );
  nor02 U1106 ( .Y(n3441), .A0(n5340), .A1(n5203) );
  nor02 U1107 ( .Y(n3442), .A0(n5222), .A1(n5430) );
  nor02 U1108 ( .Y(n3440), .A0(n3441), .A1(n3442) );
  inv01 U1109 ( .Y(s_fracta_28_o_19_), .A(n3443) );
  nor02 U1110 ( .Y(n3444), .A0(n4878), .A1(n5203) );
  nor02 U1111 ( .Y(n3445), .A0(n5223), .A1(n5441) );
  nor02 U1112 ( .Y(n3443), .A0(n3444), .A1(n3445) );
  inv01 U1113 ( .Y(s_fracta_28_o_17_), .A(n3446) );
  nor02 U1114 ( .Y(n3447), .A0(n5349), .A1(n5203) );
  nor02 U1115 ( .Y(n3448), .A0(n5222), .A1(n5443) );
  nor02 U1116 ( .Y(n3446), .A0(n3447), .A1(n3448) );
  inv01 U1117 ( .Y(s_fracta_28_o_20_), .A(n3449) );
  nor02 U1118 ( .Y(n3450), .A0(n4863), .A1(n5202) );
  nor02 U1119 ( .Y(n3451), .A0(n5223), .A1(n5436) );
  nor02 U1120 ( .Y(n3449), .A0(n3450), .A1(n3451) );
  inv01 U1121 ( .Y(s_fracta_28_o_16_), .A(n3452) );
  nor02 U1122 ( .Y(n3453), .A0(n5351), .A1(n5202) );
  nor02 U1123 ( .Y(n3454), .A0(n5222), .A1(n5444) );
  nor02 U1124 ( .Y(n3452), .A0(n3453), .A1(n3454) );
  inv01 U1125 ( .Y(s_fracta_28_o_26_), .A(n3455) );
  nor02 U1126 ( .Y(n3456), .A0(n5041), .A1(n5426) );
  nor02 U1127 ( .Y(n3457), .A0(n5425), .A1(n5222) );
  nor02 U1128 ( .Y(n3455), .A0(n3456), .A1(n3457) );
  ao21 U1129 ( .Y(n3458), .A0(n5224), .A1(n5201), .B0(n5237) );
  inv01 U1130 ( .Y(n3459), .A(n3458) );
  or03 U1131 ( .Y(n3460), .A0(n5242), .A1(n5240), .A2(n5241) );
  inv01 U1132 ( .Y(n3461), .A(n3460) );
  inv04 U1133 ( .Y(exp_o[4]), .A(n4463) );
  nand03 U1134 ( .Y(n3462), .A0(n5199), .A1(n5288), .A2(n5289) );
  inv02 U1135 ( .Y(n3463), .A(n3462) );
  nand02 U1136 ( .Y(s_fracta_28_o_8_), .A0(n3464), .A1(n3465) );
  inv01 U1137 ( .Y(n3466), .A(n____return128) );
  inv01 U1138 ( .Y(n3467), .A(n5223) );
  inv01 U1139 ( .Y(n3468), .A(n5319) );
  inv01 U1140 ( .Y(n3469), .A(n5373) );
  nand02 U1141 ( .Y(n3470), .A0(n3466), .A1(n3467) );
  nand02 U1142 ( .Y(n3471), .A0(n3466), .A1(n3468) );
  nand02 U1143 ( .Y(n3472), .A0(n3467), .A1(n3469) );
  nand02 U1144 ( .Y(n3473), .A0(n3468), .A1(n3469) );
  nand02 U1145 ( .Y(n3474), .A0(n3470), .A1(n3471) );
  inv01 U1146 ( .Y(n3464), .A(n3474) );
  nand02 U1147 ( .Y(n3475), .A0(n3472), .A1(n3473) );
  inv01 U1148 ( .Y(n3465), .A(n3475) );
  nand02 U1149 ( .Y(s_fracta_28_o_12_), .A0(n3476), .A1(n3477) );
  inv01 U1150 ( .Y(n3478), .A(n3327) );
  inv01 U1151 ( .Y(n3479), .A(n5223) );
  inv01 U1152 ( .Y(n3480), .A(n4743) );
  inv01 U1153 ( .Y(n3481), .A(n5451) );
  nand02 U1154 ( .Y(n3482), .A0(n3478), .A1(n3479) );
  nand02 U1155 ( .Y(n3483), .A0(n3478), .A1(n3480) );
  nand02 U1156 ( .Y(n3484), .A0(n3479), .A1(n3481) );
  nand02 U1157 ( .Y(n3485), .A0(n3480), .A1(n3481) );
  nand02 U1158 ( .Y(n3486), .A0(n3482), .A1(n3483) );
  inv01 U1159 ( .Y(n3476), .A(n3486) );
  nand02 U1160 ( .Y(n3487), .A0(n3484), .A1(n3485) );
  inv01 U1161 ( .Y(n3477), .A(n3487) );
  nand02 U1162 ( .Y(s_fracta_28_o_7_), .A0(n3488), .A1(n3489) );
  inv01 U1163 ( .Y(n3490), .A(n3327) );
  inv01 U1164 ( .Y(n3491), .A(n5223) );
  inv01 U1165 ( .Y(n3492), .A(n4733) );
  inv01 U1166 ( .Y(n3493), .A(n5381) );
  nand02 U1167 ( .Y(n3494), .A0(n3490), .A1(n3491) );
  nand02 U1168 ( .Y(n3495), .A0(n3490), .A1(n3492) );
  nand02 U1169 ( .Y(n3496), .A0(n3491), .A1(n3493) );
  nand02 U1170 ( .Y(n3497), .A0(n3492), .A1(n3493) );
  nand02 U1171 ( .Y(n3498), .A0(n3494), .A1(n3495) );
  inv01 U1172 ( .Y(n3488), .A(n3498) );
  nand02 U1173 ( .Y(n3499), .A0(n3496), .A1(n3497) );
  inv01 U1174 ( .Y(n3489), .A(n3499) );
  nand02 U1175 ( .Y(s_exp_o389_3_), .A0(n3500), .A1(n3501) );
  inv01 U1176 ( .Y(n3502), .A(n3327) );
  inv01 U1177 ( .Y(n3503), .A(n5223) );
  inv01 U1178 ( .Y(n3504), .A(n4913) );
  inv01 U1179 ( .Y(n3505), .A(n4935) );
  nand02 U1180 ( .Y(n3506), .A0(n3502), .A1(n3503) );
  nand02 U1181 ( .Y(n3507), .A0(n3502), .A1(n3504) );
  nand02 U1182 ( .Y(n3508), .A0(n3503), .A1(n3505) );
  nand02 U1183 ( .Y(n3509), .A0(n3504), .A1(n3505) );
  nand02 U1184 ( .Y(n3510), .A0(n3506), .A1(n3507) );
  inv01 U1185 ( .Y(n3500), .A(n3510) );
  nand02 U1186 ( .Y(n3511), .A0(n3508), .A1(n3509) );
  inv01 U1187 ( .Y(n3501), .A(n3511) );
  nand02 U1188 ( .Y(s_fractb_28_o_8_), .A0(n3512), .A1(n3513) );
  inv01 U1189 ( .Y(n3514), .A(n3327) );
  inv01 U1190 ( .Y(n3515), .A(n5222) );
  inv01 U1191 ( .Y(n3516), .A(n5318) );
  inv01 U1192 ( .Y(n3517), .A(n5319) );
  nand02 U1193 ( .Y(n3518), .A0(n3514), .A1(n3515) );
  nand02 U1194 ( .Y(n3519), .A0(n3514), .A1(n3516) );
  nand02 U1195 ( .Y(n3520), .A0(n3515), .A1(n3517) );
  nand02 U1196 ( .Y(n3521), .A0(n3516), .A1(n3517) );
  nand02 U1197 ( .Y(n3522), .A0(n3518), .A1(n3519) );
  inv01 U1198 ( .Y(n3512), .A(n3522) );
  nand02 U1199 ( .Y(n3523), .A0(n3520), .A1(n3521) );
  inv01 U1200 ( .Y(n3513), .A(n3523) );
  nand02 U1201 ( .Y(s_fractb_28_o_10_), .A0(n3524), .A1(n3525) );
  inv01 U1202 ( .Y(n3526), .A(n____return128) );
  inv01 U1203 ( .Y(n3527), .A(n5222) );
  inv01 U1204 ( .Y(n3528), .A(n5359) );
  inv01 U1205 ( .Y(n3529), .A(n4735) );
  nand02 U1206 ( .Y(n3530), .A0(n3526), .A1(n3527) );
  nand02 U1207 ( .Y(n3531), .A0(n3526), .A1(n3528) );
  nand02 U1208 ( .Y(n3532), .A0(n3527), .A1(n3529) );
  nand02 U1209 ( .Y(n3533), .A0(n3528), .A1(n3529) );
  nand02 U1210 ( .Y(n3534), .A0(n3530), .A1(n3531) );
  inv01 U1211 ( .Y(n3524), .A(n3534) );
  nand02 U1212 ( .Y(n3535), .A0(n3532), .A1(n3533) );
  inv01 U1213 ( .Y(n3525), .A(n3535) );
  nand02 U1214 ( .Y(s_exp_o389_5_), .A0(n3536), .A1(n3537) );
  inv01 U1215 ( .Y(n3538), .A(n____return128) );
  inv01 U1216 ( .Y(n3539), .A(n5222) );
  inv01 U1217 ( .Y(n3540), .A(n4919) );
  inv01 U1218 ( .Y(n3541), .A(n4933) );
  nand02 U1219 ( .Y(n3542), .A0(n3538), .A1(n3539) );
  nand02 U1220 ( .Y(n3543), .A0(n3538), .A1(n3540) );
  nand02 U1221 ( .Y(n3544), .A0(n3539), .A1(n3541) );
  nand02 U1222 ( .Y(n3545), .A0(n3540), .A1(n3541) );
  nand02 U1223 ( .Y(n3546), .A0(n3542), .A1(n3543) );
  inv01 U1224 ( .Y(n3536), .A(n3546) );
  nand02 U1225 ( .Y(n3547), .A0(n3544), .A1(n3545) );
  inv01 U1226 ( .Y(n3537), .A(n3547) );
  nand02 U1227 ( .Y(s_fracta_28_o_9_), .A0(n3548), .A1(n3549) );
  inv01 U1228 ( .Y(n3550), .A(n____return128) );
  inv01 U1229 ( .Y(n3551), .A(n5222) );
  inv01 U1230 ( .Y(n3552), .A(n5317) );
  inv01 U1231 ( .Y(n3553), .A(n5361) );
  nand02 U1232 ( .Y(n3554), .A0(n3550), .A1(n3551) );
  nand02 U1233 ( .Y(n3555), .A0(n3550), .A1(n3552) );
  nand02 U1234 ( .Y(n3556), .A0(n3551), .A1(n3553) );
  nand02 U1235 ( .Y(n3557), .A0(n3552), .A1(n3553) );
  nand02 U1236 ( .Y(n3558), .A0(n3554), .A1(n3555) );
  inv01 U1237 ( .Y(n3548), .A(n3558) );
  nand02 U1238 ( .Y(n3559), .A0(n3556), .A1(n3557) );
  inv01 U1239 ( .Y(n3549), .A(n3559) );
  nand02 U1240 ( .Y(s_fracta_28_o_13_), .A0(n3560), .A1(n3561) );
  inv01 U1241 ( .Y(n3562), .A(n3327) );
  inv01 U1242 ( .Y(n3563), .A(n5223) );
  inv01 U1243 ( .Y(n3564), .A(n4739) );
  inv01 U1244 ( .Y(n3565), .A(n5448) );
  nand02 U1245 ( .Y(n3566), .A0(n3562), .A1(n3563) );
  nand02 U1246 ( .Y(n3567), .A0(n3562), .A1(n3564) );
  nand02 U1247 ( .Y(n3568), .A0(n3563), .A1(n3565) );
  nand02 U1248 ( .Y(n3569), .A0(n3564), .A1(n3565) );
  nand02 U1249 ( .Y(n3570), .A0(n3566), .A1(n3567) );
  inv01 U1250 ( .Y(n3560), .A(n3570) );
  nand02 U1251 ( .Y(n3571), .A0(n3568), .A1(n3569) );
  inv01 U1252 ( .Y(n3561), .A(n3571) );
  nand02 U1253 ( .Y(s_fractb_28_o_14_), .A0(n3572), .A1(n3573) );
  inv01 U1254 ( .Y(n3574), .A(n3327) );
  inv01 U1255 ( .Y(n3575), .A(n5223) );
  inv01 U1256 ( .Y(n3576), .A(n5354) );
  inv01 U1257 ( .Y(n3577), .A(n4737) );
  nand02 U1258 ( .Y(n3578), .A0(n3574), .A1(n3575) );
  nand02 U1259 ( .Y(n3579), .A0(n3574), .A1(n3576) );
  nand02 U1260 ( .Y(n3580), .A0(n3575), .A1(n3577) );
  nand02 U1261 ( .Y(n3581), .A0(n3576), .A1(n3577) );
  nand02 U1262 ( .Y(n3582), .A0(n3578), .A1(n3579) );
  inv01 U1263 ( .Y(n3572), .A(n3582) );
  nand02 U1264 ( .Y(n3583), .A0(n3580), .A1(n3581) );
  inv01 U1265 ( .Y(n3573), .A(n3583) );
  nand02 U1266 ( .Y(s_exp_o389_2_), .A0(n3584), .A1(n3585) );
  inv01 U1267 ( .Y(n3586), .A(n3327) );
  inv01 U1268 ( .Y(n3587), .A(n5223) );
  inv01 U1269 ( .Y(n3588), .A(n4922) );
  inv01 U1270 ( .Y(n3589), .A(n4939) );
  nand02 U1271 ( .Y(n3590), .A0(n3586), .A1(n3587) );
  nand02 U1272 ( .Y(n3591), .A0(n3586), .A1(n3588) );
  nand02 U1273 ( .Y(n3592), .A0(n3587), .A1(n3589) );
  nand02 U1274 ( .Y(n3593), .A0(n3588), .A1(n3589) );
  nand02 U1275 ( .Y(n3594), .A0(n3590), .A1(n3591) );
  inv01 U1276 ( .Y(n3584), .A(n3594) );
  nand02 U1277 ( .Y(n3595), .A0(n3592), .A1(n3593) );
  inv01 U1278 ( .Y(n3585), .A(n3595) );
  nand02 U1279 ( .Y(s_fracta_28_o_10_), .A0(n3596), .A1(n3597) );
  inv01 U1280 ( .Y(n3598), .A(n3327) );
  inv01 U1281 ( .Y(n3599), .A(n5223) );
  inv01 U1282 ( .Y(n3600), .A(n4735) );
  inv01 U1283 ( .Y(n3601), .A(n5456) );
  nand02 U1284 ( .Y(n3602), .A0(n3598), .A1(n3599) );
  nand02 U1285 ( .Y(n3603), .A0(n3598), .A1(n3600) );
  nand02 U1286 ( .Y(n3604), .A0(n3599), .A1(n3601) );
  nand02 U1287 ( .Y(n3605), .A0(n3600), .A1(n3601) );
  nand02 U1288 ( .Y(n3606), .A0(n3602), .A1(n3603) );
  inv01 U1289 ( .Y(n3596), .A(n3606) );
  nand02 U1290 ( .Y(n3607), .A0(n3604), .A1(n3605) );
  inv01 U1291 ( .Y(n3597), .A(n3607) );
  nand02 U1292 ( .Y(s_exp_o389_7_), .A0(n3608), .A1(n3609) );
  inv01 U1293 ( .Y(n3610), .A(n____return128) );
  inv01 U1294 ( .Y(n3611), .A(n5222) );
  inv01 U1295 ( .Y(n3612), .A(n4925) );
  inv01 U1296 ( .Y(n3613), .A(n4943) );
  nand02 U1297 ( .Y(n3614), .A0(n3610), .A1(n3611) );
  nand02 U1298 ( .Y(n3615), .A0(n3610), .A1(n3612) );
  nand02 U1299 ( .Y(n3616), .A0(n3611), .A1(n3613) );
  nand02 U1300 ( .Y(n3617), .A0(n3612), .A1(n3613) );
  nand02 U1301 ( .Y(n3618), .A0(n3614), .A1(n3615) );
  inv01 U1302 ( .Y(n3608), .A(n3618) );
  nand02 U1303 ( .Y(n3619), .A0(n3616), .A1(n3617) );
  inv01 U1304 ( .Y(n3609), .A(n3619) );
  nand02 U1305 ( .Y(s_exp_o389_4_), .A0(n3620), .A1(n3621) );
  inv01 U1306 ( .Y(n3622), .A(n3327) );
  inv01 U1307 ( .Y(n3623), .A(n5222) );
  inv01 U1308 ( .Y(n3624), .A(n4928) );
  inv01 U1309 ( .Y(n3625), .A(n4941) );
  nand02 U1310 ( .Y(n3626), .A0(n3622), .A1(n3623) );
  nand02 U1311 ( .Y(n3627), .A0(n3622), .A1(n3624) );
  nand02 U1312 ( .Y(n3628), .A0(n3623), .A1(n3625) );
  nand02 U1313 ( .Y(n3629), .A0(n3624), .A1(n3625) );
  nand02 U1314 ( .Y(n3630), .A0(n3626), .A1(n3627) );
  inv01 U1315 ( .Y(n3620), .A(n3630) );
  nand02 U1316 ( .Y(n3631), .A0(n3628), .A1(n3629) );
  inv01 U1317 ( .Y(n3621), .A(n3631) );
  nand02 U1318 ( .Y(s_fractb_28_o_5_), .A0(n3632), .A1(n3633) );
  inv01 U1319 ( .Y(n3634), .A(n3327) );
  inv01 U1320 ( .Y(n3635), .A(n5222) );
  inv01 U1321 ( .Y(n3636), .A(n5322) );
  inv01 U1322 ( .Y(n3637), .A(n5323) );
  nand02 U1323 ( .Y(n3638), .A0(n3634), .A1(n3635) );
  nand02 U1324 ( .Y(n3639), .A0(n3634), .A1(n3636) );
  nand02 U1325 ( .Y(n3640), .A0(n3635), .A1(n3637) );
  nand02 U1326 ( .Y(n3641), .A0(n3636), .A1(n3637) );
  nand02 U1327 ( .Y(n3642), .A0(n3638), .A1(n3639) );
  inv01 U1328 ( .Y(n3632), .A(n3642) );
  nand02 U1329 ( .Y(n3643), .A0(n3640), .A1(n3641) );
  inv01 U1330 ( .Y(n3633), .A(n3643) );
  nand02 U1331 ( .Y(s_fractb_28_o_6_), .A0(n3644), .A1(n3645) );
  inv01 U1332 ( .Y(n3646), .A(n3327) );
  inv01 U1333 ( .Y(n3647), .A(n5222) );
  inv01 U1334 ( .Y(n3648), .A(n5321) );
  inv01 U1335 ( .Y(n3649), .A(n4741) );
  nand02 U1336 ( .Y(n3650), .A0(n3646), .A1(n3647) );
  nand02 U1337 ( .Y(n3651), .A0(n3646), .A1(n3648) );
  nand02 U1338 ( .Y(n3652), .A0(n3647), .A1(n3649) );
  nand02 U1339 ( .Y(n3653), .A0(n3648), .A1(n3649) );
  nand02 U1340 ( .Y(n3654), .A0(n3650), .A1(n3651) );
  inv01 U1341 ( .Y(n3644), .A(n3654) );
  nand02 U1342 ( .Y(n3655), .A0(n3652), .A1(n3653) );
  inv01 U1343 ( .Y(n3645), .A(n3655) );
  nand02 U1344 ( .Y(s_fractb_28_o_11_), .A0(n3656), .A1(n3657) );
  inv01 U1345 ( .Y(n3658), .A(n____return128) );
  inv01 U1346 ( .Y(n3659), .A(n5223) );
  inv01 U1347 ( .Y(n3660), .A(n5357) );
  inv01 U1348 ( .Y(n3661), .A(n5358) );
  nand02 U1349 ( .Y(n3662), .A0(n3658), .A1(n3659) );
  nand02 U1350 ( .Y(n3663), .A0(n3658), .A1(n3660) );
  nand02 U1351 ( .Y(n3664), .A0(n3659), .A1(n3661) );
  nand02 U1352 ( .Y(n3665), .A0(n3660), .A1(n3661) );
  nand02 U1353 ( .Y(n3666), .A0(n3662), .A1(n3663) );
  inv01 U1354 ( .Y(n3656), .A(n3666) );
  nand02 U1355 ( .Y(n3667), .A0(n3664), .A1(n3665) );
  inv01 U1356 ( .Y(n3657), .A(n3667) );
  nand02 U1357 ( .Y(s_exp_o389_0_), .A0(n3668), .A1(n3669) );
  inv01 U1358 ( .Y(n3670), .A(n____return128) );
  inv01 U1359 ( .Y(n3671), .A(n5223) );
  inv01 U1360 ( .Y(n3672), .A(n5469) );
  inv01 U1361 ( .Y(n3673), .A(n4957) );
  nand02 U1362 ( .Y(n3674), .A0(n3670), .A1(n3671) );
  nand02 U1363 ( .Y(n3675), .A0(n3670), .A1(n3672) );
  nand02 U1364 ( .Y(n3676), .A0(n3671), .A1(n3673) );
  nand02 U1365 ( .Y(n3677), .A0(n3672), .A1(n3673) );
  nand02 U1366 ( .Y(n3678), .A0(n3674), .A1(n3675) );
  inv01 U1367 ( .Y(n3668), .A(n3678) );
  nand02 U1368 ( .Y(n3679), .A0(n3676), .A1(n3677) );
  inv01 U1369 ( .Y(n3669), .A(n3679) );
  nand02 U1370 ( .Y(s_fractb_28_o_13_), .A0(n3680), .A1(n3681) );
  inv01 U1371 ( .Y(n3682), .A(n____return128) );
  inv01 U1372 ( .Y(n3683), .A(n5223) );
  inv01 U1373 ( .Y(n3684), .A(n5355) );
  inv01 U1374 ( .Y(n3685), .A(n4739) );
  nand02 U1375 ( .Y(n3686), .A0(n3682), .A1(n3683) );
  nand02 U1376 ( .Y(n3687), .A0(n3682), .A1(n3684) );
  nand02 U1377 ( .Y(n3688), .A0(n3683), .A1(n3685) );
  nand02 U1378 ( .Y(n3689), .A0(n3684), .A1(n3685) );
  nand02 U1379 ( .Y(n3690), .A0(n3686), .A1(n3687) );
  inv01 U1380 ( .Y(n3680), .A(n3690) );
  nand02 U1381 ( .Y(n3691), .A0(n3688), .A1(n3689) );
  inv01 U1382 ( .Y(n3681), .A(n3691) );
  nand02 U1383 ( .Y(s_exp_o389_1_), .A0(n3692), .A1(n3693) );
  inv01 U1384 ( .Y(n3694), .A(n____return128) );
  inv01 U1385 ( .Y(n3695), .A(n5223) );
  inv01 U1386 ( .Y(n3696), .A(n4916) );
  inv01 U1387 ( .Y(n3697), .A(n4931) );
  nand02 U1388 ( .Y(n3698), .A0(n3694), .A1(n3695) );
  nand02 U1389 ( .Y(n3699), .A0(n3694), .A1(n3696) );
  nand02 U1390 ( .Y(n3700), .A0(n3695), .A1(n3697) );
  nand02 U1391 ( .Y(n3701), .A0(n3696), .A1(n3697) );
  nand02 U1392 ( .Y(n3702), .A0(n3698), .A1(n3699) );
  inv01 U1393 ( .Y(n3692), .A(n3702) );
  nand02 U1394 ( .Y(n3703), .A0(n3700), .A1(n3701) );
  inv01 U1395 ( .Y(n3693), .A(n3703) );
  nand02 U1396 ( .Y(s_fracta_28_o_14_), .A0(n3704), .A1(n3705) );
  inv01 U1397 ( .Y(n3706), .A(n3327) );
  inv01 U1398 ( .Y(n3707), .A(n5222) );
  inv01 U1399 ( .Y(n3708), .A(n4737) );
  inv01 U1400 ( .Y(n3709), .A(n5446) );
  nand02 U1401 ( .Y(n3710), .A0(n3706), .A1(n3707) );
  nand02 U1402 ( .Y(n3711), .A0(n3706), .A1(n3708) );
  nand02 U1403 ( .Y(n3712), .A0(n3707), .A1(n3709) );
  nand02 U1404 ( .Y(n3713), .A0(n3708), .A1(n3709) );
  nand02 U1405 ( .Y(n3714), .A0(n3710), .A1(n3711) );
  inv01 U1406 ( .Y(n3704), .A(n3714) );
  nand02 U1407 ( .Y(n3715), .A0(n3712), .A1(n3713) );
  inv01 U1408 ( .Y(n3705), .A(n3715) );
  nand02 U1409 ( .Y(s_fractb_28_o_9_), .A0(n3716), .A1(n3717) );
  inv01 U1410 ( .Y(n3718), .A(n____return128) );
  inv01 U1411 ( .Y(n3719), .A(n5222) );
  inv01 U1412 ( .Y(n3720), .A(n5316) );
  inv01 U1413 ( .Y(n3721), .A(n5317) );
  nand02 U1414 ( .Y(n3722), .A0(n3718), .A1(n3719) );
  nand02 U1415 ( .Y(n3723), .A0(n3718), .A1(n3720) );
  nand02 U1416 ( .Y(n3724), .A0(n3719), .A1(n3721) );
  nand02 U1417 ( .Y(n3725), .A0(n3720), .A1(n3721) );
  nand02 U1418 ( .Y(n3726), .A0(n3722), .A1(n3723) );
  inv01 U1419 ( .Y(n3716), .A(n3726) );
  nand02 U1420 ( .Y(n3727), .A0(n3724), .A1(n3725) );
  inv01 U1421 ( .Y(n3717), .A(n3727) );
  nand02 U1422 ( .Y(s_fracta_28_o_3_), .A0(n3728), .A1(n3729) );
  inv01 U1423 ( .Y(n3730), .A(n____return128) );
  inv01 U1424 ( .Y(n3731), .A(n5222) );
  inv01 U1425 ( .Y(n3732), .A(n5327) );
  inv01 U1426 ( .Y(n3733), .A(n5408) );
  nand02 U1427 ( .Y(n3734), .A0(n3730), .A1(n3731) );
  nand02 U1428 ( .Y(n3735), .A0(n3730), .A1(n3732) );
  nand02 U1429 ( .Y(n3736), .A0(n3731), .A1(n3733) );
  nand02 U1430 ( .Y(n3737), .A0(n3732), .A1(n3733) );
  nand02 U1431 ( .Y(n3738), .A0(n3734), .A1(n3735) );
  inv01 U1432 ( .Y(n3728), .A(n3738) );
  nand02 U1433 ( .Y(n3739), .A0(n3736), .A1(n3737) );
  inv01 U1434 ( .Y(n3729), .A(n3739) );
  nand02 U1435 ( .Y(s_exp_o389_6_), .A0(n3740), .A1(n3741) );
  inv01 U1436 ( .Y(n3742), .A(n3327) );
  inv01 U1437 ( .Y(n3743), .A(n5223) );
  inv01 U1438 ( .Y(n3744), .A(n4910) );
  inv01 U1439 ( .Y(n3745), .A(n4937) );
  nand02 U1440 ( .Y(n3746), .A0(n3742), .A1(n3743) );
  nand02 U1441 ( .Y(n3747), .A0(n3742), .A1(n3744) );
  nand02 U1442 ( .Y(n3748), .A0(n3743), .A1(n3745) );
  nand02 U1443 ( .Y(n3749), .A0(n3744), .A1(n3745) );
  nand02 U1444 ( .Y(n3750), .A0(n3746), .A1(n3747) );
  inv01 U1445 ( .Y(n3740), .A(n3750) );
  nand02 U1446 ( .Y(n3751), .A0(n3748), .A1(n3749) );
  inv01 U1447 ( .Y(n3741), .A(n3751) );
  nand02 U1448 ( .Y(s_fractb_28_o_12_), .A0(n3752), .A1(n3753) );
  inv01 U1449 ( .Y(n3754), .A(n____return128) );
  inv01 U1450 ( .Y(n3755), .A(n5223) );
  inv01 U1451 ( .Y(n3756), .A(n5356) );
  inv01 U1452 ( .Y(n3757), .A(n4743) );
  nand02 U1453 ( .Y(n3758), .A0(n3754), .A1(n3755) );
  nand02 U1454 ( .Y(n3759), .A0(n3754), .A1(n3756) );
  nand02 U1455 ( .Y(n3760), .A0(n3755), .A1(n3757) );
  nand02 U1456 ( .Y(n3761), .A0(n3756), .A1(n3757) );
  nand02 U1457 ( .Y(n3762), .A0(n3758), .A1(n3759) );
  inv01 U1458 ( .Y(n3752), .A(n3762) );
  nand02 U1459 ( .Y(n3763), .A0(n3760), .A1(n3761) );
  inv01 U1460 ( .Y(n3753), .A(n3763) );
  nand02 U1461 ( .Y(s_fractb_28_o_7_), .A0(n3764), .A1(n3765) );
  inv01 U1462 ( .Y(n3766), .A(n3327) );
  inv01 U1463 ( .Y(n3767), .A(n5223) );
  inv01 U1464 ( .Y(n3768), .A(n5320) );
  inv01 U1465 ( .Y(n3769), .A(n4733) );
  nand02 U1466 ( .Y(n3770), .A0(n3766), .A1(n3767) );
  nand02 U1467 ( .Y(n3771), .A0(n3766), .A1(n3768) );
  nand02 U1468 ( .Y(n3772), .A0(n3767), .A1(n3769) );
  nand02 U1469 ( .Y(n3773), .A0(n3768), .A1(n3769) );
  nand02 U1470 ( .Y(n3774), .A0(n3770), .A1(n3771) );
  inv01 U1471 ( .Y(n3764), .A(n3774) );
  nand02 U1472 ( .Y(n3775), .A0(n3772), .A1(n3773) );
  inv01 U1473 ( .Y(n3765), .A(n3775) );
  nand02 U1474 ( .Y(s_fractb_28_o_15_), .A0(n3776), .A1(n3777) );
  inv01 U1475 ( .Y(n3778), .A(n3327) );
  inv01 U1476 ( .Y(n3779), .A(n5222) );
  inv01 U1477 ( .Y(n3780), .A(n5352) );
  inv01 U1478 ( .Y(n3781), .A(n5353) );
  nand02 U1479 ( .Y(n3782), .A0(n3778), .A1(n3779) );
  nand02 U1480 ( .Y(n3783), .A0(n3778), .A1(n3780) );
  nand02 U1481 ( .Y(n3784), .A0(n3779), .A1(n3781) );
  nand02 U1482 ( .Y(n3785), .A0(n3780), .A1(n3781) );
  nand02 U1483 ( .Y(n3786), .A0(n3782), .A1(n3783) );
  inv01 U1484 ( .Y(n3776), .A(n3786) );
  nand02 U1485 ( .Y(n3787), .A0(n3784), .A1(n3785) );
  inv01 U1486 ( .Y(n3777), .A(n3787) );
  nand02 U1487 ( .Y(s_fractb_28_o_3_), .A0(n3788), .A1(n3789) );
  inv01 U1488 ( .Y(n3790), .A(n3327) );
  inv01 U1489 ( .Y(n3791), .A(n5222) );
  inv01 U1490 ( .Y(n3792), .A(n5326) );
  inv01 U1491 ( .Y(n3793), .A(n5327) );
  nand02 U1492 ( .Y(n3794), .A0(n3790), .A1(n3791) );
  nand02 U1493 ( .Y(n3795), .A0(n3790), .A1(n3792) );
  nand02 U1494 ( .Y(n3796), .A0(n3791), .A1(n3793) );
  nand02 U1495 ( .Y(n3797), .A0(n3792), .A1(n3793) );
  nand02 U1496 ( .Y(n3798), .A0(n3794), .A1(n3795) );
  inv01 U1497 ( .Y(n3788), .A(n3798) );
  nand02 U1498 ( .Y(n3799), .A0(n3796), .A1(n3797) );
  inv01 U1499 ( .Y(n3789), .A(n3799) );
  nand02 U1500 ( .Y(s_fractb_28_o_4_), .A0(n3800), .A1(n3801) );
  inv01 U1501 ( .Y(n3802), .A(n3327) );
  inv01 U1502 ( .Y(n3803), .A(n5222) );
  inv01 U1503 ( .Y(n3804), .A(n5324) );
  inv01 U1504 ( .Y(n3805), .A(n5325) );
  nand02 U1505 ( .Y(n3806), .A0(n3802), .A1(n3803) );
  nand02 U1506 ( .Y(n3807), .A0(n3802), .A1(n3804) );
  nand02 U1507 ( .Y(n3808), .A0(n3803), .A1(n3805) );
  nand02 U1508 ( .Y(n3809), .A0(n3804), .A1(n3805) );
  nand02 U1509 ( .Y(n3810), .A0(n3806), .A1(n3807) );
  inv01 U1510 ( .Y(n3800), .A(n3810) );
  nand02 U1511 ( .Y(n3811), .A0(n3808), .A1(n3809) );
  inv01 U1512 ( .Y(n3801), .A(n3811) );
  nand02 U1513 ( .Y(s_fracta_28_o_11_), .A0(n3812), .A1(n3813) );
  inv01 U1514 ( .Y(n3814), .A(n3327) );
  inv01 U1515 ( .Y(n3815), .A(n5222) );
  inv01 U1516 ( .Y(n3816), .A(n5358) );
  inv01 U1517 ( .Y(n3817), .A(n5453) );
  nand02 U1518 ( .Y(n3818), .A0(n3814), .A1(n3815) );
  nand02 U1519 ( .Y(n3819), .A0(n3814), .A1(n3816) );
  nand02 U1520 ( .Y(n3820), .A0(n3815), .A1(n3817) );
  nand02 U1521 ( .Y(n3821), .A0(n3816), .A1(n3817) );
  nand02 U1522 ( .Y(n3822), .A0(n3818), .A1(n3819) );
  inv01 U1523 ( .Y(n3812), .A(n3822) );
  nand02 U1524 ( .Y(n3823), .A0(n3820), .A1(n3821) );
  inv01 U1525 ( .Y(n3813), .A(n3823) );
  nand02 U1526 ( .Y(s_fracta_28_o_6_), .A0(n3824), .A1(n3825) );
  inv01 U1527 ( .Y(n3826), .A(n3327) );
  inv01 U1528 ( .Y(n3827), .A(n5222) );
  inv01 U1529 ( .Y(n3828), .A(n4741) );
  inv01 U1530 ( .Y(n3829), .A(n5389) );
  nand02 U1531 ( .Y(n3830), .A0(n3826), .A1(n3827) );
  nand02 U1532 ( .Y(n3831), .A0(n3826), .A1(n3828) );
  nand02 U1533 ( .Y(n3832), .A0(n3827), .A1(n3829) );
  nand02 U1534 ( .Y(n3833), .A0(n3828), .A1(n3829) );
  nand02 U1535 ( .Y(n3834), .A0(n3830), .A1(n3831) );
  inv01 U1536 ( .Y(n3824), .A(n3834) );
  nand02 U1537 ( .Y(n3835), .A0(n3832), .A1(n3833) );
  inv01 U1538 ( .Y(n3825), .A(n3835) );
  nand02 U1539 ( .Y(s_fracta_28_o_4_), .A0(n3836), .A1(n3837) );
  inv01 U1540 ( .Y(n3838), .A(n3327) );
  inv01 U1541 ( .Y(n3839), .A(n5222) );
  inv01 U1542 ( .Y(n3840), .A(n5325) );
  inv01 U1543 ( .Y(n3841), .A(n5403) );
  nand02 U1544 ( .Y(n3842), .A0(n3838), .A1(n3839) );
  nand02 U1545 ( .Y(n3843), .A0(n3838), .A1(n3840) );
  nand02 U1546 ( .Y(n3844), .A0(n3839), .A1(n3841) );
  nand02 U1547 ( .Y(n3845), .A0(n3840), .A1(n3841) );
  nand02 U1548 ( .Y(n3846), .A0(n3842), .A1(n3843) );
  inv01 U1549 ( .Y(n3836), .A(n3846) );
  nand02 U1550 ( .Y(n3847), .A0(n3844), .A1(n3845) );
  inv01 U1551 ( .Y(n3837), .A(n3847) );
  nand02 U1552 ( .Y(s_fracta_28_o_5_), .A0(n3848), .A1(n3849) );
  inv01 U1553 ( .Y(n3850), .A(n3327) );
  inv01 U1554 ( .Y(n3851), .A(n5222) );
  inv01 U1555 ( .Y(n3852), .A(n5323) );
  inv01 U1556 ( .Y(n3853), .A(n5398) );
  nand02 U1557 ( .Y(n3854), .A0(n3850), .A1(n3851) );
  nand02 U1558 ( .Y(n3855), .A0(n3850), .A1(n3852) );
  nand02 U1559 ( .Y(n3856), .A0(n3851), .A1(n3853) );
  nand02 U1560 ( .Y(n3857), .A0(n3852), .A1(n3853) );
  nand02 U1561 ( .Y(n3858), .A0(n3854), .A1(n3855) );
  inv01 U1562 ( .Y(n3848), .A(n3858) );
  nand02 U1563 ( .Y(n3859), .A0(n3856), .A1(n3857) );
  inv01 U1564 ( .Y(n3849), .A(n3859) );
  nand02 U1565 ( .Y(s_fracta_28_o_15_), .A0(n3860), .A1(n3861) );
  inv01 U1566 ( .Y(n3862), .A(n3327) );
  inv01 U1567 ( .Y(n3863), .A(n5222) );
  inv01 U1568 ( .Y(n3864), .A(n5353) );
  inv01 U1569 ( .Y(n3865), .A(n5445) );
  nand02 U1570 ( .Y(n3866), .A0(n3862), .A1(n3863) );
  nand02 U1571 ( .Y(n3867), .A0(n3862), .A1(n3864) );
  nand02 U1572 ( .Y(n3868), .A0(n3863), .A1(n3865) );
  nand02 U1573 ( .Y(n3869), .A0(n3864), .A1(n3865) );
  nand02 U1574 ( .Y(n3870), .A0(n3866), .A1(n3867) );
  inv01 U1575 ( .Y(n3860), .A(n3870) );
  nand02 U1576 ( .Y(n3871), .A0(n3868), .A1(n3869) );
  inv01 U1577 ( .Y(n3861), .A(n3871) );
  or03 U1578 ( .Y(n3872), .A0(n5237), .A1(n5235), .A2(n5236) );
  inv01 U1579 ( .Y(n3873), .A(n3872) );
  or03 U1580 ( .Y(n3874), .A0(n5228), .A1(n5226), .A2(n5227) );
  inv01 U1581 ( .Y(n3875), .A(n3874) );
  nand02 U1582 ( .Y(s_fractb_28_o_21_), .A0(n3876), .A1(n3877) );
  inv01 U1583 ( .Y(n3878), .A(n5204) );
  inv01 U1584 ( .Y(n3879), .A(n4860) );
  inv01 U1585 ( .Y(n3880), .A(n5342) );
  inv01 U1586 ( .Y(n3881), .A(n3327) );
  nand02 U1587 ( .Y(n3876), .A0(n3878), .A1(n3879) );
  nand02 U1588 ( .Y(n3877), .A0(n3880), .A1(n3881) );
  nand02 U1589 ( .Y(s_fractb_28_o_18_), .A0(n3882), .A1(n3883) );
  inv01 U1590 ( .Y(n3884), .A(n5205) );
  inv01 U1591 ( .Y(n3885), .A(n5347) );
  inv01 U1592 ( .Y(n3886), .A(n5346) );
  inv01 U1593 ( .Y(n3887), .A(n3327) );
  nand02 U1594 ( .Y(n3882), .A0(n3884), .A1(n3885) );
  nand02 U1595 ( .Y(n3883), .A0(n3886), .A1(n3887) );
  nand02 U1596 ( .Y(s_fractb_28_o_23_), .A0(n3888), .A1(n3889) );
  inv01 U1597 ( .Y(n3890), .A(n4876) );
  inv01 U1598 ( .Y(n3891), .A(n5337) );
  inv01 U1599 ( .Y(n3892), .A(n5336) );
  inv01 U1600 ( .Y(n3893), .A(n3327) );
  nand02 U1601 ( .Y(n3888), .A0(n3890), .A1(n3891) );
  nand02 U1602 ( .Y(n3889), .A0(n3892), .A1(n3893) );
  nand02 U1603 ( .Y(s_fractb_28_o_19_), .A0(n3894), .A1(n3895) );
  inv01 U1604 ( .Y(n3896), .A(n5204) );
  inv01 U1605 ( .Y(n3897), .A(n4878) );
  inv01 U1606 ( .Y(n3898), .A(n5345) );
  inv01 U1607 ( .Y(n3899), .A(n3327) );
  nand02 U1608 ( .Y(n3894), .A0(n3896), .A1(n3897) );
  nand02 U1609 ( .Y(n3895), .A0(n3898), .A1(n3899) );
  nand02 U1610 ( .Y(s_fractb_28_o_17_), .A0(n3900), .A1(n3901) );
  inv01 U1611 ( .Y(n3902), .A(n5204) );
  inv01 U1612 ( .Y(n3903), .A(n5349) );
  inv01 U1613 ( .Y(n3904), .A(n5348) );
  inv01 U1614 ( .Y(n3905), .A(n3327) );
  nand02 U1615 ( .Y(n3900), .A0(n3902), .A1(n3903) );
  nand02 U1616 ( .Y(n3901), .A0(n3904), .A1(n3905) );
  nand02 U1617 ( .Y(s_fractb_28_o_16_), .A0(n3906), .A1(n3907) );
  inv01 U1618 ( .Y(n3908), .A(n5204) );
  inv01 U1619 ( .Y(n3909), .A(n5351) );
  inv01 U1620 ( .Y(n3910), .A(n5350) );
  inv01 U1621 ( .Y(n3911), .A(n3327) );
  nand02 U1622 ( .Y(n3906), .A0(n3908), .A1(n3909) );
  nand02 U1623 ( .Y(n3907), .A0(n3910), .A1(n3911) );
  nand02 U1624 ( .Y(s_fractb_28_o_24_), .A0(n3912), .A1(n3913) );
  inv01 U1625 ( .Y(n3914), .A(n4876) );
  inv01 U1626 ( .Y(n3915), .A(n5335) );
  inv01 U1627 ( .Y(n3916), .A(n5334) );
  inv01 U1628 ( .Y(n3917), .A(n____return128) );
  nand02 U1629 ( .Y(n3912), .A0(n3914), .A1(n3915) );
  nand02 U1630 ( .Y(n3913), .A0(n3916), .A1(n3917) );
  nand02 U1631 ( .Y(s_fractb_28_o_26_), .A0(n3918), .A1(n3919) );
  inv01 U1632 ( .Y(n3920), .A(n4876) );
  inv01 U1633 ( .Y(n3921), .A(n5330) );
  inv01 U1634 ( .Y(n3922), .A(n5329) );
  inv01 U1635 ( .Y(n3923), .A(n____return128) );
  nand02 U1636 ( .Y(n3918), .A0(n3920), .A1(n3921) );
  nand02 U1637 ( .Y(n3919), .A0(n3922), .A1(n3923) );
  nand02 U1638 ( .Y(s_fractb_28_o_22_), .A0(n3924), .A1(n3925) );
  inv01 U1639 ( .Y(n3926), .A(n5205) );
  inv01 U1640 ( .Y(n3927), .A(n5340) );
  inv01 U1641 ( .Y(n3928), .A(n5339) );
  inv01 U1642 ( .Y(n3929), .A(n____return128) );
  nand02 U1643 ( .Y(n3924), .A0(n3926), .A1(n3927) );
  nand02 U1644 ( .Y(n3925), .A0(n3928), .A1(n3929) );
  nand02 U1645 ( .Y(s_fractb_28_o_20_), .A0(n3930), .A1(n3931) );
  inv01 U1646 ( .Y(n3932), .A(n5205) );
  inv01 U1647 ( .Y(n3933), .A(n4863) );
  inv01 U1648 ( .Y(n3934), .A(n5343) );
  inv01 U1649 ( .Y(n3935), .A(n____return128) );
  nand02 U1650 ( .Y(n3930), .A0(n3932), .A1(n3933) );
  nand02 U1651 ( .Y(n3931), .A0(n3934), .A1(n3935) );
  nand02 U1652 ( .Y(s_fractb_28_o_25_), .A0(n3936), .A1(n3937) );
  inv01 U1653 ( .Y(n3938), .A(n4876) );
  inv01 U1654 ( .Y(n3939), .A(n5333) );
  inv01 U1655 ( .Y(n3940), .A(n5332) );
  inv01 U1656 ( .Y(n3941), .A(n____return128) );
  nand02 U1657 ( .Y(n3936), .A0(n3938), .A1(n3939) );
  nand02 U1658 ( .Y(n3937), .A0(n3940), .A1(n3941) );
  buf02 U1659 ( .Y(n4876), .A(n5331) );
  inv02 U1660 ( .Y(n5340), .A(n5396) );
  nand02 U1661 ( .Y(n3942), .A0(n5310), .A1(n5152) );
  inv02 U1662 ( .Y(n3943), .A(n3942) );
  nand02 U1663 ( .Y(U403_U4_Z_1), .A0(n3944), .A1(n3945) );
  inv01 U1664 ( .Y(n3946), .A(n____return128) );
  inv01 U1665 ( .Y(n3947), .A(n5223) );
  inv01 U1666 ( .Y(n3948), .A(n4931) );
  inv01 U1667 ( .Y(n3949), .A(n4916) );
  nand02 U1668 ( .Y(n3950), .A0(n3946), .A1(n3947) );
  nand02 U1669 ( .Y(n3951), .A0(n3946), .A1(n3948) );
  nand02 U1670 ( .Y(n3952), .A0(n3947), .A1(n3949) );
  nand02 U1671 ( .Y(n3953), .A0(n3948), .A1(n3949) );
  nand02 U1672 ( .Y(n3954), .A0(n3950), .A1(n3951) );
  inv01 U1673 ( .Y(n3944), .A(n3954) );
  nand02 U1674 ( .Y(n3955), .A0(n3952), .A1(n3953) );
  inv01 U1675 ( .Y(n3945), .A(n3955) );
  nand02 U1676 ( .Y(U403_U4_Z_6), .A0(n3956), .A1(n3957) );
  inv01 U1677 ( .Y(n3958), .A(n____return128) );
  inv01 U1678 ( .Y(n3959), .A(n5223) );
  inv01 U1679 ( .Y(n3960), .A(n4937) );
  inv01 U1680 ( .Y(n3961), .A(n4910) );
  nand02 U1681 ( .Y(n3962), .A0(n3958), .A1(n3959) );
  nand02 U1682 ( .Y(n3963), .A0(n3958), .A1(n3960) );
  nand02 U1683 ( .Y(n3964), .A0(n3959), .A1(n3961) );
  nand02 U1684 ( .Y(n3965), .A0(n3960), .A1(n3961) );
  nand02 U1685 ( .Y(n3966), .A0(n3962), .A1(n3963) );
  inv01 U1686 ( .Y(n3956), .A(n3966) );
  nand02 U1687 ( .Y(n3967), .A0(n3964), .A1(n3965) );
  inv01 U1688 ( .Y(n3957), .A(n3967) );
  nand02 U1689 ( .Y(U403_U4_Z_4), .A0(n3968), .A1(n3969) );
  inv01 U1690 ( .Y(n3970), .A(n3327) );
  inv01 U1691 ( .Y(n3971), .A(n5223) );
  inv01 U1692 ( .Y(n3972), .A(n4941) );
  inv01 U1693 ( .Y(n3973), .A(n4928) );
  nand02 U1694 ( .Y(n3974), .A0(n3970), .A1(n3971) );
  nand02 U1695 ( .Y(n3975), .A0(n3970), .A1(n3972) );
  nand02 U1696 ( .Y(n3976), .A0(n3971), .A1(n3973) );
  nand02 U1697 ( .Y(n3977), .A0(n3972), .A1(n3973) );
  nand02 U1698 ( .Y(n3978), .A0(n3974), .A1(n3975) );
  inv01 U1699 ( .Y(n3968), .A(n3978) );
  nand02 U1700 ( .Y(n3979), .A0(n3976), .A1(n3977) );
  inv01 U1701 ( .Y(n3969), .A(n3979) );
  nand02 U1702 ( .Y(U403_U4_Z_5), .A0(n3980), .A1(n3981) );
  inv01 U1703 ( .Y(n3982), .A(n____return128) );
  inv01 U1704 ( .Y(n3983), .A(n5223) );
  inv01 U1705 ( .Y(n3984), .A(n4933) );
  inv01 U1706 ( .Y(n3985), .A(n4919) );
  nand02 U1707 ( .Y(n3986), .A0(n3982), .A1(n3983) );
  nand02 U1708 ( .Y(n3987), .A0(n3982), .A1(n3984) );
  nand02 U1709 ( .Y(n3988), .A0(n3983), .A1(n3985) );
  nand02 U1710 ( .Y(n3989), .A0(n3984), .A1(n3985) );
  nand02 U1711 ( .Y(n3990), .A0(n3986), .A1(n3987) );
  inv01 U1712 ( .Y(n3980), .A(n3990) );
  nand02 U1713 ( .Y(n3991), .A0(n3988), .A1(n3989) );
  inv01 U1714 ( .Y(n3981), .A(n3991) );
  nand02 U1715 ( .Y(U403_U4_Z_3), .A0(n3992), .A1(n3993) );
  inv01 U1716 ( .Y(n3994), .A(n____return128) );
  inv01 U1717 ( .Y(n3995), .A(n5222) );
  inv01 U1718 ( .Y(n3996), .A(n4935) );
  inv01 U1719 ( .Y(n3997), .A(n4913) );
  nand02 U1720 ( .Y(n3998), .A0(n3994), .A1(n3995) );
  nand02 U1721 ( .Y(n3999), .A0(n3994), .A1(n3996) );
  nand02 U1722 ( .Y(n4000), .A0(n3995), .A1(n3997) );
  nand02 U1723 ( .Y(n4001), .A0(n3996), .A1(n3997) );
  nand02 U1724 ( .Y(n4002), .A0(n3998), .A1(n3999) );
  inv01 U1725 ( .Y(n3992), .A(n4002) );
  nand02 U1726 ( .Y(n4003), .A0(n4000), .A1(n4001) );
  inv01 U1727 ( .Y(n3993), .A(n4003) );
  nand02 U1728 ( .Y(U403_U4_Z_2), .A0(n4004), .A1(n4005) );
  inv01 U1729 ( .Y(n4007), .A(n5222) );
  inv01 U1730 ( .Y(n4008), .A(n4939) );
  inv01 U1731 ( .Y(n4009), .A(n4922) );
  nand02 U1732 ( .Y(n4010), .A0(n4006), .A1(n4007) );
  nand02 U1733 ( .Y(n4011), .A0(n4006), .A1(n4008) );
  nand02 U1734 ( .Y(n4012), .A0(n4007), .A1(n4009) );
  nand02 U1735 ( .Y(n4013), .A0(n4008), .A1(n4009) );
  nand02 U1736 ( .Y(n4014), .A0(n4010), .A1(n4011) );
  inv01 U1737 ( .Y(n4004), .A(n4014) );
  nand02 U1738 ( .Y(n4015), .A0(n4012), .A1(n4013) );
  inv01 U1739 ( .Y(n4005), .A(n4015) );
  nor02 U1740 ( .Y(n5300), .A0(n5228), .A1(n4016) );
  nor02 U1741 ( .Y(n4017), .A0(n5227), .A1(n5226) );
  inv01 U1742 ( .Y(n4016), .A(n4017) );
  nand02 U1743 ( .Y(U403_U4_Z_7), .A0(n4018), .A1(n4019) );
  inv01 U1744 ( .Y(n4020), .A(n3327) );
  inv01 U1745 ( .Y(n4021), .A(n5222) );
  inv01 U1746 ( .Y(n4022), .A(n4943) );
  inv01 U1747 ( .Y(n4023), .A(n4925) );
  nand02 U1748 ( .Y(n4024), .A0(n4020), .A1(n4021) );
  nand02 U1749 ( .Y(n4025), .A0(n4020), .A1(n4022) );
  nand02 U1750 ( .Y(n4026), .A0(n4021), .A1(n4023) );
  nand02 U1751 ( .Y(n4027), .A0(n4022), .A1(n4023) );
  nand02 U1752 ( .Y(n4028), .A0(n4024), .A1(n4025) );
  inv01 U1753 ( .Y(n4018), .A(n4028) );
  nand02 U1754 ( .Y(n4029), .A0(n4026), .A1(n4027) );
  inv01 U1755 ( .Y(n4019), .A(n4029) );
  inv01 U1756 ( .Y(n5423), .A(n4030) );
  nor02 U1757 ( .Y(n4031), .A0(n5201), .A1(n4929) );
  nor02 U1758 ( .Y(n4032), .A0(n5284), .A1(n5219) );
  nor02 U1759 ( .Y(n4033), .A0(n5180), .A1(n5220) );
  nor02 U1760 ( .Y(n4030), .A0(n4033), .A1(n4034) );
  nor02 U1761 ( .Y(n4035), .A0(n4031), .A1(n4032) );
  inv01 U1762 ( .Y(n4034), .A(n4035) );
  inv01 U1763 ( .Y(n5414), .A(n4036) );
  nor02 U1764 ( .Y(n4037), .A0(n5284), .A1(n5220) );
  nor02 U1765 ( .Y(n4038), .A0(n5201), .A1(n5219) );
  inv01 U1766 ( .Y(n4039), .A(n3394) );
  nor02 U1767 ( .Y(n4036), .A0(n4039), .A1(n4040) );
  nor02 U1768 ( .Y(n4041), .A0(n4037), .A1(n4038) );
  inv01 U1769 ( .Y(n4040), .A(n4041) );
  inv02 U1770 ( .Y(n5284), .A(n5462) );
  nand02 U1771 ( .Y(n4042), .A0(n5141), .A1(n5285) );
  inv02 U1772 ( .Y(n4043), .A(n4042) );
  nand02 U1773 ( .Y(n4044), .A0(n3396), .A1(n5150) );
  inv02 U1774 ( .Y(n4045), .A(n4044) );
  nand02 U1775 ( .Y(n4046), .A0(n5304), .A1(n5143) );
  inv02 U1776 ( .Y(n4047), .A(n4046) );
  nand02 U1777 ( .Y(n5367), .A0(n4048), .A1(n4049) );
  inv02 U1778 ( .Y(n4050), .A(n5372) );
  inv02 U1779 ( .Y(n4051), .A(n5371) );
  inv02 U1780 ( .Y(n4052), .A(n5369) );
  inv02 U1781 ( .Y(n4053), .A(n5216) );
  inv02 U1782 ( .Y(n4054), .A(n3408) );
  inv02 U1783 ( .Y(n4055), .A(n5218) );
  nand02 U1784 ( .Y(n4056), .A0(n4052), .A1(n4057) );
  nand02 U1785 ( .Y(n4058), .A0(n4053), .A1(n4059) );
  nand02 U1786 ( .Y(n4060), .A0(n4054), .A1(n4061) );
  nand02 U1787 ( .Y(n4062), .A0(n4054), .A1(n4063) );
  nand02 U1788 ( .Y(n4064), .A0(n4055), .A1(n4065) );
  nand02 U1789 ( .Y(n4066), .A0(n4055), .A1(n4067) );
  nand02 U1790 ( .Y(n4068), .A0(n4055), .A1(n4069) );
  nand02 U1791 ( .Y(n4070), .A0(n4055), .A1(n4071) );
  nand02 U1792 ( .Y(n4072), .A0(n4050), .A1(n4051) );
  inv01 U1793 ( .Y(n4057), .A(n4072) );
  nand02 U1794 ( .Y(n4073), .A0(n4050), .A1(n4051) );
  inv01 U1795 ( .Y(n4059), .A(n4073) );
  nand02 U1796 ( .Y(n4074), .A0(n4050), .A1(n4052) );
  inv01 U1797 ( .Y(n4061), .A(n4074) );
  nand02 U1798 ( .Y(n4075), .A0(n4050), .A1(n4053) );
  inv01 U1799 ( .Y(n4063), .A(n4075) );
  nand02 U1800 ( .Y(n4076), .A0(n4051), .A1(n4052) );
  inv01 U1801 ( .Y(n4065), .A(n4076) );
  nand02 U1802 ( .Y(n4077), .A0(n4051), .A1(n4053) );
  inv01 U1803 ( .Y(n4067), .A(n4077) );
  nand02 U1804 ( .Y(n4078), .A0(n4052), .A1(n4054) );
  inv01 U1805 ( .Y(n4069), .A(n4078) );
  nand02 U1806 ( .Y(n4079), .A0(n4053), .A1(n4054) );
  inv01 U1807 ( .Y(n4071), .A(n4079) );
  nand02 U1808 ( .Y(n4080), .A0(n4056), .A1(n4058) );
  inv01 U1809 ( .Y(n4081), .A(n4080) );
  nand02 U1810 ( .Y(n4082), .A0(n4060), .A1(n4062) );
  inv01 U1811 ( .Y(n4083), .A(n4082) );
  nand02 U1812 ( .Y(n4084), .A0(n4081), .A1(n4083) );
  inv01 U1813 ( .Y(n4048), .A(n4084) );
  nand02 U1814 ( .Y(n4085), .A0(n4064), .A1(n4066) );
  inv01 U1815 ( .Y(n4086), .A(n4085) );
  nand02 U1816 ( .Y(n4087), .A0(n4068), .A1(n4070) );
  inv01 U1817 ( .Y(n4088), .A(n4087) );
  nand02 U1818 ( .Y(n4089), .A0(n4086), .A1(n4088) );
  inv01 U1819 ( .Y(n4049), .A(n4089) );
  nand02 U1820 ( .Y(n5385), .A0(n4090), .A1(n4091) );
  inv02 U1821 ( .Y(n4092), .A(n5388) );
  inv02 U1822 ( .Y(n4093), .A(n5387) );
  inv02 U1823 ( .Y(n4094), .A(n5386) );
  inv02 U1824 ( .Y(n4095), .A(n5216) );
  inv02 U1825 ( .Y(n4096), .A(n3407) );
  inv02 U1826 ( .Y(n4097), .A(n5218) );
  nand02 U1827 ( .Y(n4098), .A0(n4094), .A1(n4099) );
  nand02 U1828 ( .Y(n4100), .A0(n4095), .A1(n4101) );
  nand02 U1829 ( .Y(n4102), .A0(n4096), .A1(n4103) );
  nand02 U1830 ( .Y(n4104), .A0(n4096), .A1(n4105) );
  nand02 U1831 ( .Y(n4106), .A0(n4097), .A1(n4107) );
  nand02 U1832 ( .Y(n4108), .A0(n4097), .A1(n4109) );
  nand02 U1833 ( .Y(n4110), .A0(n4097), .A1(n4111) );
  nand02 U1834 ( .Y(n4112), .A0(n4097), .A1(n4113) );
  nand02 U1835 ( .Y(n4114), .A0(n4092), .A1(n4093) );
  inv01 U1836 ( .Y(n4099), .A(n4114) );
  nand02 U1837 ( .Y(n4115), .A0(n4092), .A1(n4093) );
  inv01 U1838 ( .Y(n4101), .A(n4115) );
  nand02 U1839 ( .Y(n4116), .A0(n4092), .A1(n4094) );
  inv01 U1840 ( .Y(n4103), .A(n4116) );
  nand02 U1841 ( .Y(n4117), .A0(n4092), .A1(n4095) );
  inv01 U1842 ( .Y(n4105), .A(n4117) );
  nand02 U1843 ( .Y(n4118), .A0(n4093), .A1(n4094) );
  inv01 U1844 ( .Y(n4107), .A(n4118) );
  nand02 U1845 ( .Y(n4119), .A0(n4093), .A1(n4095) );
  inv01 U1846 ( .Y(n4109), .A(n4119) );
  nand02 U1847 ( .Y(n4120), .A0(n4094), .A1(n4096) );
  inv01 U1848 ( .Y(n4111), .A(n4120) );
  nand02 U1849 ( .Y(n4121), .A0(n4095), .A1(n4096) );
  inv01 U1850 ( .Y(n4113), .A(n4121) );
  nand02 U1851 ( .Y(n4122), .A0(n4098), .A1(n4100) );
  inv01 U1852 ( .Y(n4123), .A(n4122) );
  nand02 U1853 ( .Y(n4124), .A0(n4102), .A1(n4104) );
  inv01 U1854 ( .Y(n4125), .A(n4124) );
  nand02 U1855 ( .Y(n4126), .A0(n4123), .A1(n4125) );
  inv01 U1856 ( .Y(n4090), .A(n4126) );
  nand02 U1857 ( .Y(n4127), .A0(n4106), .A1(n4108) );
  inv01 U1858 ( .Y(n4128), .A(n4127) );
  nand02 U1859 ( .Y(n4129), .A0(n4110), .A1(n4112) );
  inv01 U1860 ( .Y(n4130), .A(n4129) );
  nand02 U1861 ( .Y(n4131), .A0(n4128), .A1(n4130) );
  inv01 U1862 ( .Y(n4091), .A(n4131) );
  nand02 U1863 ( .Y(n5405), .A0(n4132), .A1(n4133) );
  inv02 U1864 ( .Y(n4134), .A(n5407) );
  inv02 U1865 ( .Y(n4135), .A(n5406) );
  inv02 U1866 ( .Y(n4136), .A(n5375) );
  inv02 U1867 ( .Y(n4137), .A(n5216) );
  inv02 U1868 ( .Y(n4138), .A(n5197) );
  inv02 U1869 ( .Y(n4139), .A(n5218) );
  nand02 U1870 ( .Y(n4140), .A0(n4136), .A1(n4141) );
  nand02 U1871 ( .Y(n4142), .A0(n4137), .A1(n4143) );
  nand02 U1872 ( .Y(n4144), .A0(n4138), .A1(n4145) );
  nand02 U1873 ( .Y(n4146), .A0(n4138), .A1(n4147) );
  nand02 U1874 ( .Y(n4148), .A0(n4139), .A1(n4149) );
  nand02 U1875 ( .Y(n4150), .A0(n4139), .A1(n4151) );
  nand02 U1876 ( .Y(n4152), .A0(n4139), .A1(n4153) );
  nand02 U1877 ( .Y(n4154), .A0(n4139), .A1(n4155) );
  nand02 U1878 ( .Y(n4156), .A0(n4134), .A1(n4135) );
  inv01 U1879 ( .Y(n4141), .A(n4156) );
  nand02 U1880 ( .Y(n4157), .A0(n4134), .A1(n4135) );
  inv01 U1881 ( .Y(n4143), .A(n4157) );
  nand02 U1882 ( .Y(n4158), .A0(n4134), .A1(n4136) );
  inv01 U1883 ( .Y(n4145), .A(n4158) );
  nand02 U1884 ( .Y(n4159), .A0(n4134), .A1(n4137) );
  inv01 U1885 ( .Y(n4147), .A(n4159) );
  nand02 U1886 ( .Y(n4160), .A0(n4135), .A1(n4136) );
  inv01 U1887 ( .Y(n4149), .A(n4160) );
  nand02 U1888 ( .Y(n4161), .A0(n4135), .A1(n4137) );
  inv01 U1889 ( .Y(n4151), .A(n4161) );
  nand02 U1890 ( .Y(n4162), .A0(n4136), .A1(n4138) );
  inv01 U1891 ( .Y(n4153), .A(n4162) );
  nand02 U1892 ( .Y(n4163), .A0(n4137), .A1(n4138) );
  inv01 U1893 ( .Y(n4155), .A(n4163) );
  nand02 U1894 ( .Y(n4164), .A0(n4140), .A1(n4142) );
  inv01 U1895 ( .Y(n4165), .A(n4164) );
  nand02 U1896 ( .Y(n4166), .A0(n4144), .A1(n4146) );
  inv01 U1897 ( .Y(n4167), .A(n4166) );
  nand02 U1898 ( .Y(n4168), .A0(n4165), .A1(n4167) );
  inv01 U1899 ( .Y(n4132), .A(n4168) );
  nand02 U1900 ( .Y(n4169), .A0(n4148), .A1(n4150) );
  inv01 U1901 ( .Y(n4170), .A(n4169) );
  nand02 U1902 ( .Y(n4171), .A0(n4152), .A1(n4154) );
  inv01 U1903 ( .Y(n4172), .A(n4171) );
  nand02 U1904 ( .Y(n4173), .A0(n4170), .A1(n4172) );
  inv01 U1905 ( .Y(n4133), .A(n4173) );
  nand02 U1906 ( .Y(n5421), .A0(n4174), .A1(n4175) );
  inv02 U1907 ( .Y(n4176), .A(n5395) );
  inv02 U1908 ( .Y(n4177), .A(n5423) );
  inv02 U1909 ( .Y(n4178), .A(n5422) );
  inv02 U1910 ( .Y(n4179), .A(n5197) );
  inv02 U1911 ( .Y(n4180), .A(n5218) );
  inv02 U1912 ( .Y(n4181), .A(n5216) );
  nand02 U1913 ( .Y(n4182), .A0(n4178), .A1(n4183) );
  nand02 U1914 ( .Y(n4184), .A0(n4179), .A1(n4185) );
  nand02 U1915 ( .Y(n4186), .A0(n4180), .A1(n4187) );
  nand02 U1916 ( .Y(n4188), .A0(n4180), .A1(n4189) );
  nand02 U1917 ( .Y(n4190), .A0(n4181), .A1(n4191) );
  nand02 U1918 ( .Y(n4192), .A0(n4181), .A1(n4193) );
  nand02 U1919 ( .Y(n4194), .A0(n4181), .A1(n4195) );
  nand02 U1920 ( .Y(n4196), .A0(n4181), .A1(n4197) );
  nand02 U1921 ( .Y(n4198), .A0(n4176), .A1(n4177) );
  inv01 U1922 ( .Y(n4183), .A(n4198) );
  nand02 U1923 ( .Y(n4199), .A0(n4176), .A1(n4177) );
  inv01 U1924 ( .Y(n4185), .A(n4199) );
  nand02 U1925 ( .Y(n4200), .A0(n4176), .A1(n4178) );
  inv01 U1926 ( .Y(n4187), .A(n4200) );
  nand02 U1927 ( .Y(n4201), .A0(n4176), .A1(n4179) );
  inv01 U1928 ( .Y(n4189), .A(n4201) );
  nand02 U1929 ( .Y(n4202), .A0(n4177), .A1(n4178) );
  inv01 U1930 ( .Y(n4191), .A(n4202) );
  nand02 U1931 ( .Y(n4203), .A0(n4177), .A1(n4179) );
  inv01 U1932 ( .Y(n4193), .A(n4203) );
  nand02 U1933 ( .Y(n4204), .A0(n4178), .A1(n4180) );
  inv01 U1934 ( .Y(n4195), .A(n4204) );
  nand02 U1935 ( .Y(n4205), .A0(n4179), .A1(n4180) );
  inv01 U1936 ( .Y(n4197), .A(n4205) );
  nand02 U1937 ( .Y(n4206), .A0(n4182), .A1(n4184) );
  inv01 U1938 ( .Y(n4207), .A(n4206) );
  nand02 U1939 ( .Y(n4208), .A0(n4186), .A1(n4188) );
  inv01 U1940 ( .Y(n4209), .A(n4208) );
  nand02 U1941 ( .Y(n4210), .A0(n4207), .A1(n4209) );
  inv01 U1942 ( .Y(n4174), .A(n4210) );
  nand02 U1943 ( .Y(n4211), .A0(n4190), .A1(n4192) );
  inv01 U1944 ( .Y(n4212), .A(n4211) );
  nand02 U1945 ( .Y(n4213), .A0(n4194), .A1(n4196) );
  inv01 U1946 ( .Y(n4214), .A(n4213) );
  nand02 U1947 ( .Y(n4215), .A0(n4212), .A1(n4214) );
  inv01 U1948 ( .Y(n4175), .A(n4215) );
  inv02 U1949 ( .Y(n5395), .A(n4801) );
  nand02 U1950 ( .Y(n4216), .A0(n5293), .A1(n5148) );
  inv02 U1951 ( .Y(n4217), .A(n4216) );
  nand02 U1952 ( .Y(n5439), .A0(n4218), .A1(n4219) );
  inv02 U1953 ( .Y(n4220), .A(n5402) );
  inv02 U1954 ( .Y(n4221), .A(n5440) );
  inv02 U1955 ( .Y(n4222), .A(n5372) );
  inv02 U1956 ( .Y(n4223), .A(n5217) );
  inv02 U1957 ( .Y(n4224), .A(n5218) );
  inv02 U1958 ( .Y(n4225), .A(n5216) );
  nand02 U1959 ( .Y(n4226), .A0(n4222), .A1(n4227) );
  nand02 U1960 ( .Y(n4228), .A0(n4223), .A1(n4229) );
  nand02 U1961 ( .Y(n4230), .A0(n4224), .A1(n4231) );
  nand02 U1962 ( .Y(n4232), .A0(n4224), .A1(n4233) );
  nand02 U1963 ( .Y(n4234), .A0(n4225), .A1(n4235) );
  nand02 U1964 ( .Y(n4236), .A0(n4225), .A1(n4237) );
  nand02 U1965 ( .Y(n4238), .A0(n4225), .A1(n4239) );
  nand02 U1966 ( .Y(n4240), .A0(n4225), .A1(n4241) );
  nand02 U1967 ( .Y(n4242), .A0(n4220), .A1(n4221) );
  inv01 U1968 ( .Y(n4227), .A(n4242) );
  nand02 U1969 ( .Y(n4243), .A0(n4220), .A1(n4221) );
  inv01 U1970 ( .Y(n4229), .A(n4243) );
  nand02 U1971 ( .Y(n4244), .A0(n4220), .A1(n4222) );
  inv01 U1972 ( .Y(n4231), .A(n4244) );
  nand02 U1973 ( .Y(n4245), .A0(n4220), .A1(n4223) );
  inv01 U1974 ( .Y(n4233), .A(n4245) );
  nand02 U1975 ( .Y(n4246), .A0(n4221), .A1(n4222) );
  inv01 U1976 ( .Y(n4235), .A(n4246) );
  nand02 U1977 ( .Y(n4247), .A0(n4221), .A1(n4223) );
  inv01 U1978 ( .Y(n4237), .A(n4247) );
  nand02 U1979 ( .Y(n4248), .A0(n4222), .A1(n4224) );
  inv01 U1980 ( .Y(n4239), .A(n4248) );
  nand02 U1981 ( .Y(n4249), .A0(n4223), .A1(n4224) );
  inv01 U1982 ( .Y(n4241), .A(n4249) );
  nand02 U1983 ( .Y(n4250), .A0(n4226), .A1(n4228) );
  inv01 U1984 ( .Y(n4251), .A(n4250) );
  nand02 U1985 ( .Y(n4252), .A0(n4230), .A1(n4232) );
  inv01 U1986 ( .Y(n4253), .A(n4252) );
  nand02 U1987 ( .Y(n4254), .A0(n4251), .A1(n4253) );
  inv01 U1988 ( .Y(n4218), .A(n4254) );
  nand02 U1989 ( .Y(n4255), .A0(n4234), .A1(n4236) );
  inv01 U1990 ( .Y(n4256), .A(n4255) );
  nand02 U1991 ( .Y(n4257), .A0(n4238), .A1(n4240) );
  inv01 U1992 ( .Y(n4258), .A(n4257) );
  nand02 U1993 ( .Y(n4259), .A0(n4256), .A1(n4258) );
  inv01 U1994 ( .Y(n4219), .A(n4259) );
  nand02 U1995 ( .Y(n5458), .A0(n4260), .A1(n4261) );
  inv02 U1996 ( .Y(n4262), .A(n5432) );
  inv02 U1997 ( .Y(n4263), .A(n4816) );
  inv02 U1998 ( .Y(n4264), .A(n5394) );
  inv02 U1999 ( .Y(n4265), .A(n5217) );
  inv02 U2000 ( .Y(n4266), .A(n5434) );
  nand02 U2001 ( .Y(n4267), .A0(n4264), .A1(n4268) );
  nand02 U2002 ( .Y(n4269), .A0(n4265), .A1(n4270) );
  nand02 U2003 ( .Y(n4271), .A0(n4266), .A1(n4272) );
  nand02 U2004 ( .Y(n4273), .A0(n4266), .A1(n4274) );
  nand02 U2005 ( .Y(n4275), .A0(n4348), .A1(n4276) );
  nand02 U2006 ( .Y(n4277), .A0(n4390), .A1(n4278) );
  nand02 U2007 ( .Y(n4279), .A0(n4348), .A1(n4280) );
  nand02 U2008 ( .Y(n4281), .A0(n4390), .A1(n4282) );
  nand02 U2009 ( .Y(n4283), .A0(n4262), .A1(n4263) );
  inv01 U2010 ( .Y(n4268), .A(n4283) );
  nand02 U2011 ( .Y(n4284), .A0(n4262), .A1(n4263) );
  inv01 U2012 ( .Y(n4270), .A(n4284) );
  nand02 U2013 ( .Y(n4285), .A0(n4262), .A1(n4264) );
  inv01 U2014 ( .Y(n4272), .A(n4285) );
  nand02 U2015 ( .Y(n4286), .A0(n4262), .A1(n4265) );
  inv01 U2016 ( .Y(n4274), .A(n4286) );
  nand02 U2017 ( .Y(n4287), .A0(n4263), .A1(n4264) );
  inv01 U2018 ( .Y(n4276), .A(n4287) );
  nand02 U2019 ( .Y(n4288), .A0(n4263), .A1(n4265) );
  inv01 U2020 ( .Y(n4278), .A(n4288) );
  nand02 U2021 ( .Y(n4289), .A0(n4264), .A1(n4266) );
  inv01 U2022 ( .Y(n4280), .A(n4289) );
  nand02 U2023 ( .Y(n4290), .A0(n4265), .A1(n4266) );
  inv01 U2024 ( .Y(n4282), .A(n4290) );
  nand02 U2025 ( .Y(n4291), .A0(n4267), .A1(n4269) );
  inv01 U2026 ( .Y(n4292), .A(n4291) );
  nand02 U2027 ( .Y(n4293), .A0(n4271), .A1(n4273) );
  inv01 U2028 ( .Y(n4294), .A(n4293) );
  nand02 U2029 ( .Y(n4295), .A0(n4292), .A1(n4294) );
  inv01 U2030 ( .Y(n4260), .A(n4295) );
  nand02 U2031 ( .Y(n4296), .A0(n4275), .A1(n4277) );
  inv01 U2032 ( .Y(n4297), .A(n4296) );
  nand02 U2033 ( .Y(n4298), .A0(n4279), .A1(n4281) );
  inv01 U2034 ( .Y(n4299), .A(n4298) );
  nand02 U2035 ( .Y(n4300), .A0(n4297), .A1(n4299) );
  inv01 U2036 ( .Y(n4261), .A(n4300) );
  buf08 U2037 ( .Y(n5217), .A(n5363) );
  nand02 U2038 ( .Y(n5460), .A0(n4301), .A1(n4302) );
  inv02 U2039 ( .Y(n4303), .A(n5463) );
  inv02 U2040 ( .Y(n4304), .A(n5375) );
  inv02 U2041 ( .Y(n4305), .A(n5279) );
  inv02 U2042 ( .Y(n4306), .A(n____return2686) );
  inv02 U2043 ( .Y(n4307), .A(n5217) );
  inv02 U2044 ( .Y(n4308), .A(n5197) );
  nand02 U2045 ( .Y(n4309), .A0(n4305), .A1(n4310) );
  nand02 U2046 ( .Y(n4311), .A0(n4306), .A1(n4312) );
  nand02 U2047 ( .Y(n4313), .A0(n4307), .A1(n4314) );
  nand02 U2048 ( .Y(n4315), .A0(n4307), .A1(n4316) );
  nand02 U2049 ( .Y(n4317), .A0(n4308), .A1(n4318) );
  nand02 U2050 ( .Y(n4319), .A0(n4308), .A1(n4320) );
  nand02 U2051 ( .Y(n4321), .A0(n4308), .A1(n4322) );
  nand02 U2052 ( .Y(n4323), .A0(n4308), .A1(n4324) );
  nand02 U2053 ( .Y(n4325), .A0(n4303), .A1(n4304) );
  inv01 U2054 ( .Y(n4310), .A(n4325) );
  nand02 U2055 ( .Y(n4326), .A0(n4303), .A1(n4304) );
  inv01 U2056 ( .Y(n4312), .A(n4326) );
  nand02 U2057 ( .Y(n4327), .A0(n4303), .A1(n4305) );
  inv01 U2058 ( .Y(n4314), .A(n4327) );
  nand02 U2059 ( .Y(n4328), .A0(n4303), .A1(n4306) );
  inv01 U2060 ( .Y(n4316), .A(n4328) );
  nand02 U2061 ( .Y(n4329), .A0(n4304), .A1(n4305) );
  inv01 U2062 ( .Y(n4318), .A(n4329) );
  nand02 U2063 ( .Y(n4330), .A0(n4304), .A1(n4306) );
  inv01 U2064 ( .Y(n4320), .A(n4330) );
  nand02 U2065 ( .Y(n4331), .A0(n4305), .A1(n4307) );
  inv01 U2066 ( .Y(n4322), .A(n4331) );
  nand02 U2067 ( .Y(n4332), .A0(n4306), .A1(n4307) );
  inv01 U2068 ( .Y(n4324), .A(n4332) );
  nand02 U2069 ( .Y(n4333), .A0(n4309), .A1(n4311) );
  inv01 U2070 ( .Y(n4334), .A(n4333) );
  nand02 U2071 ( .Y(n4335), .A0(n4313), .A1(n4315) );
  inv01 U2072 ( .Y(n4336), .A(n4335) );
  nand02 U2073 ( .Y(n4337), .A0(n4334), .A1(n4336) );
  inv01 U2074 ( .Y(n4301), .A(n4337) );
  nand02 U2075 ( .Y(n4338), .A0(n4317), .A1(n4319) );
  inv01 U2076 ( .Y(n4339), .A(n4338) );
  nand02 U2077 ( .Y(n4340), .A0(n4321), .A1(n4323) );
  inv01 U2078 ( .Y(n4341), .A(n4340) );
  nand02 U2079 ( .Y(n4342), .A0(n4339), .A1(n4341) );
  inv01 U2080 ( .Y(n4302), .A(n4342) );
  nand02 U2081 ( .Y(n5377), .A0(n4343), .A1(n4344) );
  inv02 U2082 ( .Y(n4345), .A(n5380) );
  inv02 U2083 ( .Y(n4346), .A(n5379) );
  inv02 U2084 ( .Y(n4347), .A(n5378) );
  inv02 U2085 ( .Y(n4348), .A(n5365) );
  inv02 U2086 ( .Y(n4349), .A(n5370) );
  inv02 U2087 ( .Y(n4350), .A(n5216) );
  nand02 U2088 ( .Y(n4351), .A0(n4347), .A1(n4352) );
  nand02 U2089 ( .Y(n4353), .A0(n4348), .A1(n4354) );
  nand02 U2090 ( .Y(n4355), .A0(n4349), .A1(n4356) );
  nand02 U2091 ( .Y(n4357), .A0(n4349), .A1(n4358) );
  nand02 U2092 ( .Y(n4359), .A0(n4350), .A1(n4360) );
  nand02 U2093 ( .Y(n4361), .A0(n4350), .A1(n4362) );
  nand02 U2094 ( .Y(n4363), .A0(n4350), .A1(n4364) );
  nand02 U2095 ( .Y(n4365), .A0(n4350), .A1(n4366) );
  nand02 U2096 ( .Y(n4367), .A0(n4345), .A1(n4346) );
  inv01 U2097 ( .Y(n4352), .A(n4367) );
  nand02 U2098 ( .Y(n4368), .A0(n4345), .A1(n4346) );
  inv01 U2099 ( .Y(n4354), .A(n4368) );
  nand02 U2100 ( .Y(n4369), .A0(n4345), .A1(n4347) );
  inv01 U2101 ( .Y(n4356), .A(n4369) );
  nand02 U2102 ( .Y(n4370), .A0(n4345), .A1(n4348) );
  inv01 U2103 ( .Y(n4358), .A(n4370) );
  nand02 U2104 ( .Y(n4371), .A0(n4346), .A1(n4347) );
  inv01 U2105 ( .Y(n4360), .A(n4371) );
  nand02 U2106 ( .Y(n4372), .A0(n4346), .A1(n4348) );
  inv01 U2107 ( .Y(n4362), .A(n4372) );
  nand02 U2108 ( .Y(n4373), .A0(n4347), .A1(n4349) );
  inv01 U2109 ( .Y(n4364), .A(n4373) );
  nand02 U2110 ( .Y(n4374), .A0(n4348), .A1(n4349) );
  inv01 U2111 ( .Y(n4366), .A(n4374) );
  nand02 U2112 ( .Y(n4375), .A0(n4351), .A1(n4353) );
  inv01 U2113 ( .Y(n4376), .A(n4375) );
  nand02 U2114 ( .Y(n4377), .A0(n4355), .A1(n4357) );
  inv01 U2115 ( .Y(n4378), .A(n4377) );
  nand02 U2116 ( .Y(n4379), .A0(n4376), .A1(n4378) );
  inv01 U2117 ( .Y(n4343), .A(n4379) );
  nand02 U2118 ( .Y(n4380), .A0(n4359), .A1(n4361) );
  inv01 U2119 ( .Y(n4381), .A(n4380) );
  nand02 U2120 ( .Y(n4382), .A0(n4363), .A1(n4365) );
  inv01 U2121 ( .Y(n4383), .A(n4382) );
  nand02 U2122 ( .Y(n4384), .A0(n4381), .A1(n4383) );
  inv01 U2123 ( .Y(n4344), .A(n4384) );
  nand02 U2124 ( .Y(n5393), .A0(n4385), .A1(n4386) );
  inv02 U2125 ( .Y(n4387), .A(n5197) );
  inv02 U2126 ( .Y(n4388), .A(n5395) );
  inv02 U2127 ( .Y(n4389), .A(n5394) );
  inv02 U2128 ( .Y(n4390), .A(n5365) );
  inv02 U2129 ( .Y(n4391), .A(n5218) );
  nand02 U2130 ( .Y(n4392), .A0(n4389), .A1(n4393) );
  nand02 U2131 ( .Y(n4394), .A0(n4390), .A1(n4395) );
  nand02 U2132 ( .Y(n4396), .A0(n4391), .A1(n4397) );
  nand02 U2133 ( .Y(n4398), .A0(n4391), .A1(n4399) );
  nand02 U2134 ( .Y(n4400), .A0(n5340), .A1(n4401) );
  nand02 U2135 ( .Y(n4402), .A0(n5340), .A1(n4403) );
  nand02 U2136 ( .Y(n4404), .A0(n5340), .A1(n4405) );
  nand02 U2137 ( .Y(n4406), .A0(n5340), .A1(n4407) );
  nand02 U2138 ( .Y(n4408), .A0(n4387), .A1(n4388) );
  inv01 U2139 ( .Y(n4393), .A(n4408) );
  nand02 U2140 ( .Y(n4409), .A0(n4387), .A1(n4388) );
  inv01 U2141 ( .Y(n4395), .A(n4409) );
  nand02 U2142 ( .Y(n4410), .A0(n4387), .A1(n4389) );
  inv01 U2143 ( .Y(n4397), .A(n4410) );
  nand02 U2144 ( .Y(n4411), .A0(n4387), .A1(n4390) );
  inv01 U2145 ( .Y(n4399), .A(n4411) );
  nand02 U2146 ( .Y(n4412), .A0(n4388), .A1(n4389) );
  inv01 U2147 ( .Y(n4401), .A(n4412) );
  nand02 U2148 ( .Y(n4413), .A0(n4388), .A1(n4390) );
  inv01 U2149 ( .Y(n4403), .A(n4413) );
  nand02 U2150 ( .Y(n4414), .A0(n4389), .A1(n4391) );
  inv01 U2151 ( .Y(n4405), .A(n4414) );
  nand02 U2152 ( .Y(n4415), .A0(n4390), .A1(n4391) );
  inv01 U2153 ( .Y(n4407), .A(n4415) );
  nand02 U2154 ( .Y(n4416), .A0(n4392), .A1(n4394) );
  inv01 U2155 ( .Y(n4417), .A(n4416) );
  nand02 U2156 ( .Y(n4418), .A0(n4396), .A1(n4398) );
  inv01 U2157 ( .Y(n4419), .A(n4418) );
  nand02 U2158 ( .Y(n4420), .A0(n4417), .A1(n4419) );
  inv01 U2159 ( .Y(n4385), .A(n4420) );
  nand02 U2160 ( .Y(n4421), .A0(n4400), .A1(n4402) );
  inv01 U2161 ( .Y(n4422), .A(n4421) );
  nand02 U2162 ( .Y(n4423), .A0(n4404), .A1(n4406) );
  inv01 U2163 ( .Y(n4424), .A(n4423) );
  nand02 U2164 ( .Y(n4425), .A0(n4422), .A1(n4424) );
  inv01 U2165 ( .Y(n4386), .A(n4425) );
  inv01 U2166 ( .Y(n5400), .A(n4426) );
  nor02 U2167 ( .Y(n4427), .A0(n5402), .A1(n4428) );
  nor02 U2168 ( .Y(n4429), .A0(n5402), .A1(n4430) );
  nor02 U2169 ( .Y(n4431), .A0(n5402), .A1(n4432) );
  nor02 U2170 ( .Y(n4433), .A0(n5402), .A1(n4434) );
  nor02 U2171 ( .Y(n4435), .A0(n5218), .A1(n4436) );
  nor02 U2172 ( .Y(n4437), .A0(n5218), .A1(n4438) );
  nor02 U2173 ( .Y(n4439), .A0(n5218), .A1(n4440) );
  nor02 U2174 ( .Y(n4441), .A0(n5218), .A1(n4442) );
  nor02 U2175 ( .Y(n4426), .A0(n4443), .A1(n4444) );
  nor02 U2176 ( .Y(n4445), .A0(n5372), .A1(n5401) );
  inv01 U2177 ( .Y(n4428), .A(n4445) );
  nor02 U2178 ( .Y(n4446), .A0(n5216), .A1(n5401) );
  inv01 U2179 ( .Y(n4430), .A(n4446) );
  nor02 U2180 ( .Y(n4447), .A0(n5372), .A1(n5197) );
  inv01 U2181 ( .Y(n4432), .A(n4447) );
  nor02 U2182 ( .Y(n4448), .A0(n5216), .A1(n5197) );
  inv01 U2183 ( .Y(n4434), .A(n4448) );
  nor02 U2184 ( .Y(n4449), .A0(n5372), .A1(n5401) );
  inv01 U2185 ( .Y(n4436), .A(n4449) );
  nor02 U2186 ( .Y(n4450), .A0(n5216), .A1(n5401) );
  inv01 U2187 ( .Y(n4438), .A(n4450) );
  nor02 U2188 ( .Y(n4451), .A0(n5372), .A1(n5197) );
  inv01 U2189 ( .Y(n4440), .A(n4451) );
  nor02 U2190 ( .Y(n4452), .A0(n5216), .A1(n5197) );
  inv01 U2191 ( .Y(n4442), .A(n4452) );
  nor02 U2192 ( .Y(n4453), .A0(n4427), .A1(n4429) );
  inv01 U2193 ( .Y(n4454), .A(n4453) );
  nor02 U2194 ( .Y(n4455), .A0(n4431), .A1(n4433) );
  inv01 U2195 ( .Y(n4456), .A(n4455) );
  nor02 U2196 ( .Y(n4457), .A0(n4454), .A1(n4456) );
  inv01 U2197 ( .Y(n4443), .A(n4457) );
  nor02 U2198 ( .Y(n4458), .A0(n4435), .A1(n4437) );
  inv01 U2199 ( .Y(n4459), .A(n4458) );
  nor02 U2200 ( .Y(n4460), .A0(n4439), .A1(n4441) );
  inv01 U2201 ( .Y(n4461), .A(n4460) );
  nor02 U2202 ( .Y(n4462), .A0(n4459), .A1(n4461) );
  inv01 U2203 ( .Y(n4444), .A(n4462) );
  buf08 U2204 ( .Y(n5216), .A(n5368) );
  inv02 U2205 ( .Y(n5401), .A(n4860) );
  inv02 U2206 ( .Y(n5402), .A(n4795) );
  inv08 U2207 ( .Y(n4463), .A(n5488) );
  inv01 U2208 ( .Y(n5481), .A(n4465) );
  inv01 U2209 ( .Y(n4466), .A(opb_i[23]) );
  inv01 U2210 ( .Y(n4467), .A(opb_i[24]) );
  inv01 U2211 ( .Y(n4468), .A(opb_i[25]) );
  inv01 U2212 ( .Y(n4469), .A(opb_i[26]) );
  nand02 U2213 ( .Y(n4465), .A0(n4470), .A1(n4471) );
  nand02 U2214 ( .Y(n4472), .A0(n4466), .A1(n4467) );
  inv01 U2215 ( .Y(n4470), .A(n4472) );
  nand02 U2216 ( .Y(n4473), .A0(n4468), .A1(n4469) );
  inv01 U2217 ( .Y(n4471), .A(n4473) );
  inv02 U2218 ( .Y(n5289), .A(n4474) );
  nand02 U2219 ( .Y(n4474), .A0(n5298), .A1(n4475) );
  nand02 U2220 ( .Y(n4476), .A0(n5184), .A1(n5196) );
  inv01 U2221 ( .Y(n4475), .A(n4476) );
  inv01 U2222 ( .Y(n5482), .A(n4477) );
  inv01 U2223 ( .Y(n4478), .A(opb_i[27]) );
  inv01 U2224 ( .Y(n4479), .A(opb_i[28]) );
  inv01 U2225 ( .Y(n4480), .A(opb_i[29]) );
  inv01 U2226 ( .Y(n4481), .A(opb_i[30]) );
  nand02 U2227 ( .Y(n4477), .A0(n4482), .A1(n4483) );
  nand02 U2228 ( .Y(n4484), .A0(n4478), .A1(n4479) );
  inv01 U2229 ( .Y(n4482), .A(n4484) );
  nand02 U2230 ( .Y(n4485), .A0(n4480), .A1(n4481) );
  inv01 U2231 ( .Y(n4483), .A(n4485) );
  nand02 U2232 ( .Y(n5461), .A0(n4486), .A1(n4487) );
  inv02 U2233 ( .Y(n4488), .A(n5407) );
  inv02 U2234 ( .Y(n4489), .A(n5380) );
  inv02 U2235 ( .Y(n4490), .A(n5218) );
  inv02 U2236 ( .Y(n4491), .A(n5278) );
  inv02 U2237 ( .Y(n4492), .A(n5419) );
  inv02 U2238 ( .Y(n4493), .A(n5365) );
  inv02 U2239 ( .Y(n4494), .A(n5216) );
  nand02 U2240 ( .Y(n4495), .A0(n4490), .A1(n4496) );
  nand02 U2241 ( .Y(n4497), .A0(n4491), .A1(n4498) );
  nand02 U2242 ( .Y(n4499), .A0(n4492), .A1(n4500) );
  nand02 U2243 ( .Y(n4501), .A0(n4493), .A1(n4502) );
  nand02 U2244 ( .Y(n4503), .A0(n4493), .A1(n4504) );
  nand02 U2245 ( .Y(n4505), .A0(n4493), .A1(n4506) );
  nand02 U2246 ( .Y(n4507), .A0(n4494), .A1(n4508) );
  nand02 U2247 ( .Y(n4509), .A0(n4494), .A1(n4510) );
  nand02 U2248 ( .Y(n4511), .A0(n4494), .A1(n4512) );
  nand02 U2249 ( .Y(n4513), .A0(n4494), .A1(n4514) );
  nand02 U2250 ( .Y(n4515), .A0(n4494), .A1(n4516) );
  nand02 U2251 ( .Y(n4517), .A0(n4494), .A1(n4518) );
  nand02 U2252 ( .Y(n4519), .A0(n4488), .A1(n4489) );
  inv01 U2253 ( .Y(n4496), .A(n4519) );
  nand02 U2254 ( .Y(n4520), .A0(n4488), .A1(n4489) );
  inv01 U2255 ( .Y(n4498), .A(n4520) );
  nand02 U2256 ( .Y(n4521), .A0(n4488), .A1(n4489) );
  inv01 U2257 ( .Y(n4500), .A(n4521) );
  nand02 U2258 ( .Y(n4522), .A0(n4488), .A1(n4490) );
  inv01 U2259 ( .Y(n4502), .A(n4522) );
  nand02 U2260 ( .Y(n4523), .A0(n4488), .A1(n4491) );
  inv01 U2261 ( .Y(n4504), .A(n4523) );
  nand02 U2262 ( .Y(n4524), .A0(n4488), .A1(n4492) );
  inv01 U2263 ( .Y(n4506), .A(n4524) );
  nand02 U2264 ( .Y(n4525), .A0(n4489), .A1(n4490) );
  inv01 U2265 ( .Y(n4508), .A(n4525) );
  nand02 U2266 ( .Y(n4526), .A0(n4489), .A1(n4491) );
  inv01 U2267 ( .Y(n4510), .A(n4526) );
  nand02 U2268 ( .Y(n4527), .A0(n4489), .A1(n4492) );
  inv01 U2269 ( .Y(n4512), .A(n4527) );
  nand02 U2270 ( .Y(n4528), .A0(n4490), .A1(n4493) );
  inv01 U2271 ( .Y(n4514), .A(n4528) );
  nand02 U2272 ( .Y(n4529), .A0(n4491), .A1(n4493) );
  inv01 U2273 ( .Y(n4516), .A(n4529) );
  nand02 U2274 ( .Y(n4530), .A0(n4492), .A1(n4493) );
  inv01 U2275 ( .Y(n4518), .A(n4530) );
  nand02 U2276 ( .Y(n4531), .A0(n4495), .A1(n4497) );
  inv01 U2277 ( .Y(n4532), .A(n4531) );
  nand02 U2278 ( .Y(n4533), .A0(n4499), .A1(n4532) );
  inv01 U2279 ( .Y(n4534), .A(n4533) );
  nand02 U2280 ( .Y(n4535), .A0(n4501), .A1(n4503) );
  inv01 U2281 ( .Y(n4536), .A(n4535) );
  nand02 U2282 ( .Y(n4537), .A0(n4505), .A1(n4536) );
  inv01 U2283 ( .Y(n4538), .A(n4537) );
  nand02 U2284 ( .Y(n4539), .A0(n4534), .A1(n4538) );
  inv01 U2285 ( .Y(n4486), .A(n4539) );
  nand02 U2286 ( .Y(n4540), .A0(n4507), .A1(n4509) );
  inv01 U2287 ( .Y(n4541), .A(n4540) );
  nand02 U2288 ( .Y(n4542), .A0(n4511), .A1(n4541) );
  inv01 U2289 ( .Y(n4543), .A(n4542) );
  nand02 U2290 ( .Y(n4544), .A0(n4513), .A1(n4515) );
  inv01 U2291 ( .Y(n4545), .A(n4544) );
  nand02 U2292 ( .Y(n4546), .A0(n4517), .A1(n4545) );
  inv01 U2293 ( .Y(n4547), .A(n4546) );
  nand02 U2294 ( .Y(n4548), .A0(n4543), .A1(n4547) );
  inv01 U2295 ( .Y(n4487), .A(n4548) );
  buf08 U2296 ( .Y(n5218), .A(n5338) );
  nand02 U2297 ( .Y(n5411), .A0(n4549), .A1(n4550) );
  inv02 U2298 ( .Y(n4551), .A(n5412) );
  inv02 U2299 ( .Y(n4552), .A(n5019) );
  inv01 U2300 ( .Y(n4553), .A(s_exp_diff_2_) );
  inv01 U2301 ( .Y(n4554), .A(n5382) );
  inv01 U2302 ( .Y(n4555), .A(s_exp_diff_3_) );
  inv01 U2303 ( .Y(n4556), .A(n5386) );
  nand02 U2304 ( .Y(n4557), .A0(n4553), .A1(n4558) );
  nand02 U2305 ( .Y(n4559), .A0(n4554), .A1(n4560) );
  nand02 U2306 ( .Y(n4561), .A0(n4555), .A1(n4562) );
  nand02 U2307 ( .Y(n4563), .A0(n4556), .A1(n4564) );
  nand02 U2308 ( .Y(n4565), .A0(n4556), .A1(n4566) );
  nand02 U2309 ( .Y(n4567), .A0(n4556), .A1(n4568) );
  nand02 U2310 ( .Y(n4569), .A0(n4551), .A1(n4552) );
  inv01 U2311 ( .Y(n4558), .A(n4569) );
  nand02 U2312 ( .Y(n4570), .A0(n4551), .A1(n4552) );
  inv01 U2313 ( .Y(n4560), .A(n4570) );
  nand02 U2314 ( .Y(n4571), .A0(n4551), .A1(n4552) );
  inv01 U2315 ( .Y(n4562), .A(n4571) );
  nand02 U2316 ( .Y(n4572), .A0(n4551), .A1(n4553) );
  inv01 U2317 ( .Y(n4564), .A(n4572) );
  nand02 U2318 ( .Y(n4573), .A0(n4551), .A1(n4554) );
  inv01 U2319 ( .Y(n4566), .A(n4573) );
  nand02 U2320 ( .Y(n4574), .A0(n4551), .A1(n4555) );
  inv01 U2321 ( .Y(n4568), .A(n4574) );
  nand02 U2322 ( .Y(n4575), .A0(n4557), .A1(n4559) );
  inv01 U2323 ( .Y(n4576), .A(n4575) );
  nand02 U2324 ( .Y(n4577), .A0(n4561), .A1(n4576) );
  inv01 U2325 ( .Y(n4549), .A(n4577) );
  nand02 U2326 ( .Y(n4578), .A0(n4563), .A1(n4565) );
  inv01 U2327 ( .Y(n4579), .A(n4578) );
  nand02 U2328 ( .Y(n4580), .A0(n4567), .A1(n4579) );
  inv01 U2329 ( .Y(n4550), .A(n4580) );
  inv01 U2330 ( .Y(n5484), .A(n4581) );
  inv01 U2331 ( .Y(n4582), .A(opa_i[27]) );
  inv01 U2332 ( .Y(n4583), .A(opa_i[28]) );
  inv01 U2333 ( .Y(n4584), .A(opa_i[29]) );
  inv01 U2334 ( .Y(n4585), .A(opa_i[30]) );
  nand02 U2335 ( .Y(n4581), .A0(n4586), .A1(n4587) );
  nand02 U2336 ( .Y(n4588), .A0(n4582), .A1(n4583) );
  inv01 U2337 ( .Y(n4586), .A(n4588) );
  nand02 U2338 ( .Y(n4589), .A0(n4584), .A1(n4585) );
  inv01 U2339 ( .Y(n4587), .A(n4589) );
  nor02 U2340 ( .Y(n5301), .A0(n4590), .A1(n4591) );
  nor02 U2341 ( .Y(n4592), .A0(n5302), .A1(n5233) );
  inv02 U2342 ( .Y(n4590), .A(n4592) );
  nor02 U2343 ( .Y(n4593), .A0(n5234), .A1(n5231) );
  inv01 U2344 ( .Y(n4591), .A(n4593) );
  inv01 U2345 ( .Y(n5483), .A(n4594) );
  inv01 U2346 ( .Y(n4595), .A(opa_i[23]) );
  inv01 U2347 ( .Y(n4596), .A(opa_i[24]) );
  inv01 U2348 ( .Y(n4597), .A(opa_i[25]) );
  inv01 U2349 ( .Y(n4598), .A(opa_i[26]) );
  nand02 U2350 ( .Y(n4594), .A0(n4599), .A1(n4600) );
  nand02 U2351 ( .Y(n4601), .A0(n4595), .A1(n4596) );
  inv01 U2352 ( .Y(n4599), .A(n4601) );
  nand02 U2353 ( .Y(n4602), .A0(n4597), .A1(n4598) );
  inv01 U2354 ( .Y(n4600), .A(n4602) );
  inv02 U2355 ( .Y(U403_U5_Z_1), .A(n4603) );
  nor02 U2356 ( .Y(n4604), .A0(n____return128), .A1(n4915) );
  nor02 U2357 ( .Y(n4605), .A0(n5223), .A1(n4931) );
  nor02 U2358 ( .Y(n4603), .A0(n4604), .A1(n4605) );
  inv02 U2359 ( .Y(U403_U5_Z_2), .A(n4606) );
  nor02 U2360 ( .Y(n4607), .A0(n____return128), .A1(n4921) );
  nor02 U2361 ( .Y(n4608), .A0(n5222), .A1(n4939) );
  nor02 U2362 ( .Y(n4606), .A0(n4607), .A1(n4608) );
  inv02 U2363 ( .Y(U403_U5_Z_7), .A(n4609) );
  nor02 U2364 ( .Y(n4610), .A0(n____return128), .A1(n4924) );
  nor02 U2365 ( .Y(n4611), .A0(n5223), .A1(n4943) );
  nor02 U2366 ( .Y(n4609), .A0(n4610), .A1(n4611) );
  inv02 U2367 ( .Y(U403_U5_Z_6), .A(n4612) );
  nor02 U2368 ( .Y(n4613), .A0(n____return128), .A1(n4909) );
  nor02 U2369 ( .Y(n4614), .A0(n5222), .A1(n4937) );
  nor02 U2370 ( .Y(n4612), .A0(n4613), .A1(n4614) );
  inv02 U2371 ( .Y(U403_U5_Z_4), .A(n4615) );
  nor02 U2372 ( .Y(n4616), .A0(n____return128), .A1(n4927) );
  nor02 U2373 ( .Y(n4617), .A0(n5222), .A1(n4941) );
  nor02 U2374 ( .Y(n4615), .A0(n4616), .A1(n4617) );
  inv02 U2375 ( .Y(U403_U5_Z_3), .A(n4618) );
  nor02 U2376 ( .Y(n4619), .A0(n____return128), .A1(n4912) );
  nor02 U2377 ( .Y(n4620), .A0(n5223), .A1(n4935) );
  nor02 U2378 ( .Y(n4618), .A0(n4619), .A1(n4620) );
  inv02 U2379 ( .Y(U403_U5_Z_5), .A(n4621) );
  nor02 U2380 ( .Y(n4622), .A0(n____return128), .A1(n4918) );
  nor02 U2381 ( .Y(n4623), .A0(n5223), .A1(n4933) );
  nor02 U2382 ( .Y(n4621), .A0(n4622), .A1(n4623) );
  inv02 U2383 ( .Y(U403_U5_Z_0), .A(n4624) );
  nor02 U2384 ( .Y(n4625), .A0(n____return128), .A1(n5469) );
  nor02 U2385 ( .Y(n4626), .A0(n5223), .A1(n4957) );
  nor02 U2386 ( .Y(n4624), .A0(n4625), .A1(n4626) );
  nand02 U2387 ( .Y(n5319), .A0(n4627), .A1(n4628) );
  inv02 U2388 ( .Y(n4629), .A(n5376) );
  inv01 U2389 ( .Y(n4630), .A(n5218) );
  inv01 U2390 ( .Y(n4631), .A(n5217) );
  inv01 U2391 ( .Y(n4632), .A(n5374) );
  inv01 U2392 ( .Y(n4633), .A(n5375) );
  nand02 U2393 ( .Y(n4634), .A0(n4631), .A1(n4635) );
  nand02 U2394 ( .Y(n4636), .A0(n4632), .A1(n4637) );
  nand02 U2395 ( .Y(n4638), .A0(n4633), .A1(n4639) );
  nand02 U2396 ( .Y(n4640), .A0(n4633), .A1(n4641) );
  nand02 U2397 ( .Y(n4642), .A0(n4629), .A1(n4630) );
  inv01 U2398 ( .Y(n4635), .A(n4642) );
  nand02 U2399 ( .Y(n4643), .A0(n4629), .A1(n4630) );
  inv01 U2400 ( .Y(n4637), .A(n4643) );
  nand02 U2401 ( .Y(n4644), .A0(n4629), .A1(n4631) );
  inv01 U2402 ( .Y(n4639), .A(n4644) );
  nand02 U2403 ( .Y(n4645), .A0(n4629), .A1(n4632) );
  inv01 U2404 ( .Y(n4641), .A(n4645) );
  nand02 U2405 ( .Y(n4646), .A0(n4634), .A1(n4636) );
  inv01 U2406 ( .Y(n4627), .A(n4646) );
  nand02 U2407 ( .Y(n4647), .A0(n4638), .A1(n4640) );
  inv01 U2408 ( .Y(n4628), .A(n4647) );
  nand02 U2409 ( .Y(n5323), .A0(n4648), .A1(n4649) );
  inv02 U2410 ( .Y(n4650), .A(n5399) );
  inv01 U2411 ( .Y(n4651), .A(n5365) );
  inv01 U2412 ( .Y(n4652), .A(n5217) );
  inv01 U2413 ( .Y(n4653), .A(n5369) );
  inv01 U2414 ( .Y(n4654), .A(n5362) );
  nand02 U2415 ( .Y(n4655), .A0(n4652), .A1(n4656) );
  nand02 U2416 ( .Y(n4657), .A0(n4653), .A1(n4658) );
  nand02 U2417 ( .Y(n4659), .A0(n4654), .A1(n4660) );
  nand02 U2418 ( .Y(n4661), .A0(n4654), .A1(n4662) );
  nand02 U2419 ( .Y(n4663), .A0(n4650), .A1(n4651) );
  inv01 U2420 ( .Y(n4656), .A(n4663) );
  nand02 U2421 ( .Y(n4664), .A0(n4650), .A1(n4651) );
  inv01 U2422 ( .Y(n4658), .A(n4664) );
  nand02 U2423 ( .Y(n4665), .A0(n4650), .A1(n4652) );
  inv01 U2424 ( .Y(n4660), .A(n4665) );
  nand02 U2425 ( .Y(n4666), .A0(n4650), .A1(n4653) );
  inv01 U2426 ( .Y(n4662), .A(n4666) );
  nand02 U2427 ( .Y(n4667), .A0(n4655), .A1(n4657) );
  inv01 U2428 ( .Y(n4648), .A(n4667) );
  nand02 U2429 ( .Y(n4668), .A0(n4659), .A1(n4661) );
  inv01 U2430 ( .Y(n4649), .A(n4668) );
  nand02 U2431 ( .Y(n5325), .A0(n4669), .A1(n4670) );
  inv02 U2432 ( .Y(n4671), .A(n5404) );
  inv01 U2433 ( .Y(n4672), .A(n5365) );
  inv01 U2434 ( .Y(n4673), .A(n5217) );
  inv01 U2435 ( .Y(n4674), .A(n5380) );
  inv01 U2436 ( .Y(n4675), .A(n5374) );
  nand02 U2437 ( .Y(n4676), .A0(n4673), .A1(n4677) );
  nand02 U2438 ( .Y(n4678), .A0(n4674), .A1(n4679) );
  nand02 U2439 ( .Y(n4680), .A0(n4675), .A1(n4681) );
  nand02 U2440 ( .Y(n4682), .A0(n4675), .A1(n4683) );
  nand02 U2441 ( .Y(n4684), .A0(n4671), .A1(n4672) );
  inv01 U2442 ( .Y(n4677), .A(n4684) );
  nand02 U2443 ( .Y(n4685), .A0(n4671), .A1(n4672) );
  inv01 U2444 ( .Y(n4679), .A(n4685) );
  nand02 U2445 ( .Y(n4686), .A0(n4671), .A1(n4673) );
  inv01 U2446 ( .Y(n4681), .A(n4686) );
  nand02 U2447 ( .Y(n4687), .A0(n4671), .A1(n4674) );
  inv01 U2448 ( .Y(n4683), .A(n4687) );
  nand02 U2449 ( .Y(n4688), .A0(n4676), .A1(n4678) );
  inv01 U2450 ( .Y(n4669), .A(n4688) );
  nand02 U2451 ( .Y(n4689), .A0(n4680), .A1(n4682) );
  inv01 U2452 ( .Y(n4670), .A(n4689) );
  nand02 U2453 ( .Y(n5317), .A0(n4690), .A1(n4691) );
  inv02 U2454 ( .Y(n4692), .A(n5366) );
  inv01 U2455 ( .Y(n4693), .A(n5365) );
  inv01 U2456 ( .Y(n4694), .A(n5217) );
  inv01 U2457 ( .Y(n4695), .A(n5362) );
  inv01 U2458 ( .Y(n4696), .A(n5364) );
  nand02 U2459 ( .Y(n4697), .A0(n4694), .A1(n4698) );
  nand02 U2460 ( .Y(n4699), .A0(n4695), .A1(n4700) );
  nand02 U2461 ( .Y(n4701), .A0(n4696), .A1(n4702) );
  nand02 U2462 ( .Y(n4703), .A0(n4696), .A1(n4704) );
  nand02 U2463 ( .Y(n4705), .A0(n4692), .A1(n4693) );
  inv01 U2464 ( .Y(n4698), .A(n4705) );
  nand02 U2465 ( .Y(n4706), .A0(n4692), .A1(n4693) );
  inv01 U2466 ( .Y(n4700), .A(n4706) );
  nand02 U2467 ( .Y(n4707), .A0(n4692), .A1(n4694) );
  inv01 U2468 ( .Y(n4702), .A(n4707) );
  nand02 U2469 ( .Y(n4708), .A0(n4692), .A1(n4695) );
  inv01 U2470 ( .Y(n4704), .A(n4708) );
  nand02 U2471 ( .Y(n4709), .A0(n4697), .A1(n4699) );
  inv01 U2472 ( .Y(n4690), .A(n4709) );
  nand02 U2473 ( .Y(n4710), .A0(n4701), .A1(n4703) );
  inv01 U2474 ( .Y(n4691), .A(n4710) );
  nand02 U2475 ( .Y(n5358), .A0(n4711), .A1(n4712) );
  inv02 U2476 ( .Y(n4713), .A(n5454) );
  inv01 U2477 ( .Y(n4714), .A(n5365) );
  inv01 U2478 ( .Y(n4715), .A(n5217) );
  inv01 U2479 ( .Y(n4716), .A(n5383) );
  inv01 U2480 ( .Y(n4717), .A(n5387) );
  nand02 U2481 ( .Y(n4718), .A0(n4715), .A1(n4719) );
  nand02 U2482 ( .Y(n4720), .A0(n4716), .A1(n4721) );
  nand02 U2483 ( .Y(n4722), .A0(n4717), .A1(n4723) );
  nand02 U2484 ( .Y(n4724), .A0(n4717), .A1(n4725) );
  nand02 U2485 ( .Y(n4726), .A0(n4713), .A1(n4714) );
  inv01 U2486 ( .Y(n4719), .A(n4726) );
  nand02 U2487 ( .Y(n4727), .A0(n4713), .A1(n4714) );
  inv01 U2488 ( .Y(n4721), .A(n4727) );
  nand02 U2489 ( .Y(n4728), .A0(n4713), .A1(n4715) );
  inv01 U2490 ( .Y(n4723), .A(n4728) );
  nand02 U2491 ( .Y(n4729), .A0(n4713), .A1(n4716) );
  inv01 U2492 ( .Y(n4725), .A(n4729) );
  nand02 U2493 ( .Y(n4730), .A0(n4718), .A1(n4720) );
  inv01 U2494 ( .Y(n4711), .A(n4730) );
  nand02 U2495 ( .Y(n4731), .A0(n4722), .A1(n4724) );
  inv01 U2496 ( .Y(n4712), .A(n4731) );
  ao221 U2497 ( .Y(n4732), .A0(n5382), .A1(n5217), .B0(n5383), .B1(n5365), 
        .C0(n5384) );
  inv01 U2498 ( .Y(n4733), .A(n4732) );
  ao221 U2499 ( .Y(n4734), .A0(n5390), .A1(n5218), .B0(n5391), .B1(n5216), 
        .C0(n5457) );
  inv01 U2500 ( .Y(n4735), .A(n4734) );
  ao221 U2501 ( .Y(n4736), .A0(n5432), .A1(n5217), .B0(n5365), .B1(n5434), 
        .C0(n5447) );
  inv01 U2502 ( .Y(n4737), .A(n4736) );
  ao221 U2503 ( .Y(n4738), .A0(n5364), .A1(n5217), .B0(n5371), .B1(n5365), 
        .C0(n5449) );
  inv01 U2504 ( .Y(n4739), .A(n4738) );
  ao221 U2505 ( .Y(n4740), .A0(n5390), .A1(n5368), .B0(n5391), .B1(n5217), 
        .C0(n5392) );
  inv01 U2506 ( .Y(n4741), .A(n4740) );
  ao221 U2507 ( .Y(n4742), .A0(n5374), .A1(n5216), .B0(n5380), .B1(n5218), 
        .C0(n5452) );
  inv01 U2508 ( .Y(n4743), .A(n4742) );
  inv02 U2509 ( .Y(n5462), .A(n4744) );
  nor02 U2510 ( .Y(n4745), .A0(n5324), .A1(n5223) );
  nor02 U2511 ( .Y(n4746), .A0(n5403), .A1(n____return128) );
  nor02 U2512 ( .Y(n4744), .A0(n4745), .A1(n4746) );
  nand02 U2513 ( .Y(n5344), .A0(n4747), .A1(n4748) );
  inv02 U2514 ( .Y(n4749), .A(n5438) );
  inv01 U2515 ( .Y(n4750), .A(n5365) );
  inv01 U2516 ( .Y(n4751), .A(n5197) );
  inv01 U2517 ( .Y(n4752), .A(n5437) );
  inv02 U2518 ( .Y(n4753), .A(n5369) );
  nand02 U2519 ( .Y(n4754), .A0(n4751), .A1(n4755) );
  nand02 U2520 ( .Y(n4756), .A0(n4752), .A1(n4757) );
  nand02 U2521 ( .Y(n4758), .A0(n4753), .A1(n4759) );
  nand02 U2522 ( .Y(n4760), .A0(n4753), .A1(n4761) );
  nand02 U2523 ( .Y(n4762), .A0(n4749), .A1(n4750) );
  inv02 U2524 ( .Y(n4755), .A(n4762) );
  nand02 U2525 ( .Y(n4763), .A0(n4749), .A1(n4750) );
  inv01 U2526 ( .Y(n4757), .A(n4763) );
  nand02 U2527 ( .Y(n4764), .A0(n4749), .A1(n4751) );
  inv01 U2528 ( .Y(n4759), .A(n4764) );
  nand02 U2529 ( .Y(n4765), .A0(n4749), .A1(n4752) );
  inv01 U2530 ( .Y(n4761), .A(n4765) );
  nand02 U2531 ( .Y(n4766), .A0(n4754), .A1(n4756) );
  inv02 U2532 ( .Y(n4747), .A(n4766) );
  nand02 U2533 ( .Y(n4767), .A0(n4758), .A1(n4760) );
  inv02 U2534 ( .Y(n4748), .A(n4767) );
  nand02 U2535 ( .Y(n5328), .A0(n4768), .A1(n4769) );
  inv02 U2536 ( .Y(n4770), .A(n5420) );
  inv01 U2537 ( .Y(n4771), .A(n5365) );
  inv01 U2538 ( .Y(n4772), .A(n5217) );
  inv01 U2539 ( .Y(n4773), .A(n5390) );
  inv02 U2540 ( .Y(n4774), .A(n5391) );
  nand02 U2541 ( .Y(n4775), .A0(n4772), .A1(n4776) );
  nand02 U2542 ( .Y(n4777), .A0(n4773), .A1(n4778) );
  nand02 U2543 ( .Y(n4779), .A0(n4774), .A1(n4780) );
  nand02 U2544 ( .Y(n4781), .A0(n4774), .A1(n4782) );
  nand02 U2545 ( .Y(n4783), .A0(n4770), .A1(n4771) );
  inv02 U2546 ( .Y(n4776), .A(n4783) );
  nand02 U2547 ( .Y(n4784), .A0(n4770), .A1(n4771) );
  inv01 U2548 ( .Y(n4778), .A(n4784) );
  nand02 U2549 ( .Y(n4785), .A0(n4770), .A1(n4772) );
  inv01 U2550 ( .Y(n4780), .A(n4785) );
  nand02 U2551 ( .Y(n4786), .A0(n4770), .A1(n4773) );
  inv01 U2552 ( .Y(n4782), .A(n4786) );
  nand02 U2553 ( .Y(n4787), .A0(n4775), .A1(n4777) );
  inv02 U2554 ( .Y(n4768), .A(n4787) );
  nand02 U2555 ( .Y(n4788), .A0(n4779), .A1(n4781) );
  inv02 U2556 ( .Y(n4769), .A(n4788) );
  inv04 U2557 ( .Y(n5365), .A(n5213) );
  inv01 U2558 ( .Y(n5388), .A(n4789) );
  nor02 U2559 ( .Y(n4790), .A0(n5190), .A1(n5220) );
  nor02 U2560 ( .Y(n4791), .A0(n5164), .A1(n5219) );
  inv01 U2561 ( .Y(n4792), .A(n3333) );
  nor02 U2562 ( .Y(n4789), .A0(n4792), .A1(n4793) );
  nor02 U2563 ( .Y(n4794), .A0(n4790), .A1(n4791) );
  inv01 U2564 ( .Y(n4793), .A(n4794) );
  nor02 U2565 ( .Y(n4796), .A0(n5154), .A1(n5220) );
  nor02 U2566 ( .Y(n4797), .A0(n5150), .A1(n5219) );
  inv01 U2567 ( .Y(n4798), .A(n3404) );
  nor02 U2568 ( .Y(n4795), .A0(n4798), .A1(n4799) );
  nor02 U2569 ( .Y(n4800), .A0(n4796), .A1(n4797) );
  inv01 U2570 ( .Y(n4799), .A(n4800) );
  nor02 U2571 ( .Y(n4802), .A0(n5150), .A1(n5220) );
  nor02 U2572 ( .Y(n4803), .A0(n5190), .A1(n5219) );
  inv01 U2573 ( .Y(n4804), .A(n3329) );
  nor02 U2574 ( .Y(n4801), .A0(n4804), .A1(n4805) );
  nor02 U2575 ( .Y(n4806), .A0(n4802), .A1(n4803) );
  inv01 U2576 ( .Y(n4805), .A(n4806) );
  nand02 U2577 ( .Y(n5407), .A0(n3392), .A1(n4807) );
  inv01 U2578 ( .Y(n4808), .A(n5220) );
  inv01 U2579 ( .Y(n4809), .A(n5201) );
  inv01 U2580 ( .Y(n4810), .A(n5219) );
  inv01 U2581 ( .Y(n4811), .A(n5154) );
  nand02 U2582 ( .Y(n4812), .A0(n4808), .A1(n4809) );
  nand02 U2583 ( .Y(n4813), .A0(n4810), .A1(n4811) );
  nand02 U2584 ( .Y(n4814), .A0(n4812), .A1(n4813) );
  inv01 U2585 ( .Y(n4807), .A(n4814) );
  inv02 U2586 ( .Y(n5201), .A(n5200) );
  and02 U2587 ( .Y(n4816), .A0(n5212), .A1(n5197) );
  buf04 U2588 ( .Y(n5197), .A(n5397) );
  nand02 U2589 ( .Y(n5353), .A0(n4817), .A1(n4818) );
  inv02 U2590 ( .Y(n4819), .A(n5217) );
  inv02 U2591 ( .Y(n4820), .A(n5218) );
  inv02 U2592 ( .Y(n4821), .A(n5216) );
  inv02 U2593 ( .Y(n4822), .A(n5383) );
  inv02 U2594 ( .Y(n4823), .A(n5382) );
  inv02 U2595 ( .Y(n4824), .A(n5387) );
  nand02 U2596 ( .Y(n4825), .A0(n4821), .A1(n4826) );
  nand02 U2597 ( .Y(n4827), .A0(n4822), .A1(n4828) );
  nand02 U2598 ( .Y(n4829), .A0(n4823), .A1(n4830) );
  nand02 U2599 ( .Y(n4831), .A0(n4823), .A1(n4832) );
  nand02 U2600 ( .Y(n4833), .A0(n4824), .A1(n4834) );
  nand02 U2601 ( .Y(n4835), .A0(n4824), .A1(n4836) );
  nand02 U2602 ( .Y(n4837), .A0(n4824), .A1(n4838) );
  nand02 U2603 ( .Y(n4839), .A0(n4824), .A1(n4840) );
  nand02 U2604 ( .Y(n4841), .A0(n4819), .A1(n4820) );
  inv01 U2605 ( .Y(n4826), .A(n4841) );
  nand02 U2606 ( .Y(n4842), .A0(n4819), .A1(n4820) );
  inv01 U2607 ( .Y(n4828), .A(n4842) );
  nand02 U2608 ( .Y(n4843), .A0(n4819), .A1(n4821) );
  inv01 U2609 ( .Y(n4830), .A(n4843) );
  nand02 U2610 ( .Y(n4844), .A0(n4819), .A1(n4822) );
  inv01 U2611 ( .Y(n4832), .A(n4844) );
  nand02 U2612 ( .Y(n4845), .A0(n4820), .A1(n4821) );
  inv01 U2613 ( .Y(n4834), .A(n4845) );
  nand02 U2614 ( .Y(n4846), .A0(n4820), .A1(n4822) );
  inv01 U2615 ( .Y(n4836), .A(n4846) );
  nand02 U2616 ( .Y(n4847), .A0(n4821), .A1(n4823) );
  inv01 U2617 ( .Y(n4838), .A(n4847) );
  nand02 U2618 ( .Y(n4848), .A0(n4822), .A1(n4823) );
  inv01 U2619 ( .Y(n4840), .A(n4848) );
  nand02 U2620 ( .Y(n4849), .A0(n4825), .A1(n4827) );
  inv01 U2621 ( .Y(n4850), .A(n4849) );
  nand02 U2622 ( .Y(n4851), .A0(n4829), .A1(n4831) );
  inv01 U2623 ( .Y(n4852), .A(n4851) );
  nand02 U2624 ( .Y(n4853), .A0(n4850), .A1(n4852) );
  inv01 U2625 ( .Y(n4817), .A(n4853) );
  nand02 U2626 ( .Y(n4854), .A0(n4833), .A1(n4835) );
  inv01 U2627 ( .Y(n4855), .A(n4854) );
  nand02 U2628 ( .Y(n4856), .A0(n4837), .A1(n4839) );
  inv01 U2629 ( .Y(n4857), .A(n4856) );
  nand02 U2630 ( .Y(n4858), .A0(n4855), .A1(n4857) );
  inv01 U2631 ( .Y(n4818), .A(n4858) );
  ao22 U2632 ( .Y(n4859), .A0(n5371), .A1(n5209), .B0(n5364), .B1(n5212) );
  inv02 U2633 ( .Y(n4860), .A(n4859) );
  nand02 U2634 ( .Y(n4861), .A0(n5218), .A1(n5223) );
  ao22 U2635 ( .Y(n4862), .A0(n5378), .A1(n5212), .B0(n5379), .B1(n5209) );
  inv02 U2636 ( .Y(n4863), .A(n4862) );
  nand02 U2637 ( .Y(U403_U4_Z_0), .A0(n4864), .A1(n4865) );
  inv01 U2638 ( .Y(n4866), .A(n3327) );
  inv01 U2639 ( .Y(n4867), .A(n5223) );
  inv01 U2640 ( .Y(n4868), .A(n4957) );
  inv01 U2641 ( .Y(n4869), .A(n5469) );
  nand02 U2642 ( .Y(n4870), .A0(n4866), .A1(n4867) );
  nand02 U2643 ( .Y(n4871), .A0(n4866), .A1(n4868) );
  nand02 U2644 ( .Y(n4872), .A0(n4867), .A1(n4869) );
  nand02 U2645 ( .Y(n4873), .A0(n4868), .A1(n4869) );
  nand02 U2646 ( .Y(n4874), .A0(n4870), .A1(n4871) );
  inv02 U2647 ( .Y(n4864), .A(n4874) );
  nand02 U2648 ( .Y(n4875), .A0(n4872), .A1(n4873) );
  inv02 U2649 ( .Y(n4865), .A(n4875) );
  ao22 U2650 ( .Y(n4877), .A0(n5387), .A1(n5211), .B0(n5383), .B1(n5212) );
  inv02 U2651 ( .Y(n4878), .A(n4877) );
  inv02 U2652 ( .Y(n5390), .A(n4879) );
  nor02 U2653 ( .Y(n4880), .A0(n5186), .A1(n5220) );
  nor02 U2654 ( .Y(n4881), .A0(n5160), .A1(n5219) );
  inv01 U2655 ( .Y(n4882), .A(n5459) );
  nor02 U2656 ( .Y(n4879), .A0(n4882), .A1(n4883) );
  nor02 U2657 ( .Y(n4884), .A0(n4880), .A1(n4881) );
  inv01 U2658 ( .Y(n4883), .A(n4884) );
  buf04 U2659 ( .Y(n4885), .A(n5450) );
  inv02 U2660 ( .Y(n5386), .A(n4886) );
  nor02 U2661 ( .Y(n4887), .A0(n5160), .A1(n5220) );
  nor02 U2662 ( .Y(n4888), .A0(n5143), .A1(n5219) );
  inv01 U2663 ( .Y(n4889), .A(n5455) );
  nor02 U2664 ( .Y(n4886), .A0(n4889), .A1(n4890) );
  nor02 U2665 ( .Y(n4891), .A0(n4887), .A1(n4888) );
  inv01 U2666 ( .Y(n4890), .A(n4891) );
  inv02 U2667 ( .Y(n5375), .A(n4892) );
  nor02 U2668 ( .Y(n4893), .A0(n5164), .A1(n5220) );
  nor02 U2669 ( .Y(n4894), .A0(n5148), .A1(n5219) );
  inv01 U2670 ( .Y(n4895), .A(n3353) );
  nor02 U2671 ( .Y(n4892), .A0(n4895), .A1(n4896) );
  nor02 U2672 ( .Y(n4897), .A0(n4893), .A1(n4894) );
  inv01 U2673 ( .Y(n4896), .A(n4897) );
  inv02 U2674 ( .Y(n5372), .A(n4898) );
  nor02 U2675 ( .Y(n4899), .A0(n5148), .A1(n5220) );
  nor02 U2676 ( .Y(n4900), .A0(n5186), .A1(n5219) );
  inv01 U2677 ( .Y(n4901), .A(n3377) );
  nor02 U2678 ( .Y(n4898), .A0(n4901), .A1(n4902) );
  nor02 U2679 ( .Y(n4903), .A0(n4899), .A1(n4900) );
  inv01 U2680 ( .Y(n4902), .A(n4903) );
  inv02 U2681 ( .Y(n5469), .A(opb_i[23]) );
  ao22 U2682 ( .Y(n4904), .A0(n5467), .A1(n5329), .B0(n5425), .B1(n5468) );
  inv02 U2683 ( .Y(n4905), .A(n4904) );
  ao22 U2684 ( .Y(n4906), .A0(n5467), .A1(n5223), .B0(n5468), .B1(
        n____return128) );
  inv02 U2685 ( .Y(n4907), .A(n4906) );
  inv02 U2686 ( .Y(n5288), .A(n4907) );
  buf02 U2687 ( .Y(n4908), .A(opb_i[29]) );
  inv02 U2688 ( .Y(n4909), .A(n4908) );
  inv01 U2689 ( .Y(n4910), .A(n4908) );
  buf02 U2690 ( .Y(n4911), .A(opb_i[26]) );
  inv02 U2691 ( .Y(n4912), .A(n4911) );
  inv01 U2692 ( .Y(n4913), .A(n4911) );
  buf02 U2693 ( .Y(n4914), .A(opb_i[24]) );
  inv02 U2694 ( .Y(n4915), .A(n4914) );
  inv01 U2695 ( .Y(n4916), .A(n4914) );
  buf02 U2696 ( .Y(n4917), .A(opb_i[28]) );
  inv02 U2697 ( .Y(n4918), .A(n4917) );
  inv01 U2698 ( .Y(n4919), .A(n4917) );
  buf02 U2699 ( .Y(n4920), .A(opb_i[25]) );
  inv02 U2700 ( .Y(n4921), .A(n4920) );
  inv01 U2701 ( .Y(n4922), .A(n4920) );
  buf02 U2702 ( .Y(n4923), .A(opb_i[30]) );
  inv02 U2703 ( .Y(n4924), .A(n4923) );
  inv01 U2704 ( .Y(n4925), .A(n4923) );
  buf02 U2705 ( .Y(n4926), .A(opb_i[27]) );
  inv02 U2706 ( .Y(n4927), .A(n4926) );
  inv01 U2707 ( .Y(n4928), .A(n4926) );
  buf02 U2708 ( .Y(n4930), .A(opa_i[24]) );
  inv02 U2709 ( .Y(n4931), .A(n4930) );
  buf02 U2710 ( .Y(n4932), .A(opa_i[28]) );
  inv02 U2711 ( .Y(n4933), .A(n4932) );
  buf02 U2712 ( .Y(n4934), .A(opa_i[26]) );
  inv02 U2713 ( .Y(n4935), .A(n4934) );
  buf02 U2714 ( .Y(n4936), .A(opa_i[29]) );
  inv02 U2715 ( .Y(n4937), .A(n4936) );
  buf02 U2716 ( .Y(n4938), .A(opa_i[25]) );
  inv02 U2717 ( .Y(n4939), .A(n4938) );
  buf02 U2718 ( .Y(n4940), .A(opa_i[27]) );
  inv02 U2719 ( .Y(n4941), .A(n4940) );
  buf02 U2720 ( .Y(n4942), .A(opa_i[30]) );
  inv02 U2721 ( .Y(n4943), .A(n4942) );
  inv02 U2722 ( .Y(n5383), .A(n4944) );
  nor02 U2723 ( .Y(n4945), .A0(n5194), .A1(n5220) );
  nor02 U2724 ( .Y(n4946), .A0(n5162), .A1(n5219) );
  inv01 U2725 ( .Y(n4947), .A(n3337) );
  nor02 U2726 ( .Y(n4944), .A0(n4947), .A1(n4948) );
  nor02 U2727 ( .Y(n4949), .A0(n4945), .A1(n4946) );
  inv01 U2728 ( .Y(n4948), .A(n4949) );
  inv02 U2729 ( .Y(n5391), .A(n4950) );
  nor02 U2730 ( .Y(n4951), .A0(n5158), .A1(n5220) );
  nor02 U2731 ( .Y(n4952), .A0(n5141), .A1(n5219) );
  inv01 U2732 ( .Y(n4953), .A(n3369) );
  nor02 U2733 ( .Y(n4950), .A0(n4953), .A1(n4954) );
  nor02 U2734 ( .Y(n4955), .A0(n4951), .A1(n4952) );
  inv01 U2735 ( .Y(n4954), .A(n4955) );
  buf02 U2736 ( .Y(n4956), .A(opa_i[23]) );
  inv02 U2737 ( .Y(n4957), .A(n4956) );
  inv02 U2738 ( .Y(n5369), .A(n4958) );
  nor02 U2739 ( .Y(n4959), .A0(n5182), .A1(n5220) );
  nor02 U2740 ( .Y(n4960), .A0(n5158), .A1(n5219) );
  inv01 U2741 ( .Y(n4961), .A(n3351) );
  nor02 U2742 ( .Y(n4958), .A0(n4961), .A1(n4962) );
  nor02 U2743 ( .Y(n4963), .A0(n4959), .A1(n4960) );
  inv01 U2744 ( .Y(n4962), .A(n4963) );
  inv02 U2745 ( .Y(n5378), .A(n4964) );
  nor02 U2746 ( .Y(n4965), .A0(n5162), .A1(n5220) );
  nor02 U2747 ( .Y(n4966), .A0(n5156), .A1(n5219) );
  inv01 U2748 ( .Y(n4967), .A(n3381) );
  nor02 U2749 ( .Y(n4964), .A0(n4967), .A1(n4968) );
  nor02 U2750 ( .Y(n4969), .A0(n4965), .A1(n4966) );
  inv01 U2751 ( .Y(n4968), .A(n4969) );
  inv02 U2752 ( .Y(n5374), .A(n4970) );
  nor02 U2753 ( .Y(n4971), .A0(n5188), .A1(n5220) );
  nor02 U2754 ( .Y(n4972), .A0(n5166), .A1(n5219) );
  inv01 U2755 ( .Y(n4973), .A(n3331) );
  nor02 U2756 ( .Y(n4970), .A0(n4973), .A1(n4974) );
  nor02 U2757 ( .Y(n4975), .A0(n4971), .A1(n4972) );
  inv01 U2758 ( .Y(n4974), .A(n4975) );
  nand02 U2759 ( .Y(n5351), .A0(n4976), .A1(n4977) );
  inv02 U2760 ( .Y(n4978), .A(n5210) );
  inv02 U2761 ( .Y(n4979), .A(n5019) );
  inv02 U2762 ( .Y(n4980), .A(n5212) );
  inv02 U2763 ( .Y(n4981), .A(n5374) );
  inv02 U2764 ( .Y(n4982), .A(n5379) );
  inv02 U2765 ( .Y(n4983), .A(n5378) );
  nand02 U2766 ( .Y(n4984), .A0(n4980), .A1(n4985) );
  nand02 U2767 ( .Y(n4986), .A0(n4981), .A1(n4987) );
  nand02 U2768 ( .Y(n4988), .A0(n4982), .A1(n4989) );
  nand02 U2769 ( .Y(n4990), .A0(n4982), .A1(n4991) );
  nand02 U2770 ( .Y(n4992), .A0(n4983), .A1(n4993) );
  nand02 U2771 ( .Y(n4994), .A0(n4983), .A1(n4995) );
  nand02 U2772 ( .Y(n4996), .A0(n4983), .A1(n4997) );
  nand02 U2773 ( .Y(n4998), .A0(n4983), .A1(n4999) );
  nand02 U2774 ( .Y(n5000), .A0(n4978), .A1(n4979) );
  inv01 U2775 ( .Y(n4985), .A(n5000) );
  nand02 U2776 ( .Y(n5001), .A0(n4978), .A1(n4979) );
  inv01 U2777 ( .Y(n4987), .A(n5001) );
  nand02 U2778 ( .Y(n5002), .A0(n4978), .A1(n4980) );
  inv01 U2779 ( .Y(n4989), .A(n5002) );
  nand02 U2780 ( .Y(n5003), .A0(n4978), .A1(n4981) );
  inv01 U2781 ( .Y(n4991), .A(n5003) );
  nand02 U2782 ( .Y(n5004), .A0(n4979), .A1(n4980) );
  inv01 U2783 ( .Y(n4993), .A(n5004) );
  nand02 U2784 ( .Y(n5005), .A0(n4979), .A1(n4981) );
  inv01 U2785 ( .Y(n4995), .A(n5005) );
  nand02 U2786 ( .Y(n5006), .A0(n4980), .A1(n4982) );
  inv01 U2787 ( .Y(n4997), .A(n5006) );
  nand02 U2788 ( .Y(n5007), .A0(n4981), .A1(n4982) );
  inv01 U2789 ( .Y(n4999), .A(n5007) );
  nand02 U2790 ( .Y(n5008), .A0(n4984), .A1(n4986) );
  inv02 U2791 ( .Y(n5009), .A(n5008) );
  nand02 U2792 ( .Y(n5010), .A0(n4988), .A1(n4990) );
  inv02 U2793 ( .Y(n5011), .A(n5010) );
  nand02 U2794 ( .Y(n5012), .A0(n5009), .A1(n5011) );
  inv02 U2795 ( .Y(n4976), .A(n5012) );
  nand02 U2796 ( .Y(n5013), .A0(n4992), .A1(n4994) );
  inv02 U2797 ( .Y(n5014), .A(n5013) );
  nand02 U2798 ( .Y(n5015), .A0(n4996), .A1(n4998) );
  inv01 U2799 ( .Y(n5016), .A(n5015) );
  nand02 U2800 ( .Y(n5017), .A0(n5014), .A1(n5016) );
  inv02 U2801 ( .Y(n4977), .A(n5017) );
  inv02 U2802 ( .Y(n5210), .A(n5208) );
  nand02 U2803 ( .Y(n5018), .A0(s_exp_diff_3_), .A1(n5433) );
  inv02 U2804 ( .Y(n5019), .A(n5018) );
  inv02 U2805 ( .Y(n5432), .A(n5020) );
  nor02 U2806 ( .Y(n5021), .A0(n5184), .A1(n5220) );
  nor02 U2807 ( .Y(n5022), .A0(n5196), .A1(n5219) );
  inv01 U2808 ( .Y(n5023), .A(n3335) );
  nor02 U2809 ( .Y(n5020), .A0(n5023), .A1(n5024) );
  nor02 U2810 ( .Y(n5025), .A0(n5021), .A1(n5022) );
  inv01 U2811 ( .Y(n5024), .A(n5025) );
  inv02 U2812 ( .Y(n5362), .A(n5026) );
  nor02 U2813 ( .Y(n5027), .A0(n5166), .A1(n5220) );
  nor02 U2814 ( .Y(n5028), .A0(n5152), .A1(n5219) );
  inv01 U2815 ( .Y(n5029), .A(n3375) );
  nor02 U2816 ( .Y(n5026), .A0(n5029), .A1(n5030) );
  nor02 U2817 ( .Y(n5031), .A0(n5027), .A1(n5028) );
  inv01 U2818 ( .Y(n5030), .A(n5031) );
  inv02 U2819 ( .Y(n5364), .A(n5032) );
  nor02 U2820 ( .Y(n5033), .A0(n5156), .A1(n5220) );
  nor02 U2821 ( .Y(n5034), .A0(n5184), .A1(n5219) );
  inv01 U2822 ( .Y(n5035), .A(n3371) );
  nor02 U2823 ( .Y(n5032), .A0(n5035), .A1(n5036) );
  nor02 U2824 ( .Y(n5037), .A0(n5033), .A1(n5034) );
  inv01 U2825 ( .Y(n5036), .A(n5037) );
  nand02 U2826 ( .Y(n5347), .A0(n5038), .A1(n5039) );
  inv02 U2827 ( .Y(n5040), .A(n5212) );
  inv02 U2828 ( .Y(n5041), .A(n5434) );
  inv02 U2829 ( .Y(n5042), .A(n5211) );
  inv02 U2830 ( .Y(n5043), .A(n5432) );
  inv02 U2831 ( .Y(n5044), .A(n5019) );
  inv02 U2832 ( .Y(n5045), .A(n5394) );
  nand02 U2833 ( .Y(n5046), .A0(n5042), .A1(n5047) );
  nand02 U2834 ( .Y(n5048), .A0(n5043), .A1(n5049) );
  nand02 U2835 ( .Y(n5050), .A0(n5044), .A1(n5051) );
  nand02 U2836 ( .Y(n5052), .A0(n5044), .A1(n5053) );
  nand02 U2837 ( .Y(n5054), .A0(n5045), .A1(n5055) );
  nand02 U2838 ( .Y(n5056), .A0(n5045), .A1(n5057) );
  nand02 U2839 ( .Y(n5058), .A0(n5045), .A1(n5059) );
  nand02 U2840 ( .Y(n5060), .A0(n5045), .A1(n5061) );
  nand02 U2841 ( .Y(n5062), .A0(n5040), .A1(n5041) );
  inv01 U2842 ( .Y(n5047), .A(n5062) );
  nand02 U2843 ( .Y(n5063), .A0(n5040), .A1(n5041) );
  inv01 U2844 ( .Y(n5049), .A(n5063) );
  nand02 U2845 ( .Y(n5064), .A0(n5040), .A1(n5042) );
  inv01 U2846 ( .Y(n5051), .A(n5064) );
  nand02 U2847 ( .Y(n5065), .A0(n5040), .A1(n5043) );
  inv01 U2848 ( .Y(n5053), .A(n5065) );
  nand02 U2849 ( .Y(n5066), .A0(n5041), .A1(n5042) );
  inv01 U2850 ( .Y(n5055), .A(n5066) );
  nand02 U2851 ( .Y(n5067), .A0(n5041), .A1(n5043) );
  inv01 U2852 ( .Y(n5057), .A(n5067) );
  nand02 U2853 ( .Y(n5068), .A0(n5042), .A1(n5044) );
  inv01 U2854 ( .Y(n5059), .A(n5068) );
  nand02 U2855 ( .Y(n5069), .A0(n5043), .A1(n5044) );
  inv01 U2856 ( .Y(n5061), .A(n5069) );
  nand02 U2857 ( .Y(n5070), .A0(n5046), .A1(n5048) );
  inv02 U2858 ( .Y(n5071), .A(n5070) );
  nand02 U2859 ( .Y(n5072), .A0(n5050), .A1(n5052) );
  inv02 U2860 ( .Y(n5073), .A(n5072) );
  nand02 U2861 ( .Y(n5074), .A0(n5071), .A1(n5073) );
  inv02 U2862 ( .Y(n5038), .A(n5074) );
  nand02 U2863 ( .Y(n5075), .A0(n5054), .A1(n5056) );
  inv02 U2864 ( .Y(n5076), .A(n5075) );
  nand02 U2865 ( .Y(n5077), .A0(n5058), .A1(n5060) );
  inv01 U2866 ( .Y(n5078), .A(n5077) );
  nand02 U2867 ( .Y(n5079), .A0(n5076), .A1(n5078) );
  inv02 U2868 ( .Y(n5039), .A(n5079) );
  nand02 U2869 ( .Y(n5349), .A0(n5080), .A1(n5081) );
  inv02 U2870 ( .Y(n5082), .A(n5210) );
  inv02 U2871 ( .Y(n5083), .A(n5019) );
  inv02 U2872 ( .Y(n5084), .A(n5212) );
  inv02 U2873 ( .Y(n5085), .A(n5362) );
  inv02 U2874 ( .Y(n5086), .A(n5371) );
  inv02 U2875 ( .Y(n5087), .A(n5364) );
  nand02 U2876 ( .Y(n5088), .A0(n5084), .A1(n5089) );
  nand02 U2877 ( .Y(n5090), .A0(n5085), .A1(n5091) );
  nand02 U2878 ( .Y(n5092), .A0(n5086), .A1(n5093) );
  nand02 U2879 ( .Y(n5094), .A0(n5086), .A1(n5095) );
  nand02 U2880 ( .Y(n5096), .A0(n5087), .A1(n5097) );
  nand02 U2881 ( .Y(n5098), .A0(n5087), .A1(n5099) );
  nand02 U2882 ( .Y(n5100), .A0(n5087), .A1(n5101) );
  nand02 U2883 ( .Y(n5102), .A0(n5087), .A1(n5103) );
  nand02 U2884 ( .Y(n5104), .A0(n5082), .A1(n5083) );
  inv01 U2885 ( .Y(n5089), .A(n5104) );
  nand02 U2886 ( .Y(n5105), .A0(n5082), .A1(n5083) );
  inv01 U2887 ( .Y(n5091), .A(n5105) );
  nand02 U2888 ( .Y(n5106), .A0(n5082), .A1(n5084) );
  inv01 U2889 ( .Y(n5093), .A(n5106) );
  nand02 U2890 ( .Y(n5107), .A0(n5082), .A1(n5085) );
  inv01 U2891 ( .Y(n5095), .A(n5107) );
  nand02 U2892 ( .Y(n5108), .A0(n5083), .A1(n5084) );
  inv01 U2893 ( .Y(n5097), .A(n5108) );
  nand02 U2894 ( .Y(n5109), .A0(n5083), .A1(n5085) );
  inv01 U2895 ( .Y(n5099), .A(n5109) );
  nand02 U2896 ( .Y(n5110), .A0(n5084), .A1(n5086) );
  inv01 U2897 ( .Y(n5101), .A(n5110) );
  nand02 U2898 ( .Y(n5111), .A0(n5085), .A1(n5086) );
  inv01 U2899 ( .Y(n5103), .A(n5111) );
  nand02 U2900 ( .Y(n5112), .A0(n5088), .A1(n5090) );
  inv02 U2901 ( .Y(n5113), .A(n5112) );
  nand02 U2902 ( .Y(n5114), .A0(n5092), .A1(n5094) );
  inv01 U2903 ( .Y(n5115), .A(n5114) );
  nand02 U2904 ( .Y(n5116), .A0(n5113), .A1(n5115) );
  inv02 U2905 ( .Y(n5080), .A(n5116) );
  nand02 U2906 ( .Y(n5117), .A0(n5096), .A1(n5098) );
  inv02 U2907 ( .Y(n5118), .A(n5117) );
  nand02 U2908 ( .Y(n5119), .A0(n5100), .A1(n5102) );
  inv01 U2909 ( .Y(n5120), .A(n5119) );
  nand02 U2910 ( .Y(n5121), .A0(n5118), .A1(n5120) );
  inv02 U2911 ( .Y(n5081), .A(n5121) );
  inv02 U2912 ( .Y(n5434), .A(n5330) );
  inv02 U2913 ( .Y(n5380), .A(n5122) );
  nor02 U2914 ( .Y(n5123), .A0(n5143), .A1(n5220) );
  nor02 U2915 ( .Y(n5124), .A0(n5182), .A1(n5219) );
  inv01 U2916 ( .Y(n5125), .A(n3383) );
  nor02 U2917 ( .Y(n5122), .A0(n5125), .A1(n5126) );
  nor02 U2918 ( .Y(n5127), .A0(n5123), .A1(n5124) );
  inv01 U2919 ( .Y(n5126), .A(n5127) );
  inv02 U2920 ( .Y(n5382), .A(n5128) );
  nor02 U2921 ( .Y(n5129), .A0(n5141), .A1(n5220) );
  nor02 U2922 ( .Y(n5130), .A0(n5188), .A1(n5219) );
  inv01 U2923 ( .Y(n5131), .A(n3373) );
  nor02 U2924 ( .Y(n5128), .A0(n5131), .A1(n5132) );
  nor02 U2925 ( .Y(n5133), .A0(n5129), .A1(n5130) );
  inv01 U2926 ( .Y(n5132), .A(n5133) );
  inv02 U2927 ( .Y(n5394), .A(n5134) );
  nor02 U2928 ( .Y(n5135), .A0(n5152), .A1(n5220) );
  nor02 U2929 ( .Y(n5136), .A0(n5194), .A1(n5219) );
  inv01 U2930 ( .Y(n5137), .A(n3379) );
  nor02 U2931 ( .Y(n5134), .A0(n5137), .A1(n5138) );
  nor02 U2932 ( .Y(n5139), .A0(n5135), .A1(n5136) );
  inv01 U2933 ( .Y(n5138), .A(n5139) );
  inv02 U2934 ( .Y(n5194), .A(n5193) );
  ao22 U2935 ( .Y(n5140), .A0(opa_i[13]), .A1(n5223), .B0(opb_i[13]), .B1(
        n____return128) );
  inv02 U2936 ( .Y(n5141), .A(n5140) );
  inv02 U2937 ( .Y(n5286), .A(n5141) );
  ao22 U2938 ( .Y(n5142), .A0(opa_i[10]), .A1(n5223), .B0(opb_i[10]), .B1(
        n____return128) );
  inv02 U2939 ( .Y(n5143), .A(n5142) );
  inv02 U2940 ( .Y(n5371), .A(n5144) );
  nor02 U2941 ( .Y(n5145), .A0(n4907), .A1(n5220) );
  nor02 U2942 ( .Y(n5146), .A0(n5199), .A1(n4885) );
  nor02 U2943 ( .Y(n5144), .A0(n5145), .A1(n5146) );
  inv02 U2944 ( .Y(n5305), .A(n5143) );
  ao22 U2945 ( .Y(n5147), .A0(opa_i[7]), .A1(n5222), .B0(opb_i[7]), .B1(
        n____return128) );
  inv02 U2946 ( .Y(n5148), .A(n5147) );
  ao22 U2947 ( .Y(n5149), .A0(opa_i[4]), .A1(n5222), .B0(opb_i[4]), .B1(
        n____return128) );
  inv02 U2948 ( .Y(n5150), .A(n5149) );
  inv02 U2949 ( .Y(n5294), .A(n5148) );
  inv02 U2950 ( .Y(n5306), .A(n5150) );
  ao22 U2951 ( .Y(n5151), .A0(opa_i[16]), .A1(n5223), .B0(opb_i[16]), .B1(
        n____return128) );
  inv02 U2952 ( .Y(n5152), .A(n5151) );
  inv02 U2953 ( .Y(n5311), .A(n5152) );
  ao22 U2954 ( .Y(n5153), .A0(opa_i[3]), .A1(n5223), .B0(opb_i[3]), .B1(
        n____return128) );
  inv02 U2955 ( .Y(n5154), .A(n5153) );
  inv02 U2956 ( .Y(n5283), .A(n5154) );
  ao22 U2957 ( .Y(n5155), .A0(opa_i[19]), .A1(n5222), .B0(opb_i[19]), .B1(
        n____return128) );
  inv02 U2958 ( .Y(n5156), .A(n5155) );
  inv02 U2959 ( .Y(n5292), .A(n5156) );
  ao22 U2960 ( .Y(n5157), .A0(opa_i[12]), .A1(n5223), .B0(opb_i[12]), .B1(
        n____return128) );
  inv02 U2961 ( .Y(n5158), .A(n5157) );
  ao22 U2962 ( .Y(n5159), .A0(opa_i[9]), .A1(n5223), .B0(opb_i[9]), .B1(
        n____return128) );
  inv02 U2963 ( .Y(n5160), .A(n5159) );
  inv02 U2964 ( .Y(n5308), .A(n5158) );
  inv02 U2965 ( .Y(n5296), .A(n5160) );
  ao22 U2966 ( .Y(n5161), .A0(opa_i[18]), .A1(n5223), .B0(opb_i[18]), .B1(
        n____return128) );
  inv02 U2967 ( .Y(n5162), .A(n5161) );
  ao22 U2968 ( .Y(n5163), .A0(opa_i[6]), .A1(n5223), .B0(opb_i[6]), .B1(
        n____return128) );
  inv02 U2969 ( .Y(n5164), .A(n5163) );
  inv02 U2970 ( .Y(n5315), .A(n5162) );
  inv02 U2971 ( .Y(n5309), .A(n5164) );
  ao22 U2972 ( .Y(n5165), .A0(opa_i[15]), .A1(n5222), .B0(opb_i[15]), .B1(
        n____return128) );
  inv02 U2973 ( .Y(n5166), .A(n5165) );
  inv02 U2974 ( .Y(n5287), .A(n5166) );
  inv02 U2975 ( .Y(n5387), .A(n5167) );
  nor02 U2976 ( .Y(n5168), .A0(n5196), .A1(n5220) );
  nor02 U2977 ( .Y(n5169), .A0(n5199), .A1(n5219) );
  inv01 U2978 ( .Y(n5170), .A(n3355) );
  nor02 U2979 ( .Y(n5167), .A0(n5170), .A1(n5171) );
  nor02 U2980 ( .Y(n5172), .A0(n5168), .A1(n5169) );
  inv01 U2981 ( .Y(n5171), .A(n5172) );
  inv02 U2982 ( .Y(n5337), .A(n5387) );
  inv02 U2983 ( .Y(n5379), .A(n5173) );
  nor02 U2984 ( .Y(n5174), .A0(n5196), .A1(n4885) );
  nor02 U2985 ( .Y(n5175), .A0(n4907), .A1(n5219) );
  nor02 U2986 ( .Y(n5176), .A0(n5199), .A1(n5220) );
  nor02 U2987 ( .Y(n5173), .A0(n5176), .A1(n5177) );
  nor02 U2988 ( .Y(n5178), .A0(n5174), .A1(n5175) );
  inv01 U2989 ( .Y(n5177), .A(n5178) );
  inv02 U2990 ( .Y(n5335), .A(n5379) );
  inv02 U2991 ( .Y(n5199), .A(n5198) );
  inv02 U2992 ( .Y(n5196), .A(n5195) );
  ao22 U2993 ( .Y(n5179), .A0(opa_i[0]), .A1(n5223), .B0(opb_i[0]), .B1(
        n____return128) );
  inv02 U2994 ( .Y(n5180), .A(n5179) );
  inv02 U2995 ( .Y(n5278), .A(n5180) );
  ao22 U2996 ( .Y(n5181), .A0(opa_i[11]), .A1(n5222), .B0(opb_i[11]), .B1(
        n____return128) );
  inv02 U2997 ( .Y(n5182), .A(n5181) );
  inv02 U2998 ( .Y(n5299), .A(n5182) );
  ao22 U2999 ( .Y(n5183), .A0(opa_i[20]), .A1(n5223), .B0(opb_i[20]), .B1(
        n____return128) );
  inv02 U3000 ( .Y(n5184), .A(n5183) );
  ao22 U3001 ( .Y(n5185), .A0(opa_i[8]), .A1(n5222), .B0(opb_i[8]), .B1(
        n____return128) );
  inv02 U3002 ( .Y(n5186), .A(n5185) );
  ao22 U3003 ( .Y(n5187), .A0(opa_i[14]), .A1(n5223), .B0(opb_i[14]), .B1(
        n____return128) );
  inv02 U3004 ( .Y(n5188), .A(n5187) );
  ao22 U3005 ( .Y(n5189), .A0(opa_i[5]), .A1(n5222), .B0(opb_i[5]), .B1(
        n____return128) );
  inv02 U3006 ( .Y(n5190), .A(n5189) );
  inv02 U3007 ( .Y(n5307), .A(n5184) );
  inv02 U3008 ( .Y(n5303), .A(n5186) );
  inv02 U3009 ( .Y(n5313), .A(n5188) );
  inv02 U3010 ( .Y(n5295), .A(n5190) );
  or02 U3011 ( .Y(n5191), .A0(n5464), .A1(s_exp_diff_4_) );
  inv02 U3012 ( .Y(n5192), .A(n5191) );
  ao22 U3013 ( .Y(n5193), .A0(opa_i[17]), .A1(n5222), .B0(opb_i[17]), .B1(
        n____return128) );
  inv02 U3014 ( .Y(n5290), .A(n5194) );
  ao22 U3015 ( .Y(n5195), .A0(opa_i[21]), .A1(n5222), .B0(opb_i[21]), .B1(
        n____return128) );
  ao22 U3016 ( .Y(n5198), .A0(opa_i[22]), .A1(n5222), .B0(opb_i[22]), .B1(
        n____return128) );
  ao22 U3017 ( .Y(n5200), .A0(opa_i[2]), .A1(n5222), .B0(opb_i[2]), .B1(
        n____return128) );
  buf02 U3018 ( .Y(n5202), .A(n5431) );
  buf02 U3019 ( .Y(n5203), .A(n5431) );
  buf02 U3020 ( .Y(n5204), .A(n5341) );
  buf02 U3021 ( .Y(n5205), .A(n5341) );
  buf04 U3022 ( .Y(n5206), .A(n5472) );
  inv04 U3023 ( .Y(n5470), .A(n4905) );
  buf04 U3024 ( .Y(n5207), .A(n5473) );
  inv02 U3025 ( .Y(n5208), .A(n5415) );
  inv02 U3026 ( .Y(n5209), .A(n5208) );
  inv02 U3027 ( .Y(n5211), .A(n5208) );
  buf04 U3028 ( .Y(n5212), .A(n5413) );
  nand02 U3029 ( .Y(n5213), .A0(s_exp_diff_3_), .A1(n5214) );
  nand02 U3030 ( .Y(n5215), .A0(s_exp_diff_2_), .A1(n5192) );
  inv01 U3031 ( .Y(n5214), .A(n5215) );
  inv08 U3032 ( .Y(n5418), .A(n4885) );
  inv08 U3033 ( .Y(n5419), .A(n4929) );
  buf16 U3034 ( .Y(n5219), .A(n5416) );
  buf16 U3035 ( .Y(n5220), .A(n5417) );
  buf12 U3036 ( .Y(n5221), .A(n____return128) );
  inv16 U3037 ( .Y(n5222), .A(n5221) );
  inv16 U3038 ( .Y(n5223), .A(n5221) );
  inv01 U3039 ( .Y(n5274), .A(n5228) );
  nor02 U3040 ( .Y(n5273), .A0(n5232), .A1(n5229) );
  nor02 U3041 ( .Y(n5272), .A0(n5233), .A1(n5231) );
  inv01 U3042 ( .Y(n5271), .A(n5278) );
  and02 U3043 ( .Y(n5224), .A0(n5283), .A1(n5284) );
  nor02 U3044 ( .Y(n5282), .A0(n5239), .A1(n3463) );
  inv01 U3045 ( .Y(n5281), .A(n5241) );
  inv01 U3046 ( .Y(n5280), .A(n5240) );
  inv01 U3047 ( .Y(n5263), .A(n3424) );
  inv01 U3048 ( .Y(n5262), .A(n5229) );
  nor02 U3049 ( .Y(n5261), .A0(n5232), .A1(n5233) );
  nor02 U3050 ( .Y(n5260), .A0(n5234), .A1(n4305) );
  nand02 U3051 ( .Y(n5267), .A0(n5180), .A1(n5268) );
  nor02 U3052 ( .Y(n5266), .A0(n5239), .A1(n5235) );
  inv01 U3053 ( .Y(n5265), .A(n5242) );
  inv01 U3054 ( .Y(n5264), .A(n5240) );
  nand03 U3055 ( .Y(n5245), .A0(n5247), .A1(n3875), .A2(n5246) );
  inv01 U3056 ( .Y(n5247), .A(n5229) );
  inv01 U3057 ( .Y(n5246), .A(n4305) );
  nand03 U3058 ( .Y(n5244), .A0(n5249), .A1(n3873), .A2(n5248) );
  nor02 U3059 ( .Y(n5249), .A0(n3463), .A1(n5239) );
  nor02 U3060 ( .Y(n5248), .A0(n5243), .A1(n3424) );
  inv01 U3061 ( .Y(n5255), .A(n5226) );
  inv01 U3062 ( .Y(n5254), .A(n5230) );
  nor02 U3063 ( .Y(n5253), .A0(n5231), .A1(n5232) );
  nor02 U3064 ( .Y(n5252), .A0(n5234), .A1(n4305) );
  nand03 U3065 ( .Y(n5250), .A0(n3461), .A1(n5257), .A2(n5256) );
  nor02 U3066 ( .Y(n5257), .A0(n5238), .A1(n3463) );
  inv01 U3067 ( .Y(n5256), .A(n5243) );
  or02 U3069 ( .Y(s_rzeros_4_), .A0(n5244), .A1(n5245) );
  or02 U3070 ( .Y(s_rzeros_3_), .A0(n5250), .A1(n5251) );
  nand04 U3071 ( .Y(n5251), .A0(n5252), .A1(n5253), .A2(n5254), .A3(n5255) );
  or02 U3072 ( .Y(s_rzeros_2_), .A0(n5258), .A1(n5259) );
  nand04 U3073 ( .Y(n5259), .A0(n5260), .A1(n5261), .A2(n5262), .A3(n5263) );
  nand04 U3074 ( .Y(n5258), .A0(n5264), .A1(n5265), .A2(n5266), .A3(n5267) );
  or02 U3075 ( .Y(s_rzeros_1_), .A0(n5269), .A1(n5270) );
  nand04 U3076 ( .Y(n5270), .A0(n5271), .A1(n5272), .A2(n5273), .A3(n5274) );
  inv01 U3077 ( .Y(n5230), .A(n5275) );
  inv01 U3078 ( .Y(n5229), .A(n5276) );
  nand04 U3079 ( .Y(n5269), .A0(n5280), .A1(n5281), .A2(n5282), .A3(n3459) );
  and02 U3080 ( .Y(n5236), .A0(n5285), .A1(n5286) );
  and03 U3081 ( .Y(n5237), .A0(n5188), .A1(n5287), .A2(n4043) );
  and02 U3082 ( .Y(n5235), .A0(n3943), .A1(n5290) );
  and02 U3083 ( .Y(n5239), .A0(n5291), .A1(n5292) );
  and02 U3084 ( .Y(n5241), .A0(n5293), .A1(n5294) );
  and02 U3085 ( .Y(n5238), .A0(n4045), .A1(n5295) );
  and03 U3086 ( .Y(n5242), .A0(n5186), .A1(n5296), .A2(n4217) );
  and03 U3087 ( .Y(n5243), .A0(n5298), .A1(n5297), .A2(n5184) );
  and02 U3088 ( .Y(n5240), .A0(n4047), .A1(n5299) );
  nand04 U3089 ( .Y(s_rzeros_0_), .A0(n3419), .A1(n5180), .A2(n5300), .A3(
        n5301) );
  and02 U3090 ( .Y(n5231), .A0(n4217), .A1(n5303) );
  and02 U3091 ( .Y(n5234), .A0(n5304), .A1(n5305) );
  and02 U3092 ( .Y(n5233), .A0(n3396), .A1(n5306) );
  nand03 U3093 ( .Y(n5302), .A0(n5277), .A1(n5275), .A2(n5276) );
  nand02 U3094 ( .Y(n5276), .A0(n5298), .A1(n5307) );
  nand03 U3095 ( .Y(n5277), .A0(n5182), .A1(n5308), .A2(n4047) );
  nand03 U3096 ( .Y(n5275), .A0(n5190), .A1(n5309), .A2(n4045) );
  and02 U3097 ( .Y(n5228), .A0(n5310), .A1(n5311) );
  and02 U3098 ( .Y(n5226), .A0(n5289), .A1(n5312) );
  and02 U3099 ( .Y(n5227), .A0(n4043), .A1(n5313) );
  inv01 U3100 ( .Y(n5316), .A(opb_i[6]) );
  inv01 U3101 ( .Y(n5318), .A(opb_i[5]) );
  inv01 U3102 ( .Y(n5320), .A(opb_i[4]) );
  inv01 U3103 ( .Y(n5321), .A(opb_i[3]) );
  inv01 U3104 ( .Y(n5322), .A(opb_i[2]) );
  inv01 U3105 ( .Y(n5326), .A(opb_i[0]) );
  inv01 U3106 ( .Y(n5332), .A(opb_i[22]) );
  inv01 U3107 ( .Y(n5334), .A(opb_i[21]) );
  nand02 U3108 ( .Y(n5331), .A0(n5218), .A1(n____return128) );
  inv01 U3109 ( .Y(n5336), .A(opb_i[20]) );
  inv01 U3110 ( .Y(n5339), .A(opb_i[19]) );
  inv01 U3111 ( .Y(n5342), .A(opb_i[18]) );
  inv01 U3112 ( .Y(n5343), .A(opb_i[17]) );
  inv01 U3113 ( .Y(n5345), .A(opb_i[16]) );
  inv01 U3114 ( .Y(n5346), .A(opb_i[15]) );
  inv01 U3115 ( .Y(n5348), .A(opb_i[14]) );
  nand02 U3116 ( .Y(n5341), .A0(n5192), .A1(n____return128) );
  inv01 U3117 ( .Y(n5350), .A(opb_i[13]) );
  inv01 U3118 ( .Y(n5352), .A(opb_i[12]) );
  inv01 U3119 ( .Y(n5354), .A(opb_i[11]) );
  inv01 U3120 ( .Y(n5355), .A(opb_i[10]) );
  inv01 U3121 ( .Y(n5356), .A(opb_i[9]) );
  inv01 U3122 ( .Y(n5357), .A(opb_i[8]) );
  inv01 U3123 ( .Y(n5359), .A(opb_i[7]) );
  inv01 U3124 ( .Y(n5361), .A(opa_i[6]) );
  inv01 U3125 ( .Y(n5366), .A(n5367) );
  inv01 U3126 ( .Y(n5373), .A(opa_i[5]) );
  inv01 U3127 ( .Y(n5376), .A(n5377) );
  inv01 U3128 ( .Y(n5381), .A(opa_i[4]) );
  inv01 U3129 ( .Y(n5384), .A(n5385) );
  inv01 U3130 ( .Y(n5389), .A(opa_i[3]) );
  inv01 U3131 ( .Y(n5392), .A(n5393) );
  inv01 U3132 ( .Y(n5398), .A(opa_i[2]) );
  inv01 U3133 ( .Y(n5399), .A(n5400) );
  inv01 U3134 ( .Y(n5404), .A(n5405) );
  inv01 U3135 ( .Y(n5406), .A(n4863) );
  inv01 U3136 ( .Y(n5408), .A(opa_i[0]) );
  nand02 U3137 ( .Y(n5327), .A0(n5409), .A1(n5410) );
  mux21 U3138 ( .Y(n5410), .A0(n5411), .A1(n4878), .S0(s_exp_diff_4_) );
  ao22 U3139 ( .Y(n5412), .A0(n5212), .A1(n5414), .B0(n5211), .B1(n5388) );
  inv01 U3140 ( .Y(n5420), .A(n5421) );
  inv01 U3141 ( .Y(n5422), .A(n5347) );
  inv01 U3142 ( .Y(n5333), .A(n5371) );
  inv01 U3143 ( .Y(n5427), .A(opa_i[22]) );
  inv01 U3144 ( .Y(n5428), .A(opa_i[21]) );
  nand02 U3145 ( .Y(n5426), .A0(n5218), .A1(n5223) );
  inv01 U3146 ( .Y(n5429), .A(opa_i[20]) );
  nor02 U3147 ( .Y(n5396), .A0(n3406), .A1(s_exp_diff_3_) );
  inv01 U3148 ( .Y(n5430), .A(opa_i[19]) );
  inv01 U3149 ( .Y(n5435), .A(opa_i[18]) );
  inv01 U3150 ( .Y(n5436), .A(opa_i[17]) );
  inv01 U3151 ( .Y(n5438), .A(n5439) );
  inv01 U3152 ( .Y(n5314), .A(n5201) );
  inv01 U3153 ( .Y(n5437), .A(n5349) );
  inv01 U3154 ( .Y(n5441), .A(opa_i[16]) );
  inv01 U3155 ( .Y(n5442), .A(opa_i[15]) );
  inv01 U3156 ( .Y(n5443), .A(opa_i[14]) );
  nand02 U3157 ( .Y(n5431), .A0(n5192), .A1(n5223) );
  inv01 U3158 ( .Y(n5444), .A(opa_i[13]) );
  inv01 U3159 ( .Y(n5445), .A(opa_i[12]) );
  inv01 U3160 ( .Y(n5446), .A(opa_i[11]) );
  ao22 U3161 ( .Y(n5447), .A0(n5216), .A1(n5394), .B0(n5218), .B1(n5391) );
  inv01 U3162 ( .Y(n5448), .A(opa_i[10]) );
  ao22 U3163 ( .Y(n5449), .A0(n5218), .A1(n5369), .B0(n5216), .B1(n5362) );
  inv01 U3164 ( .Y(n5297), .A(n5196) );
  inv01 U3165 ( .Y(n5451), .A(opa_i[9]) );
  ao22 U3166 ( .Y(n5452), .A0(n5365), .A1(n5379), .B0(n5217), .B1(n5378) );
  inv01 U3167 ( .Y(n5453), .A(opa_i[8]) );
  ao22 U3168 ( .Y(n5454), .A0(n5218), .A1(n5386), .B0(n5216), .B1(n5382) );
  inv01 U3169 ( .Y(n5456), .A(opa_i[7]) );
  inv01 U3170 ( .Y(n5457), .A(n5458) );
  inv01 U3171 ( .Y(n5312), .A(n5199) );
  and02 U3172 ( .Y(n5370), .A0(n5212), .A1(n5197) );
  nand02 U3173 ( .Y(n5330), .A0(n5418), .A1(n5288) );
  and02 U3174 ( .Y(n5360), .A0(n5460), .A1(n5461) );
  and02 U3175 ( .Y(n5368), .A0(n5209), .A1(n5192) );
  and02 U3176 ( .Y(n5338), .A0(n5192), .A1(n5212) );
  inv01 U3177 ( .Y(n5463), .A(n5351) );
  nor02 U3178 ( .Y(n5415), .A0(n5433), .A1(s_exp_diff_3_) );
  nor02 U3179 ( .Y(n5413), .A0(s_exp_diff_3_), .A1(s_exp_diff_2_) );
  and02 U3180 ( .Y(n5397), .A0(s_exp_diff_4_), .A1(n5409) );
  inv01 U3181 ( .Y(n5409), .A(n5464) );
  nand02 U3182 ( .Y(n5424), .A0(s_exp_diff_1_), .A1(s_exp_diff_0_) );
  nand02 U3183 ( .Y(n5450), .A0(n5465), .A1(n5466) );
  nand02 U3184 ( .Y(n5417), .A0(s_exp_diff_0_), .A1(n5465) );
  inv01 U3185 ( .Y(n5465), .A(s_exp_diff_1_) );
  nand02 U3186 ( .Y(n5416), .A0(s_exp_diff_1_), .A1(n5466) );
  inv01 U3187 ( .Y(n5466), .A(s_exp_diff_0_) );
  and02 U3188 ( .Y(n5363), .A0(n5019), .A1(n5192) );
  nand03 U3189 ( .Y(n5464), .A0(n5486), .A1(n5487), .A2(n5485) );
  nand03 U3190 ( .Y(n5279), .A0(n5199), .A1(n5289), .A2(n4907) );
  and02 U3191 ( .Y(n5298), .A0(n5291), .A1(n5156) );
  and03 U3192 ( .Y(n5291), .A0(n5162), .A1(n3943), .A2(n5194) );
  and03 U3193 ( .Y(n5310), .A0(n5188), .A1(n4043), .A2(n5166) );
  and03 U3194 ( .Y(n5285), .A0(n5182), .A1(n5158), .A2(n4047) );
  and03 U3195 ( .Y(n5304), .A0(n5186), .A1(n5160), .A2(n4217) );
  and03 U3196 ( .Y(n5293), .A0(n5190), .A1(n5164), .A2(n4045) );
  nand03 U3197 ( .Y(n5268), .A0(n5154), .A1(n5201), .A2(n5284) );
  inv01 U3198 ( .Y(n5324), .A(opb_i[1]) );
  inv01 U3199 ( .Y(n5403), .A(opa_i[1]) );
  ao21 U3200 ( .Y(U403_U6_Z_7), .A0(n____return498_7_), .A1(n5470), .B0(n3388)
         );
  oai22 U3201 ( .Y(n5471), .A0(n4924), .A1(n5206), .B0(n4943), .B1(n5207) );
  ao21 U3202 ( .Y(U403_U6_Z_6), .A0(n____return498_6_), .A1(n5470), .B0(n3385)
         );
  oai22 U3203 ( .Y(n5474), .A0(n4909), .A1(n5206), .B0(n4937), .B1(n5207) );
  ao21 U3204 ( .Y(U403_U6_Z_5), .A0(n____return498_5_), .A1(n5470), .B0(n3390)
         );
  oai22 U3205 ( .Y(n5475), .A0(n4918), .A1(n5206), .B0(n4933), .B1(n5207) );
  ao21 U3206 ( .Y(U403_U6_Z_4), .A0(n____return498_4_), .A1(n5470), .B0(n3387)
         );
  oai22 U3207 ( .Y(n5476), .A0(n4927), .A1(n5206), .B0(n4941), .B1(n5207) );
  ao21 U3208 ( .Y(U403_U6_Z_3), .A0(n____return498_3_), .A1(n5470), .B0(n3384)
         );
  oai22 U3209 ( .Y(n5477), .A0(n4912), .A1(n5206), .B0(n4935), .B1(n5207) );
  ao21 U3210 ( .Y(U403_U6_Z_2), .A0(n____return498_2_), .A1(n5470), .B0(n3389)
         );
  oai22 U3211 ( .Y(n5478), .A0(n4921), .A1(n5206), .B0(n4939), .B1(n5207) );
  ao21 U3212 ( .Y(U403_U6_Z_1), .A0(n____return498_1_), .A1(n5470), .B0(n3386)
         );
  oai22 U3213 ( .Y(n5479), .A0(n4915), .A1(n5206), .B0(n4931), .B1(n5207) );
  ao21 U3214 ( .Y(U403_U6_Z_0), .A0(n____return498_0_), .A1(n5470), .B0(n5480)
         );
  nand02 U3215 ( .Y(n5473), .A0(n4905), .A1(n5222) );
  nand02 U3216 ( .Y(n5472), .A0(n4905), .A1(n____return128) );
  inv01 U3217 ( .Y(n5425), .A(n5467) );
  inv01 U3218 ( .Y(n5329), .A(n5468) );
  nand02 U3219 ( .Y(n5468), .A0(n5481), .A1(n5482) );
  nand02 U3220 ( .Y(n5467), .A0(n5483), .A1(n5484) );
  pre_norm_addsub_DW01_cmp2_8_1 gt_162_gt_gt ( .A({1'b0, 1'b0, 1'b0, 
        s_rzeros_4_, s_rzeros_3_, s_rzeros_2_, s_rzeros_1_, s_rzeros_0_}), .B(
        {s_exp_diff_7_, s_exp_diff_6_, s_exp_diff_5_, s_exp_diff_4_, 
        s_exp_diff_3_, s_exp_diff_2_, s_exp_diff_1_, s_exp_diff_0_}), .LEQ(
        1'b0), .TC(1'b0), .LT_LE(n____return2686) );
  pre_norm_addsub_DW01_sub_8_0 r38 ( .A({U403_U5_Z_7, U403_U5_Z_6, U403_U5_Z_5, 
        U403_U5_Z_4, U403_U5_Z_3, U403_U5_Z_2, U403_U5_Z_1, U403_U5_Z_0}), .B(
        {U403_U6_Z_7, U403_U6_Z_6, U403_U6_Z_5, U403_U6_Z_4, U403_U6_Z_3, 
        U403_U6_Z_2, U403_U6_Z_1, U403_U6_Z_0}), .CI(1'b0), .DIFF({
        s_exp_diff436_7_, s_exp_diff436_6_, s_exp_diff436_5_, s_exp_diff436_4_, 
        s_exp_diff436_3_, s_exp_diff436_2_, s_exp_diff436_1_, s_exp_diff436_0_}) );
  pre_norm_addsub_DW01_inc_8_0 r510 ( .A({U403_U4_Z_7, U403_U4_Z_6, 
        U403_U4_Z_5, U403_U4_Z_4, U403_U4_Z_3, U403_U4_Z_2, U403_U4_Z_1, 
        U403_U4_Z_0}), .SUM({n____return498_7_, n____return498_6_, 
        n____return498_5_, n____return498_4_, n____return498_3_, 
        n____return498_2_, n____return498_1_, n____return498_0_}) );
  pre_norm_addsub_DW01_cmp2_8_0 gt_110_gt_gt ( .A(opb_i[30:23]), .B(
        opa_i[30:23]), .LEQ(1'b0), .TC(1'b0), .LT_LE(n____return128) );
endmodule


module addsub_28_DW01_addsub_28_0 ( A, B, CI, ADD_SUB, SUM, CO );
  input [27:0] A;
  input [27:0] B;
  output [27:0] SUM;
  input CI, ADD_SUB;
  output CO;
  wire   carry_27_, carry_26_, carry_25_, carry_24_, carry_23_, carry_22_,
         carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, carry_6_, carry_5_, carry_4_, carry_3_,
         carry_2_, carry_1_, n763, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762;

  buf02 U4 ( .Y(SUM[27]), .A(n763) );
  inv01 U5 ( .Y(SUM[26]), .A(n2) );
  inv02 U6 ( .Y(carry_27_), .A(n3) );
  inv02 U7 ( .Y(n4), .A(n713) );
  inv02 U8 ( .Y(n5), .A(A[26]) );
  inv02 U9 ( .Y(n6), .A(carry_26_) );
  nor02 U10 ( .Y(n7), .A0(n4), .A1(n8) );
  nor02 U11 ( .Y(n9), .A0(n5), .A1(n10) );
  nor02 U12 ( .Y(n11), .A0(n6), .A1(n12) );
  nor02 U13 ( .Y(n13), .A0(n6), .A1(n14) );
  nor02 U14 ( .Y(n2), .A0(n15), .A1(n16) );
  nor02 U15 ( .Y(n17), .A0(n5), .A1(n6) );
  nor02 U16 ( .Y(n18), .A0(n4), .A1(n6) );
  nor02 U17 ( .Y(n19), .A0(n4), .A1(n5) );
  nor02 U18 ( .Y(n3), .A0(n19), .A1(n20) );
  nor02 U19 ( .Y(n21), .A0(A[26]), .A1(carry_26_) );
  inv01 U20 ( .Y(n8), .A(n21) );
  nor02 U21 ( .Y(n22), .A0(n713), .A1(carry_26_) );
  inv01 U22 ( .Y(n10), .A(n22) );
  nor02 U23 ( .Y(n23), .A0(n713), .A1(A[26]) );
  inv01 U24 ( .Y(n12), .A(n23) );
  nor02 U25 ( .Y(n24), .A0(n4), .A1(n5) );
  inv01 U26 ( .Y(n14), .A(n24) );
  nor02 U27 ( .Y(n25), .A0(n7), .A1(n9) );
  inv01 U28 ( .Y(n15), .A(n25) );
  nor02 U29 ( .Y(n26), .A0(n11), .A1(n13) );
  inv01 U30 ( .Y(n16), .A(n26) );
  nor02 U31 ( .Y(n27), .A0(n17), .A1(n18) );
  inv01 U32 ( .Y(n20), .A(n27) );
  inv01 U33 ( .Y(SUM[25]), .A(n28) );
  inv02 U34 ( .Y(carry_26_), .A(n29) );
  inv02 U35 ( .Y(n30), .A(n721) );
  inv02 U36 ( .Y(n31), .A(A[25]) );
  inv02 U37 ( .Y(n32), .A(carry_25_) );
  nor02 U38 ( .Y(n33), .A0(n30), .A1(n34) );
  nor02 U39 ( .Y(n35), .A0(n31), .A1(n36) );
  nor02 U40 ( .Y(n37), .A0(n32), .A1(n38) );
  nor02 U41 ( .Y(n39), .A0(n32), .A1(n40) );
  nor02 U42 ( .Y(n28), .A0(n41), .A1(n42) );
  nor02 U43 ( .Y(n43), .A0(n31), .A1(n32) );
  nor02 U44 ( .Y(n44), .A0(n30), .A1(n32) );
  nor02 U45 ( .Y(n45), .A0(n30), .A1(n31) );
  nor02 U46 ( .Y(n29), .A0(n45), .A1(n46) );
  nor02 U47 ( .Y(n47), .A0(A[25]), .A1(carry_25_) );
  inv01 U48 ( .Y(n34), .A(n47) );
  nor02 U49 ( .Y(n48), .A0(n721), .A1(carry_25_) );
  inv01 U50 ( .Y(n36), .A(n48) );
  nor02 U51 ( .Y(n49), .A0(n721), .A1(A[25]) );
  inv01 U52 ( .Y(n38), .A(n49) );
  nor02 U53 ( .Y(n50), .A0(n30), .A1(n31) );
  inv01 U54 ( .Y(n40), .A(n50) );
  nor02 U55 ( .Y(n51), .A0(n33), .A1(n35) );
  inv01 U56 ( .Y(n41), .A(n51) );
  nor02 U57 ( .Y(n52), .A0(n37), .A1(n39) );
  inv01 U58 ( .Y(n42), .A(n52) );
  nor02 U59 ( .Y(n53), .A0(n43), .A1(n44) );
  inv01 U60 ( .Y(n46), .A(n53) );
  inv01 U61 ( .Y(SUM[24]), .A(n54) );
  inv02 U62 ( .Y(carry_25_), .A(n55) );
  inv02 U63 ( .Y(n56), .A(n759) );
  inv02 U64 ( .Y(n57), .A(A[24]) );
  inv02 U65 ( .Y(n58), .A(carry_24_) );
  nor02 U66 ( .Y(n59), .A0(n56), .A1(n60) );
  nor02 U67 ( .Y(n61), .A0(n57), .A1(n62) );
  nor02 U68 ( .Y(n63), .A0(n58), .A1(n64) );
  nor02 U69 ( .Y(n65), .A0(n58), .A1(n66) );
  nor02 U70 ( .Y(n54), .A0(n67), .A1(n68) );
  nor02 U71 ( .Y(n69), .A0(n57), .A1(n58) );
  nor02 U72 ( .Y(n70), .A0(n56), .A1(n58) );
  nor02 U73 ( .Y(n71), .A0(n56), .A1(n57) );
  nor02 U74 ( .Y(n55), .A0(n71), .A1(n72) );
  nor02 U75 ( .Y(n73), .A0(A[24]), .A1(carry_24_) );
  inv01 U76 ( .Y(n60), .A(n73) );
  nor02 U77 ( .Y(n74), .A0(n759), .A1(carry_24_) );
  inv01 U78 ( .Y(n62), .A(n74) );
  nor02 U79 ( .Y(n75), .A0(n759), .A1(A[24]) );
  inv01 U80 ( .Y(n64), .A(n75) );
  nor02 U81 ( .Y(n76), .A0(n56), .A1(n57) );
  inv01 U82 ( .Y(n66), .A(n76) );
  nor02 U83 ( .Y(n77), .A0(n59), .A1(n61) );
  inv01 U84 ( .Y(n67), .A(n77) );
  nor02 U85 ( .Y(n78), .A0(n63), .A1(n65) );
  inv01 U86 ( .Y(n68), .A(n78) );
  nor02 U87 ( .Y(n79), .A0(n69), .A1(n70) );
  inv01 U88 ( .Y(n72), .A(n79) );
  inv02 U89 ( .Y(SUM[23]), .A(n80) );
  inv02 U90 ( .Y(carry_24_), .A(n81) );
  inv02 U91 ( .Y(n82), .A(n729) );
  inv02 U92 ( .Y(n83), .A(A[23]) );
  inv02 U93 ( .Y(n84), .A(carry_23_) );
  nor02 U94 ( .Y(n85), .A0(n82), .A1(n86) );
  nor02 U95 ( .Y(n87), .A0(n83), .A1(n88) );
  nor02 U96 ( .Y(n89), .A0(n84), .A1(n90) );
  nor02 U97 ( .Y(n91), .A0(n84), .A1(n92) );
  nor02 U98 ( .Y(n80), .A0(n93), .A1(n94) );
  nor02 U99 ( .Y(n95), .A0(n83), .A1(n84) );
  nor02 U100 ( .Y(n96), .A0(n82), .A1(n84) );
  nor02 U101 ( .Y(n97), .A0(n82), .A1(n83) );
  nor02 U102 ( .Y(n81), .A0(n97), .A1(n98) );
  nor02 U103 ( .Y(n99), .A0(A[23]), .A1(carry_23_) );
  inv01 U104 ( .Y(n86), .A(n99) );
  nor02 U105 ( .Y(n100), .A0(n729), .A1(carry_23_) );
  inv01 U106 ( .Y(n88), .A(n100) );
  nor02 U107 ( .Y(n101), .A0(n729), .A1(A[23]) );
  inv01 U108 ( .Y(n90), .A(n101) );
  nor02 U109 ( .Y(n102), .A0(n82), .A1(n83) );
  inv01 U110 ( .Y(n92), .A(n102) );
  nor02 U111 ( .Y(n103), .A0(n85), .A1(n87) );
  inv01 U112 ( .Y(n93), .A(n103) );
  nor02 U113 ( .Y(n104), .A0(n89), .A1(n91) );
  inv02 U114 ( .Y(n94), .A(n104) );
  nor02 U115 ( .Y(n105), .A0(n95), .A1(n96) );
  inv01 U116 ( .Y(n98), .A(n105) );
  inv01 U117 ( .Y(SUM[1]), .A(n106) );
  inv02 U118 ( .Y(carry_2_), .A(n107) );
  inv02 U119 ( .Y(n108), .A(n705) );
  inv02 U120 ( .Y(n109), .A(A[1]) );
  inv02 U121 ( .Y(n110), .A(carry_1_) );
  nor02 U122 ( .Y(n111), .A0(n108), .A1(n112) );
  nor02 U123 ( .Y(n113), .A0(n109), .A1(n114) );
  nor02 U124 ( .Y(n115), .A0(n110), .A1(n116) );
  nor02 U125 ( .Y(n117), .A0(n110), .A1(n118) );
  nor02 U126 ( .Y(n106), .A0(n119), .A1(n120) );
  nor02 U127 ( .Y(n121), .A0(n109), .A1(n110) );
  nor02 U128 ( .Y(n122), .A0(n108), .A1(n110) );
  nor02 U129 ( .Y(n123), .A0(n108), .A1(n109) );
  nor02 U130 ( .Y(n107), .A0(n123), .A1(n124) );
  nor02 U131 ( .Y(n125), .A0(A[1]), .A1(carry_1_) );
  inv01 U132 ( .Y(n112), .A(n125) );
  nor02 U133 ( .Y(n126), .A0(n705), .A1(carry_1_) );
  inv01 U134 ( .Y(n114), .A(n126) );
  nor02 U135 ( .Y(n127), .A0(n705), .A1(A[1]) );
  inv01 U136 ( .Y(n116), .A(n127) );
  nor02 U137 ( .Y(n128), .A0(n108), .A1(n109) );
  inv01 U138 ( .Y(n118), .A(n128) );
  nor02 U139 ( .Y(n129), .A0(n111), .A1(n113) );
  inv01 U140 ( .Y(n119), .A(n129) );
  nor02 U141 ( .Y(n130), .A0(n115), .A1(n117) );
  inv01 U142 ( .Y(n120), .A(n130) );
  nor02 U143 ( .Y(n131), .A0(n121), .A1(n122) );
  inv01 U144 ( .Y(n124), .A(n131) );
  inv01 U145 ( .Y(SUM[2]), .A(n132) );
  inv02 U146 ( .Y(carry_3_), .A(n133) );
  inv02 U147 ( .Y(n134), .A(n757) );
  inv02 U148 ( .Y(n135), .A(A[2]) );
  inv02 U149 ( .Y(n136), .A(carry_2_) );
  nor02 U150 ( .Y(n137), .A0(n134), .A1(n138) );
  nor02 U151 ( .Y(n139), .A0(n135), .A1(n140) );
  nor02 U152 ( .Y(n141), .A0(n136), .A1(n142) );
  nor02 U153 ( .Y(n143), .A0(n136), .A1(n144) );
  nor02 U154 ( .Y(n132), .A0(n145), .A1(n146) );
  nor02 U155 ( .Y(n147), .A0(n135), .A1(n136) );
  nor02 U156 ( .Y(n148), .A0(n134), .A1(n136) );
  nor02 U157 ( .Y(n149), .A0(n134), .A1(n135) );
  nor02 U158 ( .Y(n133), .A0(n149), .A1(n150) );
  nor02 U159 ( .Y(n151), .A0(A[2]), .A1(carry_2_) );
  inv01 U160 ( .Y(n138), .A(n151) );
  nor02 U161 ( .Y(n152), .A0(n757), .A1(carry_2_) );
  inv01 U162 ( .Y(n140), .A(n152) );
  nor02 U163 ( .Y(n153), .A0(n757), .A1(A[2]) );
  inv01 U164 ( .Y(n142), .A(n153) );
  nor02 U165 ( .Y(n154), .A0(n134), .A1(n135) );
  inv01 U166 ( .Y(n144), .A(n154) );
  nor02 U167 ( .Y(n155), .A0(n137), .A1(n139) );
  inv01 U168 ( .Y(n145), .A(n155) );
  nor02 U169 ( .Y(n156), .A0(n141), .A1(n143) );
  inv01 U170 ( .Y(n146), .A(n156) );
  nor02 U171 ( .Y(n157), .A0(n147), .A1(n148) );
  inv01 U172 ( .Y(n150), .A(n157) );
  inv01 U173 ( .Y(SUM[3]), .A(n158) );
  inv02 U174 ( .Y(carry_4_), .A(n159) );
  inv02 U175 ( .Y(n160), .A(n737) );
  inv02 U176 ( .Y(n161), .A(A[3]) );
  inv02 U177 ( .Y(n162), .A(carry_3_) );
  nor02 U178 ( .Y(n163), .A0(n160), .A1(n164) );
  nor02 U179 ( .Y(n165), .A0(n161), .A1(n166) );
  nor02 U180 ( .Y(n167), .A0(n162), .A1(n168) );
  nor02 U181 ( .Y(n169), .A0(n162), .A1(n170) );
  nor02 U182 ( .Y(n158), .A0(n171), .A1(n172) );
  nor02 U183 ( .Y(n173), .A0(n161), .A1(n162) );
  nor02 U184 ( .Y(n174), .A0(n160), .A1(n162) );
  nor02 U185 ( .Y(n175), .A0(n160), .A1(n161) );
  nor02 U186 ( .Y(n159), .A0(n175), .A1(n176) );
  nor02 U187 ( .Y(n177), .A0(A[3]), .A1(carry_3_) );
  inv01 U188 ( .Y(n164), .A(n177) );
  nor02 U189 ( .Y(n178), .A0(n737), .A1(carry_3_) );
  inv01 U190 ( .Y(n166), .A(n178) );
  nor02 U191 ( .Y(n179), .A0(n737), .A1(A[3]) );
  inv01 U192 ( .Y(n168), .A(n179) );
  nor02 U193 ( .Y(n180), .A0(n160), .A1(n161) );
  inv01 U194 ( .Y(n170), .A(n180) );
  nor02 U195 ( .Y(n181), .A0(n163), .A1(n165) );
  inv01 U196 ( .Y(n171), .A(n181) );
  nor02 U197 ( .Y(n182), .A0(n167), .A1(n169) );
  inv01 U198 ( .Y(n172), .A(n182) );
  nor02 U199 ( .Y(n183), .A0(n173), .A1(n174) );
  inv01 U200 ( .Y(n176), .A(n183) );
  inv01 U201 ( .Y(SUM[4]), .A(n184) );
  inv02 U202 ( .Y(carry_5_), .A(n185) );
  inv02 U203 ( .Y(n186), .A(n739) );
  inv02 U204 ( .Y(n187), .A(A[4]) );
  inv02 U205 ( .Y(n188), .A(carry_4_) );
  nor02 U206 ( .Y(n189), .A0(n186), .A1(n190) );
  nor02 U207 ( .Y(n191), .A0(n187), .A1(n192) );
  nor02 U208 ( .Y(n193), .A0(n188), .A1(n194) );
  nor02 U209 ( .Y(n195), .A0(n188), .A1(n196) );
  nor02 U210 ( .Y(n184), .A0(n197), .A1(n198) );
  nor02 U211 ( .Y(n199), .A0(n187), .A1(n188) );
  nor02 U212 ( .Y(n200), .A0(n186), .A1(n188) );
  nor02 U213 ( .Y(n201), .A0(n186), .A1(n187) );
  nor02 U214 ( .Y(n185), .A0(n201), .A1(n202) );
  nor02 U215 ( .Y(n203), .A0(A[4]), .A1(carry_4_) );
  inv01 U216 ( .Y(n190), .A(n203) );
  nor02 U217 ( .Y(n204), .A0(n739), .A1(carry_4_) );
  inv01 U218 ( .Y(n192), .A(n204) );
  nor02 U219 ( .Y(n205), .A0(n739), .A1(A[4]) );
  inv01 U220 ( .Y(n194), .A(n205) );
  nor02 U221 ( .Y(n206), .A0(n186), .A1(n187) );
  inv01 U222 ( .Y(n196), .A(n206) );
  nor02 U223 ( .Y(n207), .A0(n189), .A1(n191) );
  inv01 U224 ( .Y(n197), .A(n207) );
  nor02 U225 ( .Y(n208), .A0(n193), .A1(n195) );
  inv01 U226 ( .Y(n198), .A(n208) );
  nor02 U227 ( .Y(n209), .A0(n199), .A1(n200) );
  inv01 U228 ( .Y(n202), .A(n209) );
  inv01 U229 ( .Y(SUM[5]), .A(n210) );
  inv02 U230 ( .Y(carry_6_), .A(n211) );
  inv02 U231 ( .Y(n212), .A(n719) );
  inv02 U232 ( .Y(n213), .A(A[5]) );
  inv02 U233 ( .Y(n214), .A(carry_5_) );
  nor02 U234 ( .Y(n215), .A0(n212), .A1(n216) );
  nor02 U235 ( .Y(n217), .A0(n213), .A1(n218) );
  nor02 U236 ( .Y(n219), .A0(n214), .A1(n220) );
  nor02 U237 ( .Y(n221), .A0(n214), .A1(n222) );
  nor02 U238 ( .Y(n210), .A0(n223), .A1(n224) );
  nor02 U239 ( .Y(n225), .A0(n213), .A1(n214) );
  nor02 U240 ( .Y(n226), .A0(n212), .A1(n214) );
  nor02 U241 ( .Y(n227), .A0(n212), .A1(n213) );
  nor02 U242 ( .Y(n211), .A0(n227), .A1(n228) );
  nor02 U243 ( .Y(n229), .A0(A[5]), .A1(carry_5_) );
  inv01 U244 ( .Y(n216), .A(n229) );
  nor02 U245 ( .Y(n230), .A0(n719), .A1(carry_5_) );
  inv01 U246 ( .Y(n218), .A(n230) );
  nor02 U247 ( .Y(n231), .A0(n719), .A1(A[5]) );
  inv01 U248 ( .Y(n220), .A(n231) );
  nor02 U249 ( .Y(n232), .A0(n212), .A1(n213) );
  inv01 U250 ( .Y(n222), .A(n232) );
  nor02 U251 ( .Y(n233), .A0(n215), .A1(n217) );
  inv01 U252 ( .Y(n223), .A(n233) );
  nor02 U253 ( .Y(n234), .A0(n219), .A1(n221) );
  inv01 U254 ( .Y(n224), .A(n234) );
  nor02 U255 ( .Y(n235), .A0(n225), .A1(n226) );
  inv01 U256 ( .Y(n228), .A(n235) );
  inv01 U257 ( .Y(SUM[6]), .A(n236) );
  inv02 U258 ( .Y(carry_7_), .A(n237) );
  inv02 U259 ( .Y(n238), .A(n745) );
  inv02 U260 ( .Y(n239), .A(A[6]) );
  inv02 U261 ( .Y(n240), .A(carry_6_) );
  nor02 U262 ( .Y(n241), .A0(n238), .A1(n242) );
  nor02 U263 ( .Y(n243), .A0(n239), .A1(n244) );
  nor02 U264 ( .Y(n245), .A0(n240), .A1(n246) );
  nor02 U265 ( .Y(n247), .A0(n240), .A1(n248) );
  nor02 U266 ( .Y(n236), .A0(n249), .A1(n250) );
  nor02 U267 ( .Y(n251), .A0(n239), .A1(n240) );
  nor02 U268 ( .Y(n252), .A0(n238), .A1(n240) );
  nor02 U269 ( .Y(n253), .A0(n238), .A1(n239) );
  nor02 U270 ( .Y(n237), .A0(n253), .A1(n254) );
  nor02 U271 ( .Y(n255), .A0(A[6]), .A1(carry_6_) );
  inv01 U272 ( .Y(n242), .A(n255) );
  nor02 U273 ( .Y(n256), .A0(n745), .A1(carry_6_) );
  inv01 U274 ( .Y(n244), .A(n256) );
  nor02 U275 ( .Y(n257), .A0(n745), .A1(A[6]) );
  inv01 U276 ( .Y(n246), .A(n257) );
  nor02 U277 ( .Y(n258), .A0(n238), .A1(n239) );
  inv01 U278 ( .Y(n248), .A(n258) );
  nor02 U279 ( .Y(n259), .A0(n241), .A1(n243) );
  inv01 U280 ( .Y(n249), .A(n259) );
  nor02 U281 ( .Y(n260), .A0(n245), .A1(n247) );
  inv01 U282 ( .Y(n250), .A(n260) );
  nor02 U283 ( .Y(n261), .A0(n251), .A1(n252) );
  inv01 U284 ( .Y(n254), .A(n261) );
  inv01 U285 ( .Y(SUM[7]), .A(n262) );
  inv02 U286 ( .Y(carry_8_), .A(n263) );
  inv02 U287 ( .Y(n264), .A(n717) );
  inv02 U288 ( .Y(n265), .A(A[7]) );
  inv02 U289 ( .Y(n266), .A(carry_7_) );
  nor02 U290 ( .Y(n267), .A0(n264), .A1(n268) );
  nor02 U291 ( .Y(n269), .A0(n265), .A1(n270) );
  nor02 U292 ( .Y(n271), .A0(n266), .A1(n272) );
  nor02 U293 ( .Y(n273), .A0(n266), .A1(n274) );
  nor02 U294 ( .Y(n262), .A0(n275), .A1(n276) );
  nor02 U295 ( .Y(n277), .A0(n265), .A1(n266) );
  nor02 U296 ( .Y(n278), .A0(n264), .A1(n266) );
  nor02 U297 ( .Y(n279), .A0(n264), .A1(n265) );
  nor02 U298 ( .Y(n263), .A0(n279), .A1(n280) );
  nor02 U299 ( .Y(n281), .A0(A[7]), .A1(carry_7_) );
  inv01 U300 ( .Y(n268), .A(n281) );
  nor02 U301 ( .Y(n282), .A0(n717), .A1(carry_7_) );
  inv01 U302 ( .Y(n270), .A(n282) );
  nor02 U303 ( .Y(n283), .A0(n717), .A1(A[7]) );
  inv01 U304 ( .Y(n272), .A(n283) );
  nor02 U305 ( .Y(n284), .A0(n264), .A1(n265) );
  inv01 U306 ( .Y(n274), .A(n284) );
  nor02 U307 ( .Y(n285), .A0(n267), .A1(n269) );
  inv01 U308 ( .Y(n275), .A(n285) );
  nor02 U309 ( .Y(n286), .A0(n271), .A1(n273) );
  inv01 U310 ( .Y(n276), .A(n286) );
  nor02 U311 ( .Y(n287), .A0(n277), .A1(n278) );
  inv01 U312 ( .Y(n280), .A(n287) );
  inv01 U313 ( .Y(SUM[8]), .A(n288) );
  inv02 U314 ( .Y(carry_9_), .A(n289) );
  inv02 U315 ( .Y(n290), .A(n741) );
  inv02 U316 ( .Y(n291), .A(A[8]) );
  inv02 U317 ( .Y(n292), .A(carry_8_) );
  nor02 U318 ( .Y(n293), .A0(n290), .A1(n294) );
  nor02 U319 ( .Y(n295), .A0(n291), .A1(n296) );
  nor02 U320 ( .Y(n297), .A0(n292), .A1(n298) );
  nor02 U321 ( .Y(n299), .A0(n292), .A1(n300) );
  nor02 U322 ( .Y(n288), .A0(n301), .A1(n302) );
  nor02 U323 ( .Y(n303), .A0(n291), .A1(n292) );
  nor02 U324 ( .Y(n304), .A0(n290), .A1(n292) );
  nor02 U325 ( .Y(n305), .A0(n290), .A1(n291) );
  nor02 U326 ( .Y(n289), .A0(n305), .A1(n306) );
  nor02 U327 ( .Y(n307), .A0(A[8]), .A1(carry_8_) );
  inv01 U328 ( .Y(n294), .A(n307) );
  nor02 U329 ( .Y(n308), .A0(n741), .A1(carry_8_) );
  inv01 U330 ( .Y(n296), .A(n308) );
  nor02 U331 ( .Y(n309), .A0(n741), .A1(A[8]) );
  inv01 U332 ( .Y(n298), .A(n309) );
  nor02 U333 ( .Y(n310), .A0(n290), .A1(n291) );
  inv01 U334 ( .Y(n300), .A(n310) );
  nor02 U335 ( .Y(n311), .A0(n293), .A1(n295) );
  inv01 U336 ( .Y(n301), .A(n311) );
  nor02 U337 ( .Y(n312), .A0(n297), .A1(n299) );
  inv01 U338 ( .Y(n302), .A(n312) );
  nor02 U339 ( .Y(n313), .A0(n303), .A1(n304) );
  inv01 U340 ( .Y(n306), .A(n313) );
  inv01 U341 ( .Y(SUM[9]), .A(n314) );
  inv02 U342 ( .Y(carry_10_), .A(n315) );
  inv02 U343 ( .Y(n316), .A(n733) );
  inv02 U344 ( .Y(n317), .A(A[9]) );
  inv02 U345 ( .Y(n318), .A(carry_9_) );
  nor02 U346 ( .Y(n319), .A0(n316), .A1(n320) );
  nor02 U347 ( .Y(n321), .A0(n317), .A1(n322) );
  nor02 U348 ( .Y(n323), .A0(n318), .A1(n324) );
  nor02 U349 ( .Y(n325), .A0(n318), .A1(n326) );
  nor02 U350 ( .Y(n314), .A0(n327), .A1(n328) );
  nor02 U351 ( .Y(n329), .A0(n317), .A1(n318) );
  nor02 U352 ( .Y(n330), .A0(n316), .A1(n318) );
  nor02 U353 ( .Y(n331), .A0(n316), .A1(n317) );
  nor02 U354 ( .Y(n315), .A0(n331), .A1(n332) );
  nor02 U355 ( .Y(n333), .A0(A[9]), .A1(carry_9_) );
  inv01 U356 ( .Y(n320), .A(n333) );
  nor02 U357 ( .Y(n334), .A0(n733), .A1(carry_9_) );
  inv01 U358 ( .Y(n322), .A(n334) );
  nor02 U359 ( .Y(n335), .A0(n733), .A1(A[9]) );
  inv01 U360 ( .Y(n324), .A(n335) );
  nor02 U361 ( .Y(n336), .A0(n316), .A1(n317) );
  inv01 U362 ( .Y(n326), .A(n336) );
  nor02 U363 ( .Y(n337), .A0(n319), .A1(n321) );
  inv01 U364 ( .Y(n327), .A(n337) );
  nor02 U365 ( .Y(n338), .A0(n323), .A1(n325) );
  inv01 U366 ( .Y(n328), .A(n338) );
  nor02 U367 ( .Y(n339), .A0(n329), .A1(n330) );
  inv01 U368 ( .Y(n332), .A(n339) );
  inv02 U369 ( .Y(SUM[17]), .A(n340) );
  inv02 U370 ( .Y(carry_18_), .A(n341) );
  inv02 U371 ( .Y(n342), .A(n723) );
  inv02 U372 ( .Y(n343), .A(A[17]) );
  inv02 U373 ( .Y(n344), .A(carry_17_) );
  nor02 U374 ( .Y(n345), .A0(n342), .A1(n346) );
  nor02 U375 ( .Y(n347), .A0(n343), .A1(n348) );
  nor02 U376 ( .Y(n349), .A0(n344), .A1(n350) );
  nor02 U377 ( .Y(n351), .A0(n344), .A1(n352) );
  nor02 U378 ( .Y(n340), .A0(n353), .A1(n354) );
  nor02 U379 ( .Y(n355), .A0(n343), .A1(n344) );
  nor02 U380 ( .Y(n356), .A0(n342), .A1(n344) );
  nor02 U381 ( .Y(n357), .A0(n342), .A1(n343) );
  nor02 U382 ( .Y(n341), .A0(n357), .A1(n358) );
  nor02 U383 ( .Y(n359), .A0(A[17]), .A1(carry_17_) );
  inv01 U384 ( .Y(n346), .A(n359) );
  nor02 U385 ( .Y(n360), .A0(n723), .A1(carry_17_) );
  inv01 U386 ( .Y(n348), .A(n360) );
  nor02 U387 ( .Y(n361), .A0(n723), .A1(A[17]) );
  inv01 U388 ( .Y(n350), .A(n361) );
  nor02 U389 ( .Y(n362), .A0(n342), .A1(n343) );
  inv01 U390 ( .Y(n352), .A(n362) );
  nor02 U391 ( .Y(n363), .A0(n345), .A1(n347) );
  inv01 U392 ( .Y(n353), .A(n363) );
  nor02 U393 ( .Y(n364), .A0(n349), .A1(n351) );
  inv02 U394 ( .Y(n354), .A(n364) );
  nor02 U395 ( .Y(n365), .A0(n355), .A1(n356) );
  inv01 U396 ( .Y(n358), .A(n365) );
  inv02 U397 ( .Y(SUM[10]), .A(n366) );
  inv02 U398 ( .Y(carry_11_), .A(n367) );
  inv02 U399 ( .Y(n368), .A(n735) );
  inv02 U400 ( .Y(n369), .A(A[10]) );
  inv02 U401 ( .Y(n370), .A(carry_10_) );
  nor02 U402 ( .Y(n371), .A0(n368), .A1(n372) );
  nor02 U403 ( .Y(n373), .A0(n369), .A1(n374) );
  nor02 U404 ( .Y(n375), .A0(n370), .A1(n376) );
  nor02 U405 ( .Y(n377), .A0(n370), .A1(n378) );
  nor02 U406 ( .Y(n366), .A0(n379), .A1(n380) );
  nor02 U407 ( .Y(n381), .A0(n369), .A1(n370) );
  nor02 U408 ( .Y(n382), .A0(n368), .A1(n370) );
  nor02 U409 ( .Y(n383), .A0(n368), .A1(n369) );
  nor02 U410 ( .Y(n367), .A0(n383), .A1(n384) );
  nor02 U411 ( .Y(n385), .A0(A[10]), .A1(carry_10_) );
  inv01 U412 ( .Y(n372), .A(n385) );
  nor02 U413 ( .Y(n386), .A0(n735), .A1(carry_10_) );
  inv01 U414 ( .Y(n374), .A(n386) );
  nor02 U415 ( .Y(n387), .A0(n735), .A1(A[10]) );
  inv01 U416 ( .Y(n376), .A(n387) );
  nor02 U417 ( .Y(n388), .A0(n368), .A1(n369) );
  inv01 U418 ( .Y(n378), .A(n388) );
  nor02 U419 ( .Y(n389), .A0(n371), .A1(n373) );
  inv01 U420 ( .Y(n379), .A(n389) );
  nor02 U421 ( .Y(n390), .A0(n375), .A1(n377) );
  inv02 U422 ( .Y(n380), .A(n390) );
  nor02 U423 ( .Y(n391), .A0(n381), .A1(n382) );
  inv01 U424 ( .Y(n384), .A(n391) );
  inv01 U425 ( .Y(SUM[11]), .A(n392) );
  inv02 U426 ( .Y(carry_12_), .A(n393) );
  inv02 U427 ( .Y(n394), .A(n727) );
  inv02 U428 ( .Y(n395), .A(A[11]) );
  inv02 U429 ( .Y(n396), .A(carry_11_) );
  nor02 U430 ( .Y(n397), .A0(n394), .A1(n398) );
  nor02 U431 ( .Y(n399), .A0(n395), .A1(n400) );
  nor02 U432 ( .Y(n401), .A0(n396), .A1(n402) );
  nor02 U433 ( .Y(n403), .A0(n396), .A1(n404) );
  nor02 U434 ( .Y(n392), .A0(n405), .A1(n406) );
  nor02 U435 ( .Y(n407), .A0(n395), .A1(n396) );
  nor02 U436 ( .Y(n408), .A0(n394), .A1(n396) );
  nor02 U437 ( .Y(n409), .A0(n394), .A1(n395) );
  nor02 U438 ( .Y(n393), .A0(n409), .A1(n410) );
  nor02 U439 ( .Y(n411), .A0(A[11]), .A1(carry_11_) );
  inv01 U440 ( .Y(n398), .A(n411) );
  nor02 U441 ( .Y(n412), .A0(n727), .A1(carry_11_) );
  inv01 U442 ( .Y(n400), .A(n412) );
  nor02 U443 ( .Y(n413), .A0(n727), .A1(A[11]) );
  inv01 U444 ( .Y(n402), .A(n413) );
  nor02 U445 ( .Y(n414), .A0(n394), .A1(n395) );
  inv01 U446 ( .Y(n404), .A(n414) );
  nor02 U447 ( .Y(n415), .A0(n397), .A1(n399) );
  inv01 U448 ( .Y(n405), .A(n415) );
  nor02 U449 ( .Y(n416), .A0(n401), .A1(n403) );
  inv01 U450 ( .Y(n406), .A(n416) );
  nor02 U451 ( .Y(n417), .A0(n407), .A1(n408) );
  inv01 U452 ( .Y(n410), .A(n417) );
  inv01 U453 ( .Y(SUM[18]), .A(n418) );
  inv02 U454 ( .Y(carry_19_), .A(n419) );
  inv02 U455 ( .Y(n420), .A(n749) );
  inv02 U456 ( .Y(n421), .A(A[18]) );
  inv02 U457 ( .Y(n422), .A(carry_18_) );
  nor02 U458 ( .Y(n423), .A0(n420), .A1(n424) );
  nor02 U459 ( .Y(n425), .A0(n421), .A1(n426) );
  nor02 U460 ( .Y(n427), .A0(n422), .A1(n428) );
  nor02 U461 ( .Y(n429), .A0(n422), .A1(n430) );
  nor02 U462 ( .Y(n418), .A0(n431), .A1(n432) );
  nor02 U463 ( .Y(n433), .A0(n421), .A1(n422) );
  nor02 U464 ( .Y(n434), .A0(n420), .A1(n422) );
  nor02 U465 ( .Y(n435), .A0(n420), .A1(n421) );
  nor02 U466 ( .Y(n419), .A0(n435), .A1(n436) );
  nor02 U467 ( .Y(n437), .A0(A[18]), .A1(carry_18_) );
  inv01 U468 ( .Y(n424), .A(n437) );
  nor02 U469 ( .Y(n438), .A0(n749), .A1(carry_18_) );
  inv01 U470 ( .Y(n426), .A(n438) );
  nor02 U471 ( .Y(n439), .A0(n749), .A1(A[18]) );
  inv01 U472 ( .Y(n428), .A(n439) );
  nor02 U473 ( .Y(n440), .A0(n420), .A1(n421) );
  inv01 U474 ( .Y(n430), .A(n440) );
  nor02 U475 ( .Y(n441), .A0(n423), .A1(n425) );
  inv01 U476 ( .Y(n431), .A(n441) );
  nor02 U477 ( .Y(n442), .A0(n427), .A1(n429) );
  inv01 U478 ( .Y(n432), .A(n442) );
  nor02 U479 ( .Y(n443), .A0(n433), .A1(n434) );
  inv01 U480 ( .Y(n436), .A(n443) );
  inv01 U481 ( .Y(SUM[19]), .A(n444) );
  inv02 U482 ( .Y(carry_20_), .A(n445) );
  inv02 U483 ( .Y(n446), .A(n715) );
  inv02 U484 ( .Y(n447), .A(A[19]) );
  inv02 U485 ( .Y(n448), .A(carry_19_) );
  nor02 U486 ( .Y(n449), .A0(n446), .A1(n450) );
  nor02 U487 ( .Y(n451), .A0(n447), .A1(n452) );
  nor02 U488 ( .Y(n453), .A0(n448), .A1(n454) );
  nor02 U489 ( .Y(n455), .A0(n448), .A1(n456) );
  nor02 U490 ( .Y(n444), .A0(n457), .A1(n458) );
  nor02 U491 ( .Y(n459), .A0(n447), .A1(n448) );
  nor02 U492 ( .Y(n460), .A0(n446), .A1(n448) );
  nor02 U493 ( .Y(n461), .A0(n446), .A1(n447) );
  nor02 U494 ( .Y(n445), .A0(n461), .A1(n462) );
  nor02 U495 ( .Y(n463), .A0(A[19]), .A1(carry_19_) );
  inv01 U496 ( .Y(n450), .A(n463) );
  nor02 U497 ( .Y(n464), .A0(n715), .A1(carry_19_) );
  inv01 U498 ( .Y(n452), .A(n464) );
  nor02 U499 ( .Y(n465), .A0(n715), .A1(A[19]) );
  inv01 U500 ( .Y(n454), .A(n465) );
  nor02 U501 ( .Y(n466), .A0(n446), .A1(n447) );
  inv01 U502 ( .Y(n456), .A(n466) );
  nor02 U503 ( .Y(n467), .A0(n449), .A1(n451) );
  inv01 U504 ( .Y(n457), .A(n467) );
  nor02 U505 ( .Y(n468), .A0(n453), .A1(n455) );
  inv01 U506 ( .Y(n458), .A(n468) );
  nor02 U507 ( .Y(n469), .A0(n459), .A1(n460) );
  inv01 U508 ( .Y(n462), .A(n469) );
  inv01 U509 ( .Y(SUM[12]), .A(n470) );
  inv02 U510 ( .Y(carry_13_), .A(n471) );
  inv02 U511 ( .Y(n472), .A(n731) );
  inv02 U512 ( .Y(n473), .A(A[12]) );
  inv02 U513 ( .Y(n474), .A(carry_12_) );
  nor02 U514 ( .Y(n475), .A0(n472), .A1(n476) );
  nor02 U515 ( .Y(n477), .A0(n473), .A1(n478) );
  nor02 U516 ( .Y(n479), .A0(n474), .A1(n480) );
  nor02 U517 ( .Y(n481), .A0(n474), .A1(n482) );
  nor02 U518 ( .Y(n470), .A0(n483), .A1(n484) );
  nor02 U519 ( .Y(n485), .A0(n473), .A1(n474) );
  nor02 U520 ( .Y(n486), .A0(n472), .A1(n474) );
  nor02 U521 ( .Y(n487), .A0(n472), .A1(n473) );
  nor02 U522 ( .Y(n471), .A0(n487), .A1(n488) );
  nor02 U523 ( .Y(n489), .A0(A[12]), .A1(carry_12_) );
  inv01 U524 ( .Y(n476), .A(n489) );
  nor02 U525 ( .Y(n490), .A0(n731), .A1(carry_12_) );
  inv01 U526 ( .Y(n478), .A(n490) );
  nor02 U527 ( .Y(n491), .A0(n731), .A1(A[12]) );
  inv01 U528 ( .Y(n480), .A(n491) );
  nor02 U529 ( .Y(n492), .A0(n472), .A1(n473) );
  inv01 U530 ( .Y(n482), .A(n492) );
  nor02 U531 ( .Y(n493), .A0(n475), .A1(n477) );
  inv01 U532 ( .Y(n483), .A(n493) );
  nor02 U533 ( .Y(n494), .A0(n479), .A1(n481) );
  inv01 U534 ( .Y(n484), .A(n494) );
  nor02 U535 ( .Y(n495), .A0(n485), .A1(n486) );
  inv01 U536 ( .Y(n488), .A(n495) );
  inv01 U537 ( .Y(SUM[13]), .A(n496) );
  inv02 U538 ( .Y(carry_14_), .A(n497) );
  inv02 U539 ( .Y(n498), .A(n707) );
  inv02 U540 ( .Y(n499), .A(A[13]) );
  inv02 U541 ( .Y(n500), .A(carry_13_) );
  nor02 U542 ( .Y(n501), .A0(n498), .A1(n502) );
  nor02 U543 ( .Y(n503), .A0(n499), .A1(n504) );
  nor02 U544 ( .Y(n505), .A0(n500), .A1(n506) );
  nor02 U545 ( .Y(n507), .A0(n500), .A1(n508) );
  nor02 U546 ( .Y(n496), .A0(n509), .A1(n510) );
  nor02 U547 ( .Y(n511), .A0(n499), .A1(n500) );
  nor02 U548 ( .Y(n512), .A0(n498), .A1(n500) );
  nor02 U549 ( .Y(n513), .A0(n498), .A1(n499) );
  nor02 U550 ( .Y(n497), .A0(n513), .A1(n514) );
  nor02 U551 ( .Y(n515), .A0(A[13]), .A1(carry_13_) );
  inv01 U552 ( .Y(n502), .A(n515) );
  nor02 U553 ( .Y(n516), .A0(n707), .A1(carry_13_) );
  inv01 U554 ( .Y(n504), .A(n516) );
  nor02 U555 ( .Y(n517), .A0(n707), .A1(A[13]) );
  inv01 U556 ( .Y(n506), .A(n517) );
  nor02 U557 ( .Y(n518), .A0(n498), .A1(n499) );
  inv01 U558 ( .Y(n508), .A(n518) );
  nor02 U559 ( .Y(n519), .A0(n501), .A1(n503) );
  inv01 U560 ( .Y(n509), .A(n519) );
  nor02 U561 ( .Y(n520), .A0(n505), .A1(n507) );
  inv01 U562 ( .Y(n510), .A(n520) );
  nor02 U563 ( .Y(n521), .A0(n511), .A1(n512) );
  inv01 U564 ( .Y(n514), .A(n521) );
  inv01 U565 ( .Y(SUM[20]), .A(n522) );
  inv02 U566 ( .Y(carry_21_), .A(n523) );
  inv02 U567 ( .Y(n524), .A(n753) );
  inv02 U568 ( .Y(n525), .A(A[20]) );
  inv02 U569 ( .Y(n526), .A(carry_20_) );
  nor02 U570 ( .Y(n527), .A0(n524), .A1(n528) );
  nor02 U571 ( .Y(n529), .A0(n525), .A1(n530) );
  nor02 U572 ( .Y(n531), .A0(n526), .A1(n532) );
  nor02 U573 ( .Y(n533), .A0(n526), .A1(n534) );
  nor02 U574 ( .Y(n522), .A0(n535), .A1(n536) );
  nor02 U575 ( .Y(n537), .A0(n525), .A1(n526) );
  nor02 U576 ( .Y(n538), .A0(n524), .A1(n526) );
  nor02 U577 ( .Y(n539), .A0(n524), .A1(n525) );
  nor02 U578 ( .Y(n523), .A0(n539), .A1(n540) );
  nor02 U579 ( .Y(n541), .A0(A[20]), .A1(carry_20_) );
  inv01 U580 ( .Y(n528), .A(n541) );
  nor02 U581 ( .Y(n542), .A0(n753), .A1(carry_20_) );
  inv01 U582 ( .Y(n530), .A(n542) );
  nor02 U583 ( .Y(n543), .A0(n753), .A1(A[20]) );
  inv01 U584 ( .Y(n532), .A(n543) );
  nor02 U585 ( .Y(n544), .A0(n524), .A1(n525) );
  inv01 U586 ( .Y(n534), .A(n544) );
  nor02 U587 ( .Y(n545), .A0(n527), .A1(n529) );
  inv01 U588 ( .Y(n535), .A(n545) );
  nor02 U589 ( .Y(n546), .A0(n531), .A1(n533) );
  inv01 U590 ( .Y(n536), .A(n546) );
  nor02 U591 ( .Y(n547), .A0(n537), .A1(n538) );
  inv01 U592 ( .Y(n540), .A(n547) );
  inv02 U593 ( .Y(SUM[21]), .A(n548) );
  inv02 U594 ( .Y(carry_22_), .A(n549) );
  inv02 U595 ( .Y(n550), .A(n725) );
  inv02 U596 ( .Y(n551), .A(A[21]) );
  inv02 U597 ( .Y(n552), .A(carry_21_) );
  nor02 U598 ( .Y(n553), .A0(n550), .A1(n554) );
  nor02 U599 ( .Y(n555), .A0(n551), .A1(n556) );
  nor02 U600 ( .Y(n557), .A0(n552), .A1(n558) );
  nor02 U601 ( .Y(n559), .A0(n552), .A1(n560) );
  nor02 U602 ( .Y(n548), .A0(n561), .A1(n562) );
  nor02 U603 ( .Y(n563), .A0(n551), .A1(n552) );
  nor02 U604 ( .Y(n564), .A0(n550), .A1(n552) );
  nor02 U605 ( .Y(n565), .A0(n550), .A1(n551) );
  nor02 U606 ( .Y(n549), .A0(n565), .A1(n566) );
  nor02 U607 ( .Y(n567), .A0(A[21]), .A1(carry_21_) );
  inv01 U608 ( .Y(n554), .A(n567) );
  nor02 U609 ( .Y(n568), .A0(n725), .A1(carry_21_) );
  inv01 U610 ( .Y(n556), .A(n568) );
  nor02 U611 ( .Y(n569), .A0(n725), .A1(A[21]) );
  inv01 U612 ( .Y(n558), .A(n569) );
  nor02 U613 ( .Y(n570), .A0(n550), .A1(n551) );
  inv01 U614 ( .Y(n560), .A(n570) );
  nor02 U615 ( .Y(n571), .A0(n553), .A1(n555) );
  inv01 U616 ( .Y(n561), .A(n571) );
  nor02 U617 ( .Y(n572), .A0(n557), .A1(n559) );
  inv02 U618 ( .Y(n562), .A(n572) );
  nor02 U619 ( .Y(n573), .A0(n563), .A1(n564) );
  inv01 U620 ( .Y(n566), .A(n573) );
  inv01 U621 ( .Y(SUM[14]), .A(n574) );
  inv02 U622 ( .Y(carry_15_), .A(n575) );
  inv02 U623 ( .Y(n576), .A(n747) );
  inv02 U624 ( .Y(n577), .A(A[14]) );
  inv02 U625 ( .Y(n578), .A(carry_14_) );
  nor02 U626 ( .Y(n579), .A0(n576), .A1(n580) );
  nor02 U627 ( .Y(n581), .A0(n577), .A1(n582) );
  nor02 U628 ( .Y(n583), .A0(n578), .A1(n584) );
  nor02 U629 ( .Y(n585), .A0(n578), .A1(n586) );
  nor02 U630 ( .Y(n574), .A0(n587), .A1(n588) );
  nor02 U631 ( .Y(n589), .A0(n577), .A1(n578) );
  nor02 U632 ( .Y(n590), .A0(n576), .A1(n578) );
  nor02 U633 ( .Y(n591), .A0(n576), .A1(n577) );
  nor02 U634 ( .Y(n575), .A0(n591), .A1(n592) );
  nor02 U635 ( .Y(n593), .A0(A[14]), .A1(carry_14_) );
  inv01 U636 ( .Y(n580), .A(n593) );
  nor02 U637 ( .Y(n594), .A0(n747), .A1(carry_14_) );
  inv01 U638 ( .Y(n582), .A(n594) );
  nor02 U639 ( .Y(n595), .A0(n747), .A1(A[14]) );
  inv01 U640 ( .Y(n584), .A(n595) );
  nor02 U641 ( .Y(n596), .A0(n576), .A1(n577) );
  inv01 U642 ( .Y(n586), .A(n596) );
  nor02 U643 ( .Y(n597), .A0(n579), .A1(n581) );
  inv01 U644 ( .Y(n587), .A(n597) );
  nor02 U645 ( .Y(n598), .A0(n583), .A1(n585) );
  inv01 U646 ( .Y(n588), .A(n598) );
  nor02 U647 ( .Y(n599), .A0(n589), .A1(n590) );
  inv01 U648 ( .Y(n592), .A(n599) );
  inv02 U649 ( .Y(SUM[15]), .A(n600) );
  inv02 U650 ( .Y(carry_16_), .A(n601) );
  inv02 U651 ( .Y(n602), .A(n709) );
  inv02 U652 ( .Y(n603), .A(A[15]) );
  inv02 U653 ( .Y(n604), .A(carry_15_) );
  nor02 U654 ( .Y(n605), .A0(n602), .A1(n606) );
  nor02 U655 ( .Y(n607), .A0(n603), .A1(n608) );
  nor02 U656 ( .Y(n609), .A0(n604), .A1(n610) );
  nor02 U657 ( .Y(n611), .A0(n604), .A1(n612) );
  nor02 U658 ( .Y(n600), .A0(n613), .A1(n614) );
  nor02 U659 ( .Y(n615), .A0(n603), .A1(n604) );
  nor02 U660 ( .Y(n616), .A0(n602), .A1(n604) );
  nor02 U661 ( .Y(n617), .A0(n602), .A1(n603) );
  nor02 U662 ( .Y(n601), .A0(n617), .A1(n618) );
  nor02 U663 ( .Y(n619), .A0(A[15]), .A1(carry_15_) );
  inv01 U664 ( .Y(n606), .A(n619) );
  nor02 U665 ( .Y(n620), .A0(n709), .A1(carry_15_) );
  inv01 U666 ( .Y(n608), .A(n620) );
  nor02 U667 ( .Y(n621), .A0(n709), .A1(A[15]) );
  inv01 U668 ( .Y(n610), .A(n621) );
  nor02 U669 ( .Y(n622), .A0(n602), .A1(n603) );
  inv01 U670 ( .Y(n612), .A(n622) );
  nor02 U671 ( .Y(n623), .A0(n605), .A1(n607) );
  inv01 U672 ( .Y(n613), .A(n623) );
  nor02 U673 ( .Y(n624), .A0(n609), .A1(n611) );
  inv02 U674 ( .Y(n614), .A(n624) );
  nor02 U675 ( .Y(n625), .A0(n615), .A1(n616) );
  inv01 U676 ( .Y(n618), .A(n625) );
  inv02 U677 ( .Y(SUM[22]), .A(n626) );
  inv02 U678 ( .Y(carry_23_), .A(n627) );
  inv02 U679 ( .Y(n628), .A(n743) );
  inv02 U680 ( .Y(n629), .A(A[22]) );
  inv02 U681 ( .Y(n630), .A(carry_22_) );
  nor02 U682 ( .Y(n631), .A0(n628), .A1(n632) );
  nor02 U683 ( .Y(n633), .A0(n629), .A1(n634) );
  nor02 U684 ( .Y(n635), .A0(n630), .A1(n636) );
  nor02 U685 ( .Y(n637), .A0(n630), .A1(n638) );
  nor02 U686 ( .Y(n626), .A0(n639), .A1(n640) );
  nor02 U687 ( .Y(n641), .A0(n629), .A1(n630) );
  nor02 U688 ( .Y(n642), .A0(n628), .A1(n630) );
  nor02 U689 ( .Y(n643), .A0(n628), .A1(n629) );
  nor02 U690 ( .Y(n627), .A0(n643), .A1(n644) );
  nor02 U691 ( .Y(n645), .A0(A[22]), .A1(carry_22_) );
  inv01 U692 ( .Y(n632), .A(n645) );
  nor02 U693 ( .Y(n646), .A0(n743), .A1(carry_22_) );
  inv01 U694 ( .Y(n634), .A(n646) );
  nor02 U695 ( .Y(n647), .A0(n743), .A1(A[22]) );
  inv01 U696 ( .Y(n636), .A(n647) );
  nor02 U697 ( .Y(n648), .A0(n628), .A1(n629) );
  inv01 U698 ( .Y(n638), .A(n648) );
  nor02 U699 ( .Y(n649), .A0(n631), .A1(n633) );
  inv01 U700 ( .Y(n639), .A(n649) );
  nor02 U701 ( .Y(n650), .A0(n635), .A1(n637) );
  inv01 U702 ( .Y(n640), .A(n650) );
  nor02 U703 ( .Y(n651), .A0(n641), .A1(n642) );
  inv01 U704 ( .Y(n644), .A(n651) );
  inv02 U705 ( .Y(SUM[0]), .A(n652) );
  inv02 U706 ( .Y(carry_1_), .A(n653) );
  inv02 U707 ( .Y(n654), .A(n711) );
  inv02 U708 ( .Y(n655), .A(A[0]) );
  inv02 U709 ( .Y(n656), .A(ADD_SUB) );
  nor02 U710 ( .Y(n657), .A0(n654), .A1(n658) );
  nor02 U711 ( .Y(n659), .A0(n655), .A1(n660) );
  nor02 U712 ( .Y(n661), .A0(n656), .A1(n662) );
  nor02 U713 ( .Y(n663), .A0(n656), .A1(n664) );
  nor02 U714 ( .Y(n652), .A0(n665), .A1(n666) );
  nor02 U715 ( .Y(n667), .A0(n655), .A1(n656) );
  nor02 U716 ( .Y(n668), .A0(n654), .A1(n656) );
  nor02 U717 ( .Y(n669), .A0(n654), .A1(n655) );
  nor02 U718 ( .Y(n653), .A0(n669), .A1(n670) );
  nor02 U719 ( .Y(n671), .A0(A[0]), .A1(ADD_SUB) );
  inv01 U720 ( .Y(n658), .A(n671) );
  nor02 U721 ( .Y(n672), .A0(n711), .A1(ADD_SUB) );
  inv01 U722 ( .Y(n660), .A(n672) );
  nor02 U723 ( .Y(n673), .A0(n711), .A1(A[0]) );
  inv01 U724 ( .Y(n662), .A(n673) );
  nor02 U725 ( .Y(n674), .A0(n654), .A1(n655) );
  inv01 U726 ( .Y(n664), .A(n674) );
  nor02 U727 ( .Y(n675), .A0(n657), .A1(n659) );
  inv01 U728 ( .Y(n665), .A(n675) );
  nor02 U729 ( .Y(n676), .A0(n661), .A1(n663) );
  inv01 U730 ( .Y(n666), .A(n676) );
  nor02 U731 ( .Y(n677), .A0(n667), .A1(n668) );
  inv01 U732 ( .Y(n670), .A(n677) );
  inv02 U733 ( .Y(SUM[16]), .A(n678) );
  inv02 U734 ( .Y(carry_17_), .A(n679) );
  inv02 U735 ( .Y(n680), .A(n751) );
  inv02 U736 ( .Y(n681), .A(A[16]) );
  inv02 U737 ( .Y(n682), .A(carry_16_) );
  nor02 U738 ( .Y(n683), .A0(n680), .A1(n684) );
  nor02 U739 ( .Y(n685), .A0(n681), .A1(n686) );
  nor02 U740 ( .Y(n687), .A0(n682), .A1(n688) );
  nor02 U741 ( .Y(n689), .A0(n682), .A1(n690) );
  nor02 U742 ( .Y(n678), .A0(n691), .A1(n692) );
  nor02 U743 ( .Y(n693), .A0(n681), .A1(n682) );
  nor02 U744 ( .Y(n694), .A0(n680), .A1(n682) );
  nor02 U745 ( .Y(n695), .A0(n680), .A1(n681) );
  nor02 U746 ( .Y(n679), .A0(n695), .A1(n696) );
  nor02 U747 ( .Y(n697), .A0(A[16]), .A1(carry_16_) );
  inv01 U748 ( .Y(n684), .A(n697) );
  nor02 U749 ( .Y(n698), .A0(n751), .A1(carry_16_) );
  inv01 U750 ( .Y(n686), .A(n698) );
  nor02 U751 ( .Y(n699), .A0(n751), .A1(A[16]) );
  inv01 U752 ( .Y(n688), .A(n699) );
  nor02 U753 ( .Y(n700), .A0(n680), .A1(n681) );
  inv01 U754 ( .Y(n690), .A(n700) );
  nor02 U755 ( .Y(n701), .A0(n683), .A1(n685) );
  inv01 U756 ( .Y(n691), .A(n701) );
  nor02 U757 ( .Y(n702), .A0(n687), .A1(n689) );
  inv01 U758 ( .Y(n692), .A(n702) );
  nor02 U759 ( .Y(n703), .A0(n693), .A1(n694) );
  inv01 U760 ( .Y(n696), .A(n703) );
  xor2 U761 ( .Y(n704), .A0(B[1]), .A1(n760) );
  inv02 U762 ( .Y(n705), .A(n704) );
  xor2 U763 ( .Y(n706), .A0(B[13]), .A1(n760) );
  inv02 U764 ( .Y(n707), .A(n706) );
  xor2 U765 ( .Y(n708), .A0(B[15]), .A1(n760) );
  inv02 U766 ( .Y(n709), .A(n708) );
  xor2 U767 ( .Y(n710), .A0(B[0]), .A1(n761) );
  inv02 U768 ( .Y(n711), .A(n710) );
  xor2 U769 ( .Y(n712), .A0(B[26]), .A1(n761) );
  inv02 U770 ( .Y(n713), .A(n712) );
  xor2 U771 ( .Y(n714), .A0(B[19]), .A1(n760) );
  inv02 U772 ( .Y(n715), .A(n714) );
  xor2 U773 ( .Y(n716), .A0(B[7]), .A1(n761) );
  inv02 U774 ( .Y(n717), .A(n716) );
  xor2 U775 ( .Y(n718), .A0(B[5]), .A1(n761) );
  inv02 U776 ( .Y(n719), .A(n718) );
  xor2 U777 ( .Y(n720), .A0(B[25]), .A1(n761) );
  inv02 U778 ( .Y(n721), .A(n720) );
  xor2 U779 ( .Y(n722), .A0(B[17]), .A1(n760) );
  inv02 U780 ( .Y(n723), .A(n722) );
  xor2 U781 ( .Y(n724), .A0(B[21]), .A1(n760) );
  inv02 U782 ( .Y(n725), .A(n724) );
  xor2 U783 ( .Y(n726), .A0(B[11]), .A1(n760) );
  inv02 U784 ( .Y(n727), .A(n726) );
  xor2 U785 ( .Y(n728), .A0(B[23]), .A1(n760) );
  inv02 U786 ( .Y(n729), .A(n728) );
  xor2 U787 ( .Y(n730), .A0(B[12]), .A1(n760) );
  inv02 U788 ( .Y(n731), .A(n730) );
  xor2 U789 ( .Y(n732), .A0(B[9]), .A1(n760) );
  inv02 U790 ( .Y(n733), .A(n732) );
  xor2 U791 ( .Y(n734), .A0(B[10]), .A1(n761) );
  inv02 U792 ( .Y(n735), .A(n734) );
  xor2 U793 ( .Y(n736), .A0(B[3]), .A1(n761) );
  inv02 U794 ( .Y(n737), .A(n736) );
  xor2 U795 ( .Y(n738), .A0(B[4]), .A1(n761) );
  inv02 U796 ( .Y(n739), .A(n738) );
  xor2 U797 ( .Y(n740), .A0(B[8]), .A1(n761) );
  inv02 U798 ( .Y(n741), .A(n740) );
  xor2 U799 ( .Y(n742), .A0(B[22]), .A1(n760) );
  inv02 U800 ( .Y(n743), .A(n742) );
  xor2 U801 ( .Y(n744), .A0(B[6]), .A1(n761) );
  inv02 U802 ( .Y(n745), .A(n744) );
  xor2 U803 ( .Y(n746), .A0(B[14]), .A1(n761) );
  inv02 U804 ( .Y(n747), .A(n746) );
  xor2 U805 ( .Y(n748), .A0(B[18]), .A1(n760) );
  inv02 U806 ( .Y(n749), .A(n748) );
  xor2 U807 ( .Y(n750), .A0(B[16]), .A1(n760) );
  inv02 U808 ( .Y(n751), .A(n750) );
  xor2 U809 ( .Y(n752), .A0(B[20]), .A1(n760) );
  inv02 U810 ( .Y(n753), .A(n752) );
  xor2 U811 ( .Y(n754), .A0(B[27]), .A1(n761) );
  inv02 U812 ( .Y(n755), .A(n754) );
  xor2 U813 ( .Y(n756), .A0(B[2]), .A1(n761) );
  inv02 U814 ( .Y(n757), .A(n756) );
  xor2 U815 ( .Y(n758), .A0(B[24]), .A1(n761) );
  inv02 U816 ( .Y(n759), .A(n758) );
  buf12 U817 ( .Y(n760), .A(n762) );
  buf12 U818 ( .Y(n761), .A(n762) );
  inv01 U819 ( .Y(n762), .A(ADD_SUB) );
  fadd1 U1_27 ( .S(n763), .A(A[27]), .B(n755), .CI(carry_27_) );
endmodule


module addsub_28_DW01_cmp2_28_0 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [27:0] A;
  input [27:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165;

  buf02 U6 ( .Y(n15), .A(n97) );
  nand02 U7 ( .Y(LT_LE), .A0(n16), .A1(n17) );
  nand02 U8 ( .Y(n16), .A0(B[27]), .A1(n96) );
  inv01 U9 ( .Y(n17), .A(n15) );
  inv01 U10 ( .Y(n99), .A(n18) );
  nor02 U11 ( .Y(n19), .A0(B[26]), .A1(n101) );
  nor02 U12 ( .Y(n20), .A0(B[25]), .A1(n102) );
  inv01 U13 ( .Y(n21), .A(n103) );
  nor02 U14 ( .Y(n18), .A0(n21), .A1(n22) );
  nor02 U15 ( .Y(n23), .A0(n19), .A1(n20) );
  inv01 U16 ( .Y(n22), .A(n23) );
  inv02 U17 ( .Y(n102), .A(A[25]) );
  inv02 U18 ( .Y(n101), .A(A[26]) );
  inv01 U19 ( .Y(n161), .A(n24) );
  nor02 U20 ( .Y(n25), .A0(B[2]), .A1(n159) );
  nor02 U21 ( .Y(n26), .A0(n162), .A1(n163) );
  inv01 U22 ( .Y(n27), .A(n164) );
  nor02 U23 ( .Y(n24), .A0(n27), .A1(n28) );
  nor02 U24 ( .Y(n29), .A0(n25), .A1(n26) );
  inv01 U25 ( .Y(n28), .A(n29) );
  inv01 U26 ( .Y(n160), .A(n161) );
  inv02 U27 ( .Y(n163), .A(A[1]) );
  inv02 U28 ( .Y(n159), .A(A[2]) );
  inv01 U29 ( .Y(n141), .A(n30) );
  nor02 U30 ( .Y(n31), .A0(B[9]), .A1(n142) );
  nor02 U31 ( .Y(n32), .A0(B[10]), .A1(n139) );
  inv01 U32 ( .Y(n33), .A(n143) );
  nor02 U33 ( .Y(n30), .A0(n33), .A1(n34) );
  nor02 U34 ( .Y(n35), .A0(n31), .A1(n32) );
  inv01 U35 ( .Y(n34), .A(n35) );
  inv01 U36 ( .Y(n121), .A(n36) );
  nor02 U37 ( .Y(n37), .A0(B[18]), .A1(n119) );
  nor02 U38 ( .Y(n38), .A0(B[17]), .A1(n122) );
  inv01 U39 ( .Y(n39), .A(n123) );
  nor02 U40 ( .Y(n36), .A0(n39), .A1(n40) );
  nor02 U41 ( .Y(n41), .A0(n37), .A1(n38) );
  inv01 U42 ( .Y(n40), .A(n41) );
  inv01 U43 ( .Y(n140), .A(n141) );
  inv02 U44 ( .Y(n139), .A(A[10]) );
  inv02 U45 ( .Y(n142), .A(A[9]) );
  inv01 U46 ( .Y(n120), .A(n121) );
  inv02 U47 ( .Y(n122), .A(A[17]) );
  inv02 U48 ( .Y(n119), .A(A[18]) );
  inv01 U49 ( .Y(n136), .A(n42) );
  nor02 U50 ( .Y(n43), .A0(B[12]), .A1(n134) );
  nor02 U51 ( .Y(n44), .A0(B[11]), .A1(n137) );
  inv01 U52 ( .Y(n45), .A(n138) );
  nor02 U53 ( .Y(n42), .A0(n45), .A1(n46) );
  nor02 U54 ( .Y(n47), .A0(n43), .A1(n44) );
  inv01 U55 ( .Y(n46), .A(n47) );
  inv01 U56 ( .Y(n135), .A(n136) );
  inv02 U57 ( .Y(n137), .A(A[11]) );
  inv02 U58 ( .Y(n134), .A(A[12]) );
  inv01 U59 ( .Y(n116), .A(n48) );
  nor02 U60 ( .Y(n49), .A0(B[20]), .A1(n114) );
  nor02 U61 ( .Y(n50), .A0(B[19]), .A1(n117) );
  inv01 U62 ( .Y(n51), .A(n118) );
  nor02 U63 ( .Y(n48), .A0(n51), .A1(n52) );
  nor02 U64 ( .Y(n53), .A0(n49), .A1(n50) );
  inv01 U65 ( .Y(n52), .A(n53) );
  inv01 U66 ( .Y(n131), .A(n54) );
  nor02 U67 ( .Y(n55), .A0(B[14]), .A1(n129) );
  nor02 U68 ( .Y(n56), .A0(B[13]), .A1(n132) );
  inv01 U69 ( .Y(n57), .A(n133) );
  nor02 U70 ( .Y(n54), .A0(n57), .A1(n58) );
  nor02 U71 ( .Y(n59), .A0(n55), .A1(n56) );
  inv01 U72 ( .Y(n58), .A(n59) );
  inv01 U73 ( .Y(n115), .A(n116) );
  inv02 U74 ( .Y(n117), .A(A[19]) );
  inv02 U75 ( .Y(n114), .A(A[20]) );
  inv01 U76 ( .Y(n130), .A(n131) );
  inv02 U77 ( .Y(n132), .A(A[13]) );
  inv02 U78 ( .Y(n129), .A(A[14]) );
  inv01 U79 ( .Y(n111), .A(n60) );
  nor02 U80 ( .Y(n61), .A0(B[22]), .A1(n109) );
  nor02 U81 ( .Y(n62), .A0(B[21]), .A1(n112) );
  inv01 U82 ( .Y(n63), .A(n113) );
  nor02 U83 ( .Y(n60), .A0(n63), .A1(n64) );
  nor02 U84 ( .Y(n65), .A0(n61), .A1(n62) );
  inv01 U85 ( .Y(n64), .A(n65) );
  inv01 U86 ( .Y(n156), .A(n66) );
  nor02 U87 ( .Y(n67), .A0(B[4]), .A1(n154) );
  nor02 U88 ( .Y(n68), .A0(B[3]), .A1(n157) );
  inv01 U89 ( .Y(n69), .A(n158) );
  nor02 U90 ( .Y(n66), .A0(n69), .A1(n70) );
  nor02 U91 ( .Y(n71), .A0(n67), .A1(n68) );
  inv01 U92 ( .Y(n70), .A(n71) );
  inv01 U93 ( .Y(n110), .A(n111) );
  inv02 U94 ( .Y(n112), .A(A[21]) );
  inv02 U95 ( .Y(n109), .A(A[22]) );
  inv01 U96 ( .Y(n155), .A(n156) );
  inv02 U97 ( .Y(n157), .A(A[3]) );
  inv02 U98 ( .Y(n154), .A(A[4]) );
  inv01 U99 ( .Y(n126), .A(n72) );
  nor02 U100 ( .Y(n73), .A0(B[16]), .A1(n124) );
  nor02 U101 ( .Y(n74), .A0(B[15]), .A1(n127) );
  inv01 U102 ( .Y(n75), .A(n128) );
  nor02 U103 ( .Y(n72), .A0(n75), .A1(n76) );
  nor02 U104 ( .Y(n77), .A0(n73), .A1(n74) );
  inv01 U105 ( .Y(n76), .A(n77) );
  inv01 U106 ( .Y(n151), .A(n78) );
  nor02 U107 ( .Y(n79), .A0(B[6]), .A1(n149) );
  nor02 U108 ( .Y(n80), .A0(B[5]), .A1(n152) );
  inv01 U109 ( .Y(n81), .A(n153) );
  nor02 U110 ( .Y(n78), .A0(n81), .A1(n82) );
  nor02 U111 ( .Y(n83), .A0(n79), .A1(n80) );
  inv01 U112 ( .Y(n82), .A(n83) );
  inv01 U113 ( .Y(n125), .A(n126) );
  inv02 U114 ( .Y(n127), .A(A[15]) );
  inv02 U115 ( .Y(n124), .A(A[16]) );
  inv01 U116 ( .Y(n150), .A(n151) );
  inv02 U117 ( .Y(n152), .A(A[5]) );
  inv02 U118 ( .Y(n149), .A(A[6]) );
  inv01 U119 ( .Y(n106), .A(n84) );
  nor02 U120 ( .Y(n85), .A0(B[24]), .A1(n104) );
  nor02 U121 ( .Y(n86), .A0(B[23]), .A1(n107) );
  inv01 U122 ( .Y(n87), .A(n108) );
  nor02 U123 ( .Y(n84), .A0(n87), .A1(n88) );
  nor02 U124 ( .Y(n89), .A0(n85), .A1(n86) );
  inv01 U125 ( .Y(n88), .A(n89) );
  inv01 U126 ( .Y(n146), .A(n90) );
  nor02 U127 ( .Y(n91), .A0(B[8]), .A1(n144) );
  nor02 U128 ( .Y(n92), .A0(B[7]), .A1(n147) );
  inv01 U129 ( .Y(n93), .A(n148) );
  nor02 U130 ( .Y(n90), .A0(n93), .A1(n94) );
  nor02 U131 ( .Y(n95), .A0(n91), .A1(n92) );
  inv01 U132 ( .Y(n94), .A(n95) );
  inv01 U133 ( .Y(n105), .A(n106) );
  inv02 U134 ( .Y(n107), .A(A[23]) );
  inv02 U135 ( .Y(n104), .A(A[24]) );
  inv01 U136 ( .Y(n145), .A(n146) );
  inv02 U137 ( .Y(n147), .A(A[7]) );
  inv02 U138 ( .Y(n144), .A(A[8]) );
  inv04 U139 ( .Y(n165), .A(B[0]) );
  inv04 U140 ( .Y(n98), .A(B[27]) );
  inv04 U141 ( .Y(n96), .A(A[27]) );
  aoi22 U142 ( .Y(n97), .A0(A[27]), .A1(n98), .B0(n99), .B1(n100) );
  nand02 U143 ( .Y(n100), .A0(B[26]), .A1(n101) );
  ao221 U144 ( .Y(n103), .A0(n104), .A1(B[24]), .B0(n102), .B1(B[25]), .C0(
        n105) );
  ao221 U145 ( .Y(n108), .A0(n109), .A1(B[22]), .B0(n107), .B1(B[23]), .C0(
        n110) );
  ao221 U146 ( .Y(n113), .A0(n114), .A1(B[20]), .B0(n112), .B1(B[21]), .C0(
        n115) );
  ao221 U147 ( .Y(n118), .A0(n119), .A1(B[18]), .B0(n117), .B1(B[19]), .C0(
        n120) );
  ao221 U148 ( .Y(n123), .A0(n124), .A1(B[16]), .B0(n122), .B1(B[17]), .C0(
        n125) );
  ao221 U149 ( .Y(n128), .A0(n129), .A1(B[14]), .B0(n127), .B1(B[15]), .C0(
        n130) );
  ao221 U150 ( .Y(n133), .A0(n134), .A1(B[12]), .B0(n132), .B1(B[13]), .C0(
        n135) );
  ao221 U151 ( .Y(n138), .A0(n139), .A1(B[10]), .B0(n137), .B1(B[11]), .C0(
        n140) );
  ao221 U152 ( .Y(n143), .A0(n144), .A1(B[8]), .B0(n142), .B1(B[9]), .C0(n145)
         );
  ao221 U153 ( .Y(n148), .A0(n149), .A1(B[6]), .B0(n147), .B1(B[7]), .C0(n150)
         );
  ao221 U154 ( .Y(n153), .A0(n154), .A1(B[4]), .B0(n152), .B1(B[5]), .C0(n155)
         );
  ao221 U155 ( .Y(n158), .A0(n159), .A1(B[2]), .B0(n157), .B1(B[3]), .C0(n160)
         );
  ao21 U156 ( .Y(n164), .A0(n162), .A1(n163), .B0(B[1]) );
  nor02 U157 ( .Y(n162), .A0(n165), .A1(A[0]) );
endmodule


module addsub_28 ( clk_i, fpu_op_i, fracta_i, fractb_i, signa_i, signb_i, 
        fract_o, sign_o );
  input [27:0] fracta_i;
  input [27:0] fractb_i;
  output [27:0] fract_o;
  input clk_i, fpu_op_i, signa_i, signb_i;
  output sign_o;
  wire   s_sign_o, n____return53, U42_U3_Z_0, U42_U2_Z_27, U42_U2_Z_26,
         U42_U2_Z_25, U42_U2_Z_24, U42_U2_Z_23, U42_U2_Z_22, U42_U2_Z_21,
         U42_U2_Z_20, U42_U2_Z_19, U42_U2_Z_18, U42_U2_Z_17, U42_U2_Z_16,
         U42_U2_Z_15, U42_U2_Z_14, U42_U2_Z_13, U42_U2_Z_12, U42_U2_Z_11,
         U42_U2_Z_10, U42_U2_Z_9, U42_U2_Z_8, U42_U2_Z_7, U42_U2_Z_6,
         U42_U2_Z_5, U42_U2_Z_4, U42_U2_Z_3, U42_U2_Z_2, U42_U2_Z_1,
         U42_U2_Z_0, U42_U1_Z_27, U42_U1_Z_26, U42_U1_Z_25, U42_U1_Z_24,
         U42_U1_Z_23, U42_U1_Z_22, U42_U1_Z_21, U42_U1_Z_20, U42_U1_Z_19,
         U42_U1_Z_18, U42_U1_Z_17, U42_U1_Z_16, U42_U1_Z_15, U42_U1_Z_14,
         U42_U1_Z_13, U42_U1_Z_12, U42_U1_Z_11, U42_U1_Z_10, U42_U1_Z_9,
         U42_U1_Z_8, U42_U1_Z_7, U42_U1_Z_6, U42_U1_Z_5, U42_U1_Z_4,
         U42_U1_Z_3, U42_U1_Z_2, U42_U1_Z_1, U42_U1_Z_0, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611;
  wire   [27:0] s_fract_o;

  dff fract_o_reg_27_ ( .QB(n540), .D(s_fract_o[27]), .CLK(clk_i) );
  dff fract_o_reg_26_ ( .Q(fract_o[26]), .D(s_fract_o[26]), .CLK(clk_i) );
  dff fract_o_reg_25_ ( .Q(fract_o[25]), .D(s_fract_o[25]), .CLK(clk_i) );
  dff fract_o_reg_24_ ( .Q(fract_o[24]), .D(s_fract_o[24]), .CLK(clk_i) );
  dff fract_o_reg_23_ ( .Q(fract_o[23]), .D(s_fract_o[23]), .CLK(clk_i) );
  dff fract_o_reg_22_ ( .Q(fract_o[22]), .D(s_fract_o[22]), .CLK(clk_i) );
  dff fract_o_reg_21_ ( .Q(fract_o[21]), .D(s_fract_o[21]), .CLK(clk_i) );
  dff fract_o_reg_20_ ( .Q(fract_o[20]), .D(s_fract_o[20]), .CLK(clk_i) );
  dff fract_o_reg_19_ ( .Q(fract_o[19]), .D(s_fract_o[19]), .CLK(clk_i) );
  dff fract_o_reg_18_ ( .Q(fract_o[18]), .D(s_fract_o[18]), .CLK(clk_i) );
  dff fract_o_reg_17_ ( .Q(fract_o[17]), .D(s_fract_o[17]), .CLK(clk_i) );
  dff fract_o_reg_16_ ( .Q(fract_o[16]), .D(s_fract_o[16]), .CLK(clk_i) );
  dff fract_o_reg_15_ ( .Q(fract_o[15]), .D(s_fract_o[15]), .CLK(clk_i) );
  dff fract_o_reg_14_ ( .Q(fract_o[14]), .D(s_fract_o[14]), .CLK(clk_i) );
  dff fract_o_reg_13_ ( .Q(fract_o[13]), .D(s_fract_o[13]), .CLK(clk_i) );
  dff fract_o_reg_12_ ( .Q(fract_o[12]), .D(s_fract_o[12]), .CLK(clk_i) );
  dff fract_o_reg_11_ ( .Q(fract_o[11]), .D(s_fract_o[11]), .CLK(clk_i) );
  dff fract_o_reg_10_ ( .Q(fract_o[10]), .D(s_fract_o[10]), .CLK(clk_i) );
  dff fract_o_reg_9_ ( .Q(fract_o[9]), .D(s_fract_o[9]), .CLK(clk_i) );
  dff fract_o_reg_8_ ( .Q(fract_o[8]), .D(s_fract_o[8]), .CLK(clk_i) );
  dff fract_o_reg_7_ ( .Q(fract_o[7]), .D(s_fract_o[7]), .CLK(clk_i) );
  dff fract_o_reg_6_ ( .Q(fract_o[6]), .D(s_fract_o[6]), .CLK(clk_i) );
  dff fract_o_reg_5_ ( .Q(fract_o[5]), .D(s_fract_o[5]), .CLK(clk_i) );
  dff fract_o_reg_4_ ( .Q(fract_o[4]), .D(s_fract_o[4]), .CLK(clk_i) );
  dff fract_o_reg_3_ ( .Q(fract_o[3]), .D(s_fract_o[3]), .CLK(clk_i) );
  dff fract_o_reg_2_ ( .Q(fract_o[2]), .D(s_fract_o[2]), .CLK(clk_i) );
  dff fract_o_reg_1_ ( .Q(fract_o[1]), .D(s_fract_o[1]), .CLK(clk_i) );
  dff fract_o_reg_0_ ( .Q(fract_o[0]), .D(s_fract_o[0]), .CLK(clk_i) );
  dff sign_o_reg ( .Q(sign_o), .D(s_sign_o), .CLK(clk_i) );
  nand02 U182 ( .Y(n547), .A0(n419), .A1(n420) );
  inv01 U183 ( .Y(n421), .A(signa_i) );
  inv01 U184 ( .Y(n422), .A(n463) );
  inv01 U185 ( .Y(n423), .A(n____return53) );
  nand02 U186 ( .Y(n419), .A0(n____return53), .A1(n421) );
  nand02 U187 ( .Y(n420), .A0(n422), .A1(n423) );
  buf02 U188 ( .Y(n424), .A(U42_U2_Z_19) );
  buf02 U189 ( .Y(n425), .A(U42_U2_Z_15) );
  buf02 U190 ( .Y(n426), .A(U42_U2_Z_26) );
  buf02 U191 ( .Y(n427), .A(U42_U2_Z_1) );
  buf02 U192 ( .Y(n428), .A(U42_U2_Z_9) );
  buf02 U193 ( .Y(n429), .A(U42_U2_Z_11) );
  buf02 U194 ( .Y(n430), .A(U42_U2_Z_21) );
  buf02 U195 ( .Y(n431), .A(U42_U2_Z_25) );
  buf02 U196 ( .Y(n432), .A(U42_U2_Z_3) );
  buf02 U197 ( .Y(n433), .A(U42_U2_Z_5) );
  buf02 U198 ( .Y(n434), .A(U42_U2_Z_23) );
  buf02 U199 ( .Y(n435), .A(U42_U2_Z_7) );
  buf02 U200 ( .Y(n436), .A(U42_U2_Z_16) );
  buf02 U201 ( .Y(n437), .A(U42_U2_Z_24) );
  buf02 U202 ( .Y(n438), .A(U42_U2_Z_17) );
  buf02 U203 ( .Y(n439), .A(U42_U2_Z_13) );
  buf02 U204 ( .Y(n440), .A(U42_U2_Z_22) );
  buf02 U205 ( .Y(n441), .A(U42_U2_Z_8) );
  buf02 U206 ( .Y(n442), .A(U42_U2_Z_2) );
  buf02 U207 ( .Y(n443), .A(U42_U2_Z_14) );
  buf02 U208 ( .Y(n444), .A(U42_U2_Z_4) );
  buf02 U209 ( .Y(n445), .A(U42_U2_Z_18) );
  buf02 U210 ( .Y(n446), .A(U42_U2_Z_20) );
  buf02 U211 ( .Y(n447), .A(U42_U2_Z_10) );
  buf02 U212 ( .Y(n448), .A(U42_U2_Z_12) );
  buf02 U213 ( .Y(n449), .A(U42_U2_Z_6) );
  buf02 U214 ( .Y(n450), .A(U42_U2_Z_0) );
  buf02 U215 ( .Y(n451), .A(U42_U2_Z_27) );
  nand02 U216 ( .Y(s_sign_o), .A0(n452), .A1(n453) );
  inv01 U217 ( .Y(n454), .A(n547) );
  inv01 U218 ( .Y(n455), .A(n546) );
  inv01 U219 ( .Y(n456), .A(n545) );
  nand02 U220 ( .Y(n452), .A0(n454), .A1(n455) );
  nand02 U221 ( .Y(n453), .A0(n454), .A1(n456) );
  or03 U222 ( .Y(n457), .A0(s_fract_o[21]), .A1(s_fract_o[23]), .A2(
        s_fract_o[22]) );
  inv01 U223 ( .Y(n458), .A(n457) );
  or03 U224 ( .Y(n459), .A0(n554), .A1(s_fract_o[10]), .A2(s_fract_o[0]) );
  inv01 U225 ( .Y(n460), .A(n459) );
  or03 U226 ( .Y(n461), .A0(s_fract_o[15]), .A1(s_fract_o[17]), .A2(
        s_fract_o[16]) );
  inv01 U227 ( .Y(n462), .A(n461) );
  buf02 U228 ( .Y(n463), .A(n548) );
  xor2 U229 ( .Y(n464), .A0(n463), .A1(signa_i) );
  inv01 U230 ( .Y(n465), .A(n464) );
  inv04 U231 ( .Y(fract_o[27]), .A(n540) );
  buf08 U232 ( .Y(n466), .A(n542) );
  inv02 U233 ( .Y(n542), .A(n557) );
  inv01 U234 ( .Y(n549), .A(n467) );
  inv01 U235 ( .Y(n468), .A(s_fract_o[24]) );
  inv01 U236 ( .Y(n469), .A(s_fract_o[25]) );
  inv01 U237 ( .Y(n470), .A(s_fract_o[26]) );
  inv01 U238 ( .Y(n471), .A(s_fract_o[27]) );
  nand02 U239 ( .Y(n467), .A0(n472), .A1(n473) );
  nand02 U240 ( .Y(n474), .A0(n468), .A1(n469) );
  inv01 U241 ( .Y(n472), .A(n474) );
  nand02 U242 ( .Y(n475), .A0(n470), .A1(n471) );
  inv01 U243 ( .Y(n473), .A(n475) );
  inv01 U244 ( .Y(n552), .A(n476) );
  inv01 U245 ( .Y(n477), .A(s_fract_o[11]) );
  inv01 U246 ( .Y(n478), .A(s_fract_o[12]) );
  inv01 U247 ( .Y(n479), .A(s_fract_o[13]) );
  inv01 U248 ( .Y(n480), .A(s_fract_o[14]) );
  nand02 U249 ( .Y(n476), .A0(n481), .A1(n482) );
  nand02 U250 ( .Y(n483), .A0(n477), .A1(n478) );
  inv01 U251 ( .Y(n481), .A(n483) );
  nand02 U252 ( .Y(n484), .A0(n479), .A1(n480) );
  inv01 U253 ( .Y(n482), .A(n484) );
  inv01 U254 ( .Y(n550), .A(n485) );
  inv01 U255 ( .Y(n486), .A(s_fract_o[2]) );
  inv01 U256 ( .Y(n487), .A(s_fract_o[3]) );
  inv01 U257 ( .Y(n488), .A(s_fract_o[4]) );
  inv01 U258 ( .Y(n489), .A(s_fract_o[5]) );
  nand02 U259 ( .Y(n485), .A0(n490), .A1(n491) );
  nand02 U260 ( .Y(n492), .A0(n486), .A1(n487) );
  inv01 U261 ( .Y(n490), .A(n492) );
  nand02 U262 ( .Y(n493), .A0(n488), .A1(n489) );
  inv01 U263 ( .Y(n491), .A(n493) );
  buf02 U264 ( .Y(n494), .A(U42_U1_Z_6) );
  buf02 U265 ( .Y(n495), .A(U42_U1_Z_12) );
  buf02 U266 ( .Y(n496), .A(U42_U1_Z_20) );
  buf02 U267 ( .Y(n497), .A(U42_U1_Z_0) );
  buf02 U268 ( .Y(n498), .A(U42_U1_Z_13) );
  buf02 U269 ( .Y(n499), .A(U42_U1_Z_17) );
  buf02 U270 ( .Y(n500), .A(U42_U1_Z_14) );
  buf02 U271 ( .Y(n501), .A(U42_U1_Z_11) );
  buf02 U272 ( .Y(n502), .A(U42_U1_Z_5) );
  buf02 U273 ( .Y(n503), .A(U42_U1_Z_3) );
  buf02 U274 ( .Y(n504), .A(U42_U1_Z_26) );
  buf02 U275 ( .Y(n505), .A(U42_U1_Z_24) );
  buf02 U276 ( .Y(n506), .A(U42_U1_Z_4) );
  buf02 U277 ( .Y(n507), .A(U42_U1_Z_22) );
  buf02 U278 ( .Y(n508), .A(U42_U1_Z_16) );
  buf02 U279 ( .Y(n509), .A(U42_U1_Z_23) );
  buf02 U280 ( .Y(n510), .A(U42_U1_Z_8) );
  buf02 U281 ( .Y(n511), .A(U42_U1_Z_15) );
  buf02 U282 ( .Y(n512), .A(U42_U1_Z_9) );
  buf02 U283 ( .Y(n513), .A(U42_U1_Z_10) );
  buf02 U284 ( .Y(n514), .A(U42_U1_Z_2) );
  buf02 U285 ( .Y(n515), .A(U42_U1_Z_19) );
  buf02 U286 ( .Y(n516), .A(U42_U1_Z_21) );
  buf02 U287 ( .Y(n517), .A(U42_U1_Z_7) );
  buf02 U288 ( .Y(n518), .A(U42_U1_Z_1) );
  buf02 U289 ( .Y(n519), .A(U42_U1_Z_25) );
  buf02 U290 ( .Y(n520), .A(U42_U1_Z_18) );
  buf02 U291 ( .Y(n521), .A(U42_U1_Z_27) );
  inv01 U292 ( .Y(n551), .A(n522) );
  inv01 U293 ( .Y(n523), .A(s_fract_o[6]) );
  inv01 U294 ( .Y(n524), .A(s_fract_o[7]) );
  inv01 U295 ( .Y(n525), .A(s_fract_o[8]) );
  inv01 U296 ( .Y(n526), .A(s_fract_o[9]) );
  nand02 U297 ( .Y(n522), .A0(n527), .A1(n528) );
  nand02 U298 ( .Y(n529), .A0(n523), .A1(n524) );
  inv01 U299 ( .Y(n527), .A(n529) );
  nand02 U300 ( .Y(n530), .A0(n525), .A1(n526) );
  inv01 U301 ( .Y(n528), .A(n530) );
  inv01 U302 ( .Y(n553), .A(n531) );
  inv01 U303 ( .Y(n532), .A(s_fract_o[18]) );
  inv01 U304 ( .Y(n533), .A(s_fract_o[19]) );
  inv01 U305 ( .Y(n534), .A(s_fract_o[1]) );
  inv01 U306 ( .Y(n535), .A(s_fract_o[20]) );
  nand02 U307 ( .Y(n531), .A0(n536), .A1(n537) );
  nand02 U308 ( .Y(n538), .A0(n532), .A1(n533) );
  inv01 U309 ( .Y(n536), .A(n538) );
  nand02 U310 ( .Y(n539), .A0(n534), .A1(n535) );
  inv01 U311 ( .Y(n537), .A(n539) );
  inv02 U312 ( .Y(U42_U3_Z_0), .A(n465) );
  inv16 U313 ( .Y(n543), .A(n466) );
  inv16 U314 ( .Y(n544), .A(n466) );
  and04 U315 ( .Y(n546), .A0(n458), .A1(n549), .A2(n550), .A3(n551) );
  and04 U316 ( .Y(n545), .A0(n460), .A1(n552), .A2(n462), .A3(n553) );
  and02 U317 ( .Y(n554), .A0(signa_i), .A1(signb_i) );
  mux21 U318 ( .Y(U42_U2_Z_9), .A0(n555), .A1(n556), .S0(n544) );
  mux21 U319 ( .Y(U42_U2_Z_8), .A0(n558), .A1(n559), .S0(n543) );
  mux21 U320 ( .Y(U42_U2_Z_7), .A0(n560), .A1(n561), .S0(n543) );
  mux21 U321 ( .Y(U42_U2_Z_6), .A0(n562), .A1(n563), .S0(n543) );
  mux21 U322 ( .Y(U42_U2_Z_5), .A0(n564), .A1(n565), .S0(n543) );
  mux21 U323 ( .Y(U42_U2_Z_4), .A0(n566), .A1(n567), .S0(n543) );
  mux21 U324 ( .Y(U42_U2_Z_3), .A0(n568), .A1(n569), .S0(n543) );
  mux21 U325 ( .Y(U42_U2_Z_27), .A0(n570), .A1(n571), .S0(n543) );
  mux21 U326 ( .Y(U42_U2_Z_26), .A0(n572), .A1(n573), .S0(n543) );
  mux21 U327 ( .Y(U42_U2_Z_25), .A0(n574), .A1(n575), .S0(n543) );
  mux21 U328 ( .Y(U42_U2_Z_24), .A0(n576), .A1(n577), .S0(n543) );
  mux21 U329 ( .Y(U42_U2_Z_23), .A0(n578), .A1(n579), .S0(n543) );
  mux21 U330 ( .Y(U42_U2_Z_22), .A0(n580), .A1(n581), .S0(n543) );
  mux21 U331 ( .Y(U42_U2_Z_21), .A0(n582), .A1(n583), .S0(n543) );
  mux21 U332 ( .Y(U42_U2_Z_20), .A0(n584), .A1(n585), .S0(n543) );
  mux21 U333 ( .Y(U42_U2_Z_2), .A0(n586), .A1(n587), .S0(n543) );
  mux21 U334 ( .Y(U42_U2_Z_19), .A0(n588), .A1(n589), .S0(n543) );
  mux21 U335 ( .Y(U42_U2_Z_18), .A0(n590), .A1(n591), .S0(n543) );
  mux21 U336 ( .Y(U42_U2_Z_17), .A0(n592), .A1(n593), .S0(n543) );
  mux21 U337 ( .Y(U42_U2_Z_16), .A0(n594), .A1(n595), .S0(n543) );
  mux21 U338 ( .Y(U42_U2_Z_15), .A0(n596), .A1(n597), .S0(n543) );
  mux21 U339 ( .Y(U42_U2_Z_14), .A0(n598), .A1(n599), .S0(n543) );
  mux21 U340 ( .Y(U42_U2_Z_13), .A0(n600), .A1(n601), .S0(n543) );
  mux21 U341 ( .Y(U42_U2_Z_12), .A0(n602), .A1(n603), .S0(n543) );
  mux21 U342 ( .Y(U42_U2_Z_11), .A0(n604), .A1(n605), .S0(n543) );
  mux21 U343 ( .Y(U42_U2_Z_10), .A0(n606), .A1(n607), .S0(n543) );
  mux21 U344 ( .Y(U42_U2_Z_1), .A0(n608), .A1(n609), .S0(n543) );
  mux21 U345 ( .Y(U42_U2_Z_0), .A0(n610), .A1(n611), .S0(n543) );
  mux21 U346 ( .Y(U42_U1_Z_9), .A0(n556), .A1(n555), .S0(n543) );
  inv01 U347 ( .Y(n555), .A(fractb_i[9]) );
  inv01 U348 ( .Y(n556), .A(fracta_i[9]) );
  mux21 U349 ( .Y(U42_U1_Z_8), .A0(n559), .A1(n558), .S0(n544) );
  inv01 U350 ( .Y(n558), .A(fractb_i[8]) );
  inv01 U351 ( .Y(n559), .A(fracta_i[8]) );
  mux21 U352 ( .Y(U42_U1_Z_7), .A0(n561), .A1(n560), .S0(n544) );
  inv01 U353 ( .Y(n560), .A(fractb_i[7]) );
  inv01 U354 ( .Y(n561), .A(fracta_i[7]) );
  mux21 U355 ( .Y(U42_U1_Z_6), .A0(n563), .A1(n562), .S0(n544) );
  inv01 U356 ( .Y(n562), .A(fractb_i[6]) );
  inv01 U357 ( .Y(n563), .A(fracta_i[6]) );
  mux21 U358 ( .Y(U42_U1_Z_5), .A0(n565), .A1(n564), .S0(n544) );
  inv01 U359 ( .Y(n564), .A(fractb_i[5]) );
  inv01 U360 ( .Y(n565), .A(fracta_i[5]) );
  mux21 U361 ( .Y(U42_U1_Z_4), .A0(n567), .A1(n566), .S0(n544) );
  inv01 U362 ( .Y(n566), .A(fractb_i[4]) );
  inv01 U363 ( .Y(n567), .A(fracta_i[4]) );
  mux21 U364 ( .Y(U42_U1_Z_3), .A0(n569), .A1(n568), .S0(n544) );
  inv01 U365 ( .Y(n568), .A(fractb_i[3]) );
  inv01 U366 ( .Y(n569), .A(fracta_i[3]) );
  mux21 U367 ( .Y(U42_U1_Z_27), .A0(n571), .A1(n570), .S0(n544) );
  inv01 U368 ( .Y(n570), .A(fractb_i[27]) );
  inv01 U369 ( .Y(n571), .A(fracta_i[27]) );
  mux21 U370 ( .Y(U42_U1_Z_26), .A0(n573), .A1(n572), .S0(n544) );
  inv01 U371 ( .Y(n572), .A(fractb_i[26]) );
  inv01 U372 ( .Y(n573), .A(fracta_i[26]) );
  mux21 U373 ( .Y(U42_U1_Z_25), .A0(n575), .A1(n574), .S0(n544) );
  inv01 U374 ( .Y(n574), .A(fractb_i[25]) );
  inv01 U375 ( .Y(n575), .A(fracta_i[25]) );
  mux21 U376 ( .Y(U42_U1_Z_24), .A0(n577), .A1(n576), .S0(n544) );
  inv01 U377 ( .Y(n576), .A(fractb_i[24]) );
  inv01 U378 ( .Y(n577), .A(fracta_i[24]) );
  mux21 U379 ( .Y(U42_U1_Z_23), .A0(n579), .A1(n578), .S0(n544) );
  inv01 U380 ( .Y(n578), .A(fractb_i[23]) );
  inv01 U381 ( .Y(n579), .A(fracta_i[23]) );
  mux21 U382 ( .Y(U42_U1_Z_22), .A0(n581), .A1(n580), .S0(n544) );
  inv01 U383 ( .Y(n580), .A(fractb_i[22]) );
  inv01 U384 ( .Y(n581), .A(fracta_i[22]) );
  mux21 U385 ( .Y(U42_U1_Z_21), .A0(n583), .A1(n582), .S0(n544) );
  inv01 U386 ( .Y(n582), .A(fractb_i[21]) );
  inv01 U387 ( .Y(n583), .A(fracta_i[21]) );
  mux21 U388 ( .Y(U42_U1_Z_20), .A0(n585), .A1(n584), .S0(n544) );
  inv01 U389 ( .Y(n584), .A(fractb_i[20]) );
  inv01 U390 ( .Y(n585), .A(fracta_i[20]) );
  mux21 U391 ( .Y(U42_U1_Z_2), .A0(n587), .A1(n586), .S0(n544) );
  inv01 U392 ( .Y(n586), .A(fractb_i[2]) );
  inv01 U393 ( .Y(n587), .A(fracta_i[2]) );
  mux21 U394 ( .Y(U42_U1_Z_19), .A0(n589), .A1(n588), .S0(n544) );
  inv01 U395 ( .Y(n588), .A(fractb_i[19]) );
  inv01 U396 ( .Y(n589), .A(fracta_i[19]) );
  mux21 U397 ( .Y(U42_U1_Z_18), .A0(n591), .A1(n590), .S0(n544) );
  inv01 U398 ( .Y(n590), .A(fractb_i[18]) );
  inv01 U399 ( .Y(n591), .A(fracta_i[18]) );
  mux21 U400 ( .Y(U42_U1_Z_17), .A0(n593), .A1(n592), .S0(n544) );
  inv01 U401 ( .Y(n592), .A(fractb_i[17]) );
  inv01 U402 ( .Y(n593), .A(fracta_i[17]) );
  mux21 U403 ( .Y(U42_U1_Z_16), .A0(n595), .A1(n594), .S0(n544) );
  inv01 U404 ( .Y(n594), .A(fractb_i[16]) );
  inv01 U405 ( .Y(n595), .A(fracta_i[16]) );
  mux21 U406 ( .Y(U42_U1_Z_15), .A0(n597), .A1(n596), .S0(n544) );
  inv01 U407 ( .Y(n596), .A(fractb_i[15]) );
  inv01 U408 ( .Y(n597), .A(fracta_i[15]) );
  mux21 U409 ( .Y(U42_U1_Z_14), .A0(n599), .A1(n598), .S0(n544) );
  inv01 U410 ( .Y(n598), .A(fractb_i[14]) );
  inv01 U411 ( .Y(n599), .A(fracta_i[14]) );
  mux21 U412 ( .Y(U42_U1_Z_13), .A0(n601), .A1(n600), .S0(n544) );
  inv01 U413 ( .Y(n600), .A(fractb_i[13]) );
  inv01 U414 ( .Y(n601), .A(fracta_i[13]) );
  mux21 U415 ( .Y(U42_U1_Z_12), .A0(n603), .A1(n602), .S0(n544) );
  inv01 U416 ( .Y(n602), .A(fractb_i[12]) );
  inv01 U417 ( .Y(n603), .A(fracta_i[12]) );
  mux21 U418 ( .Y(U42_U1_Z_11), .A0(n605), .A1(n604), .S0(n544) );
  inv01 U419 ( .Y(n604), .A(fractb_i[11]) );
  inv01 U420 ( .Y(n605), .A(fracta_i[11]) );
  mux21 U421 ( .Y(U42_U1_Z_10), .A0(n607), .A1(n606), .S0(n544) );
  inv01 U422 ( .Y(n606), .A(fractb_i[10]) );
  inv01 U423 ( .Y(n607), .A(fracta_i[10]) );
  mux21 U424 ( .Y(U42_U1_Z_1), .A0(n609), .A1(n608), .S0(n544) );
  inv01 U425 ( .Y(n608), .A(fractb_i[1]) );
  inv01 U426 ( .Y(n609), .A(fracta_i[1]) );
  mux21 U427 ( .Y(U42_U1_Z_0), .A0(n611), .A1(n610), .S0(n544) );
  nor02 U428 ( .Y(n557), .A0(n465), .A1(n____return53) );
  xor2 U429 ( .Y(n548), .A0(signb_i), .A1(fpu_op_i) );
  inv01 U430 ( .Y(n610), .A(fractb_i[0]) );
  inv01 U431 ( .Y(n611), .A(fracta_i[0]) );
  addsub_28_DW01_addsub_28_0 r272 ( .A({n521, n504, n519, n505, n509, n507, 
        n516, n496, n515, n520, n499, n508, n511, n500, n498, n495, n501, n513, 
        n512, n510, n517, n494, n502, n506, n503, n514, n518, n497}), .B({n451, 
        n426, n431, n437, n434, n440, n430, n446, n424, n445, n438, n436, n425, 
        n443, n439, n448, n429, n447, n428, n441, n435, n449, n433, n444, n432, 
        n442, n427, n450}), .CI(1'b0), .ADD_SUB(U42_U3_Z_0), .SUM(s_fract_o)
         );
  addsub_28_DW01_cmp2_28_0 gt_100_gt_gt ( .A(fractb_i), .B(fracta_i), .LEQ(
        1'b0), .TC(1'b0), .LT_LE(n____return53) );
endmodule


module post_norm_addsub_DW01_inc_9_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;
  wire   carry_8_, carry_7_, carry_6_, carry_5_, carry_4_, carry_3_, carry_2_;

  inv01 U5 ( .Y(SUM[0]), .A(A[0]) );
  xor2 U6 ( .Y(SUM[8]), .A0(carry_8_), .A1(A[8]) );
  hadd1 U1_1_1 ( .S(SUM[1]), .CO(carry_2_), .A(A[1]), .B(A[0]) );
  hadd1 U1_1_2 ( .S(SUM[2]), .CO(carry_3_), .A(A[2]), .B(carry_2_) );
  hadd1 U1_1_3 ( .S(SUM[3]), .CO(carry_4_), .A(A[3]), .B(carry_3_) );
  hadd1 U1_1_4 ( .S(SUM[4]), .CO(carry_5_), .A(A[4]), .B(carry_4_) );
  hadd1 U1_1_5 ( .S(SUM[5]), .CO(carry_6_), .A(A[5]), .B(carry_5_) );
  hadd1 U1_1_6 ( .S(SUM[6]), .CO(carry_7_), .A(A[6]), .B(carry_6_) );
  hadd1 U1_1_7 ( .S(SUM[7]), .CO(carry_8_), .A(A[7]), .B(carry_7_) );
endmodule


module post_norm_addsub_DW01_add_28_0 ( A, B, CI, SUM, CO );
  input [27:0] A;
  input [27:0] B;
  output [27:0] SUM;
  input CI;
  output CO;
  wire   carry_27_, A_2_, A_1_, A_0_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44;
  assign SUM[2] = A_2_;
  assign A_2_ = A[2];
  assign SUM[1] = A_1_;
  assign A_1_ = A[1];
  assign SUM[0] = A_0_;
  assign A_0_ = A[0];

  nand02 U4 ( .Y(n1), .A0(n34), .A1(A[5]) );
  inv02 U5 ( .Y(n2), .A(n1) );
  nand02 U6 ( .Y(n3), .A0(n20), .A1(A[12]) );
  inv02 U7 ( .Y(n4), .A(n3) );
  nand02 U8 ( .Y(n5), .A0(n26), .A1(A[14]) );
  inv02 U9 ( .Y(n6), .A(n5) );
  nand02 U10 ( .Y(n7), .A0(n36), .A1(A[22]) );
  inv02 U11 ( .Y(n8), .A(n7) );
  nand02 U12 ( .Y(n9), .A0(n42), .A1(A[20]) );
  inv02 U13 ( .Y(n10), .A(n9) );
  nand02 U14 ( .Y(n11), .A0(n30), .A1(A[16]) );
  inv02 U15 ( .Y(n12), .A(n11) );
  nand02 U16 ( .Y(n13), .A0(n40), .A1(A[18]) );
  inv02 U17 ( .Y(n14), .A(n13) );
  nand02 U18 ( .Y(n15), .A0(n32), .A1(A[7]) );
  inv02 U19 ( .Y(n16), .A(n15) );
  nand02 U20 ( .Y(n17), .A0(n38), .A1(A[24]) );
  inv02 U21 ( .Y(n18), .A(n17) );
  nand02 U22 ( .Y(n19), .A0(n24), .A1(A[11]) );
  inv02 U23 ( .Y(n20), .A(n19) );
  nand02 U24 ( .Y(n21), .A0(n28), .A1(A[9]) );
  inv02 U25 ( .Y(n22), .A(n21) );
  nand02 U26 ( .Y(n23), .A0(n22), .A1(A[10]) );
  inv02 U27 ( .Y(n24), .A(n23) );
  nand02 U28 ( .Y(n25), .A0(n4), .A1(A[13]) );
  inv02 U29 ( .Y(n26), .A(n25) );
  nand02 U30 ( .Y(n27), .A0(n16), .A1(A[8]) );
  inv02 U31 ( .Y(n28), .A(n27) );
  nand02 U32 ( .Y(n29), .A0(n6), .A1(A[15]) );
  inv02 U33 ( .Y(n30), .A(n29) );
  nand02 U34 ( .Y(n31), .A0(n2), .A1(A[6]) );
  inv02 U35 ( .Y(n32), .A(n31) );
  nand02 U36 ( .Y(n33), .A0(A[3]), .A1(A[4]) );
  inv02 U37 ( .Y(n34), .A(n33) );
  nand02 U38 ( .Y(n35), .A0(n10), .A1(A[21]) );
  inv02 U39 ( .Y(n36), .A(n35) );
  nand02 U40 ( .Y(n37), .A0(n8), .A1(A[23]) );
  inv02 U41 ( .Y(n38), .A(n37) );
  nand02 U42 ( .Y(n39), .A0(n12), .A1(A[17]) );
  inv02 U43 ( .Y(n40), .A(n39) );
  nand02 U44 ( .Y(n41), .A0(n14), .A1(A[19]) );
  inv02 U45 ( .Y(n42), .A(n41) );
  nand02 U46 ( .Y(n43), .A0(n18), .A1(A[25]) );
  inv02 U47 ( .Y(n44), .A(n43) );
  xor2 U48 ( .Y(SUM[27]), .A0(A[27]), .A1(carry_27_) );
  and02 U49 ( .Y(carry_27_), .A0(n44), .A1(A[26]) );
  xor2 U50 ( .Y(SUM[26]), .A0(A[26]), .A1(n44) );
  xor2 U51 ( .Y(SUM[25]), .A0(A[25]), .A1(n18) );
  xor2 U52 ( .Y(SUM[24]), .A0(A[24]), .A1(n38) );
  xor2 U53 ( .Y(SUM[23]), .A0(A[23]), .A1(n8) );
  xor2 U54 ( .Y(SUM[22]), .A0(A[22]), .A1(n36) );
  xor2 U55 ( .Y(SUM[21]), .A0(A[21]), .A1(n10) );
  xor2 U56 ( .Y(SUM[20]), .A0(A[20]), .A1(n42) );
  xor2 U57 ( .Y(SUM[19]), .A0(A[19]), .A1(n14) );
  xor2 U58 ( .Y(SUM[18]), .A0(A[18]), .A1(n40) );
  xor2 U59 ( .Y(SUM[17]), .A0(A[17]), .A1(n12) );
  xor2 U60 ( .Y(SUM[16]), .A0(A[16]), .A1(n30) );
  xor2 U61 ( .Y(SUM[15]), .A0(A[15]), .A1(n6) );
  xor2 U62 ( .Y(SUM[14]), .A0(A[14]), .A1(n26) );
  xor2 U63 ( .Y(SUM[13]), .A0(A[13]), .A1(n4) );
  xor2 U64 ( .Y(SUM[12]), .A0(A[12]), .A1(n20) );
  xor2 U65 ( .Y(SUM[11]), .A0(A[11]), .A1(n24) );
  xor2 U66 ( .Y(SUM[10]), .A0(A[10]), .A1(n22) );
  xor2 U67 ( .Y(SUM[9]), .A0(A[9]), .A1(n28) );
  xor2 U68 ( .Y(SUM[8]), .A0(A[8]), .A1(n16) );
  xor2 U69 ( .Y(SUM[7]), .A0(A[7]), .A1(n32) );
  xor2 U70 ( .Y(SUM[6]), .A0(A[6]), .A1(n2) );
  xor2 U71 ( .Y(SUM[5]), .A0(A[5]), .A1(n34) );
  xor2 U72 ( .Y(SUM[4]), .A0(A[4]), .A1(A[3]) );
  inv01 U73 ( .Y(SUM[3]), .A(A[3]) );
endmodule


module post_norm_addsub_DW01_dec_9_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;
  wire   carry_7_, carry_5_, carry_4_, carry_3_, n5, n7, n8, n9, n11, n13, n15,
         n17, n19, n21, n22, n23, n24, n25, n26, n27, n28;

  xor2 U6 ( .Y(n5), .A0(A[4]), .A1(n26) );
  inv01 U7 ( .Y(SUM[4]), .A(n5) );
  nor02 U8 ( .Y(n7), .A0(A[7]), .A1(n28) );
  inv02 U9 ( .Y(n8), .A(n7) );
  xor2 U10 ( .Y(n9), .A0(A[5]), .A1(n27) );
  inv01 U11 ( .Y(SUM[5]), .A(n9) );
  xor2 U12 ( .Y(n11), .A0(A[2]), .A1(n24) );
  inv01 U13 ( .Y(SUM[2]), .A(n11) );
  xor2 U14 ( .Y(n13), .A0(A[3]), .A1(n25) );
  inv01 U15 ( .Y(SUM[3]), .A(n13) );
  xor2 U16 ( .Y(n15), .A0(A[7]), .A1(n28) );
  inv01 U17 ( .Y(SUM[7]), .A(n15) );
  xor2 U18 ( .Y(n17), .A0(A[6]), .A1(n22) );
  inv01 U19 ( .Y(SUM[6]), .A(n17) );
  xor2 U20 ( .Y(n19), .A0(A[1]), .A1(A[0]) );
  inv01 U21 ( .Y(SUM[1]), .A(n19) );
  nor02 U22 ( .Y(n21), .A0(A[5]), .A1(n27) );
  inv02 U23 ( .Y(n22), .A(n21) );
  nor02 U24 ( .Y(n23), .A0(A[1]), .A1(A[0]) );
  inv02 U25 ( .Y(n24), .A(n23) );
  buf02 U26 ( .Y(n25), .A(carry_3_) );
  buf02 U27 ( .Y(n26), .A(carry_4_) );
  buf02 U28 ( .Y(n27), .A(carry_5_) );
  buf02 U29 ( .Y(n28), .A(carry_7_) );
  inv01 U30 ( .Y(SUM[0]), .A(A[0]) );
  or02 U1_B_2 ( .Y(carry_3_), .A0(A[2]), .A1(n24) );
  or02 U1_B_3 ( .Y(carry_4_), .A0(A[3]), .A1(n25) );
  or02 U1_B_4 ( .Y(carry_5_), .A0(A[4]), .A1(n26) );
  or02 U1_B_6 ( .Y(carry_7_), .A0(A[6]), .A1(n22) );
  xnor2 U1_A_8 ( .Y(SUM[8]), .A0(A[8]), .A1(n8) );
endmodule


module post_norm_addsub_DW01_dec_6_0 ( A, SUM );
  input [5:0] A;
  output [5:0] SUM;
  wire   carry_5_, carry_4_, carry_3_, carry_2_, n5, n7, n9, n11, n13, n15,
         n16, n17, n18, n19;

  xor2 U6 ( .Y(n5), .A0(A[4]), .A1(n18) );
  inv01 U7 ( .Y(SUM[4]), .A(n5) );
  xor2 U8 ( .Y(n7), .A0(carry_5_), .A1(A[5]) );
  inv01 U9 ( .Y(SUM[5]), .A(n7) );
  xor2 U10 ( .Y(n9), .A0(A[3]), .A1(n16) );
  inv01 U11 ( .Y(SUM[3]), .A(n9) );
  xor2 U12 ( .Y(n11), .A0(A[1]), .A1(A[0]) );
  inv01 U13 ( .Y(SUM[1]), .A(n11) );
  xor2 U14 ( .Y(n13), .A0(A[2]), .A1(n15) );
  inv01 U15 ( .Y(SUM[2]), .A(n13) );
  buf02 U16 ( .Y(n15), .A(carry_2_) );
  buf02 U17 ( .Y(n16), .A(carry_3_) );
  inv01 U18 ( .Y(n17), .A(carry_4_) );
  inv01 U19 ( .Y(n18), .A(n17) );
  inv01 U20 ( .Y(n19), .A(n17) );
  inv01 U21 ( .Y(SUM[0]), .A(A[0]) );
  or02 U1_B_1 ( .Y(carry_2_), .A0(A[1]), .A1(A[0]) );
  or02 U1_B_2 ( .Y(carry_3_), .A0(A[2]), .A1(n15) );
  or02 U1_B_3 ( .Y(carry_4_), .A0(A[3]), .A1(n16) );
  or02 U1_B_4 ( .Y(carry_5_), .A0(A[4]), .A1(n19) );
endmodule


module post_norm_addsub ( clk_i, opa_i, opb_i, fract_28_i, exp_i, sign_i, 
        fpu_op_i, rmode_i, output_o, ine_o );
  input [31:0] opa_i;
  input [31:0] opb_i;
  input [27:0] fract_28_i;
  input [7:0] exp_i;
  input [1:0] rmode_i;
  output [31:0] output_o;
  input clk_i, sign_i, fpu_op_i;
  output ine_o;
  wire   s_ine_o, s_shr1_5_, s_shr1_4_, s_shr1_3_, s_shr1_2_, s_shr1_1_,
         s_shr1_0_, s_shl11786_5_, s_shl11786_4_, s_shl11786_3_, s_shl11786_2_,
         s_shl11786_1_, s_shl11786_0_, s_shl1_4_, s_shl1_3_, s_shl1_2_,
         s_shl1_1_, s_shl1_0_, s_expo9_11794_6_, s_expo9_11794_5_,
         s_expo9_11794_4_, s_expo9_11794_3_, s_expo9_11794_2_,
         s_expo9_11794_1_, s_expo9_11794_0_, n____return1927_5_,
         n____return1927_4_, n____return1927_3_, n____return1927_2_,
         n____return1927_1_, n____return1927_0_, s_fracto28_12090_27_,
         s_fracto28_12090_26_, s_fracto28_12090_25_, s_fracto28_12090_24_,
         s_fracto28_12090_23_, s_fracto28_12090_22_, s_fracto28_12090_21_,
         s_fracto28_12090_20_, s_fracto28_12090_19_, s_fracto28_12090_18_,
         s_fracto28_12090_17_, s_fracto28_12090_16_, s_fracto28_12090_15_,
         s_fracto28_12090_14_, s_fracto28_12090_13_, s_fracto28_12090_12_,
         s_fracto28_12090_11_, s_fracto28_12090_10_, s_fracto28_12090_9_,
         s_fracto28_12090_8_, s_fracto28_12090_7_, s_fracto28_12090_6_,
         s_fracto28_12090_5_, s_fracto28_12090_4_, s_fracto28_12090_3_,
         s_fracto28_12090_2_, s_fracto28_12090_1_, s_fracto28_12090_0_,
         n2550_8_, n____return2548_7_, n____return2548_6_, n____return2548_5_,
         n____return2548_4_, n____return2548_3_, n____return2548_2_,
         n____return2548_1_, n____return2548_0_, n2768_27_,
         n____return2766_26_, n____return2766_25_, n____return2766_24_,
         n____return2766_23_, n____return2766_22_, n____return2766_21_,
         n____return2766_20_, n____return2766_19_, n____return2766_18_,
         n____return2766_17_, n____return2766_16_, n____return2766_15_,
         n____return2766_14_, n____return2766_13_, n____return2766_12_,
         n____return2766_11_, n____return2766_10_, n____return2766_9_,
         n____return2766_8_, n____return2766_7_, n____return2766_6_,
         n____return2766_5_, n____return2766_4_, n____return2766_3_,
         n____return2766_2_, n____return2766_1_, n____return2766_0_, n2866_8_,
         n____return2864_7_, n____return2864_6_, n____return2864_5_,
         n____return2864_4_, n____return2864_3_, n____return2864_2_,
         n____return2864_1_, n____return2864_0_, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114;
  wire   [31:0] s_output_o;
  wire   [8:0] s_expo9_1;
  wire   [27:0] s_fracto28_1;
  wire   [8:0] s_expo9_2;

  dff s_expo9_1_reg_8_ ( .Q(s_expo9_1[8]), .D(1'b0), .CLK(clk_i) );
  dff s_shr1_reg_5_ ( .Q(s_shr1_5_), .D(1'b0), .CLK(clk_i) );
  dff s_shr1_reg_4_ ( .Q(s_shr1_4_), .D(1'b0), .CLK(clk_i) );
  dff s_shr1_reg_3_ ( .Q(s_shr1_3_), .D(1'b0), .CLK(clk_i) );
  dff s_shr1_reg_2_ ( .Q(s_shr1_2_), .D(1'b0), .CLK(clk_i) );
  dff s_shr1_reg_1_ ( .Q(s_shr1_1_), .D(1'b0), .CLK(clk_i) );
  dff s_shl1_reg_5_ ( .QB(n8114), .D(s_shl11786_5_), .CLK(clk_i) );
  dff s_shl1_reg_4_ ( .Q(s_shl1_4_), .D(s_shl11786_4_), .CLK(clk_i) );
  dff s_shl1_reg_3_ ( .Q(s_shl1_3_), .D(s_shl11786_3_), .CLK(clk_i) );
  dff s_shl1_reg_2_ ( .Q(s_shl1_2_), .D(s_shl11786_2_), .CLK(clk_i) );
  dff s_shl1_reg_1_ ( .Q(s_shl1_1_), .D(s_shl11786_1_), .CLK(clk_i) );
  dff s_shl1_reg_0_ ( .Q(s_shl1_0_), .D(s_shl11786_0_), .CLK(clk_i) );
  dff s_expo9_1_reg_7_ ( .Q(s_expo9_1[7]), .D(n6969), .CLK(clk_i) );
  dff s_expo9_1_reg_6_ ( .Q(s_expo9_1[6]), .D(s_expo9_11794_6_), .CLK(clk_i)
         );
  dff s_expo9_1_reg_5_ ( .Q(s_expo9_1[5]), .D(s_expo9_11794_5_), .CLK(clk_i)
         );
  dff s_expo9_1_reg_4_ ( .Q(s_expo9_1[4]), .D(s_expo9_11794_4_), .CLK(clk_i)
         );
  dff s_expo9_1_reg_3_ ( .Q(s_expo9_1[3]), .D(s_expo9_11794_3_), .CLK(clk_i)
         );
  dff s_expo9_1_reg_2_ ( .Q(s_expo9_1[2]), .D(s_expo9_11794_2_), .CLK(clk_i)
         );
  dff s_expo9_1_reg_1_ ( .Q(s_expo9_1[1]), .D(s_expo9_11794_1_), .CLK(clk_i)
         );
  dff s_expo9_1_reg_0_ ( .Q(s_expo9_1[0]), .D(s_expo9_11794_0_), .CLK(clk_i)
         );
  dff s_fracto28_1_reg_27_ ( .Q(s_fracto28_1[27]), .D(s_fracto28_12090_27_), 
        .CLK(clk_i) );
  dff s_fracto28_1_reg_26_ ( .Q(s_fracto28_1[26]), .D(s_fracto28_12090_26_), 
        .CLK(clk_i) );
  dff s_fracto28_1_reg_25_ ( .Q(s_fracto28_1[25]), .D(s_fracto28_12090_25_), 
        .CLK(clk_i) );
  dff s_fracto28_1_reg_24_ ( .Q(s_fracto28_1[24]), .D(s_fracto28_12090_24_), 
        .CLK(clk_i) );
  dff s_fracto28_1_reg_23_ ( .Q(s_fracto28_1[23]), .D(s_fracto28_12090_23_), 
        .CLK(clk_i) );
  dff s_fracto28_1_reg_22_ ( .Q(s_fracto28_1[22]), .D(n4491), .CLK(clk_i) );
  dff s_fracto28_1_reg_21_ ( .Q(s_fracto28_1[21]), .D(n4495), .CLK(clk_i) );
  dff s_fracto28_1_reg_20_ ( .Q(s_fracto28_1[20]), .D(s_fracto28_12090_20_), 
        .CLK(clk_i) );
  dff s_fracto28_1_reg_19_ ( .Q(s_fracto28_1[19]), .D(s_fracto28_12090_19_), 
        .CLK(clk_i) );
  dff s_fracto28_1_reg_18_ ( .Q(s_fracto28_1[18]), .D(s_fracto28_12090_18_), 
        .CLK(clk_i) );
  dff s_fracto28_1_reg_17_ ( .Q(s_fracto28_1[17]), .D(s_fracto28_12090_17_), 
        .CLK(clk_i) );
  dff s_fracto28_1_reg_16_ ( .Q(s_fracto28_1[16]), .D(s_fracto28_12090_16_), 
        .CLK(clk_i) );
  dff s_fracto28_1_reg_15_ ( .Q(s_fracto28_1[15]), .D(s_fracto28_12090_15_), 
        .CLK(clk_i) );
  dff s_fracto28_1_reg_14_ ( .Q(s_fracto28_1[14]), .D(n4492), .CLK(clk_i) );
  dff s_fracto28_1_reg_13_ ( .Q(s_fracto28_1[13]), .D(s_fracto28_12090_13_), 
        .CLK(clk_i) );
  dff s_fracto28_1_reg_12_ ( .Q(s_fracto28_1[12]), .D(s_fracto28_12090_12_), 
        .CLK(clk_i) );
  dff s_fracto28_1_reg_11_ ( .Q(s_fracto28_1[11]), .D(s_fracto28_12090_11_), 
        .CLK(clk_i) );
  dff s_fracto28_1_reg_10_ ( .Q(s_fracto28_1[10]), .D(s_fracto28_12090_10_), 
        .CLK(clk_i) );
  dff s_fracto28_1_reg_9_ ( .Q(s_fracto28_1[9]), .D(s_fracto28_12090_9_), 
        .CLK(clk_i) );
  dff s_fracto28_1_reg_8_ ( .Q(s_fracto28_1[8]), .D(s_fracto28_12090_8_), 
        .CLK(clk_i) );
  dff s_fracto28_1_reg_7_ ( .Q(s_fracto28_1[7]), .D(s_fracto28_12090_7_), 
        .CLK(clk_i) );
  dff s_fracto28_1_reg_6_ ( .Q(s_fracto28_1[6]), .D(n4490), .CLK(clk_i) );
  dff s_fracto28_1_reg_5_ ( .Q(s_fracto28_1[5]), .D(s_fracto28_12090_5_), 
        .CLK(clk_i) );
  dff s_fracto28_1_reg_4_ ( .Q(s_fracto28_1[4]), .D(s_fracto28_12090_4_), 
        .CLK(clk_i) );
  dff s_fracto28_1_reg_3_ ( .Q(s_fracto28_1[3]), .D(s_fracto28_12090_3_), 
        .CLK(clk_i) );
  dff s_fracto28_1_reg_2_ ( .Q(s_fracto28_1[2]), .D(s_fracto28_12090_2_), 
        .CLK(clk_i) );
  dff s_fracto28_1_reg_1_ ( .Q(s_fracto28_1[1]), .D(s_fracto28_12090_1_), 
        .CLK(clk_i) );
  dff s_fracto28_1_reg_0_ ( .Q(s_fracto28_1[0]), .D(s_fracto28_12090_0_), 
        .CLK(clk_i) );
  dff output_o_reg_31_ ( .Q(output_o[31]), .D(s_output_o[31]), .CLK(clk_i) );
  dff output_o_reg_30_ ( .Q(output_o[30]), .D(s_output_o[30]), .CLK(clk_i) );
  dff output_o_reg_29_ ( .Q(output_o[29]), .D(s_output_o[29]), .CLK(clk_i) );
  dff output_o_reg_28_ ( .Q(output_o[28]), .D(s_output_o[28]), .CLK(clk_i) );
  dff output_o_reg_27_ ( .Q(output_o[27]), .D(s_output_o[27]), .CLK(clk_i) );
  dff output_o_reg_26_ ( .Q(output_o[26]), .D(s_output_o[26]), .CLK(clk_i) );
  dff output_o_reg_25_ ( .Q(output_o[25]), .D(s_output_o[25]), .CLK(clk_i) );
  dff output_o_reg_24_ ( .Q(output_o[24]), .D(s_output_o[24]), .CLK(clk_i) );
  dff output_o_reg_23_ ( .Q(output_o[23]), .D(s_output_o[23]), .CLK(clk_i) );
  dff output_o_reg_22_ ( .Q(output_o[22]), .D(s_output_o[22]), .CLK(clk_i) );
  dff output_o_reg_21_ ( .Q(output_o[21]), .D(s_output_o[21]), .CLK(clk_i) );
  dff output_o_reg_20_ ( .Q(output_o[20]), .D(s_output_o[20]), .CLK(clk_i) );
  dff output_o_reg_19_ ( .Q(output_o[19]), .D(s_output_o[19]), .CLK(clk_i) );
  dff output_o_reg_18_ ( .Q(output_o[18]), .D(s_output_o[18]), .CLK(clk_i) );
  dff output_o_reg_17_ ( .Q(output_o[17]), .D(s_output_o[17]), .CLK(clk_i) );
  dff output_o_reg_16_ ( .Q(output_o[16]), .D(s_output_o[16]), .CLK(clk_i) );
  dff output_o_reg_15_ ( .Q(output_o[15]), .D(s_output_o[15]), .CLK(clk_i) );
  dff output_o_reg_14_ ( .Q(output_o[14]), .D(s_output_o[14]), .CLK(clk_i) );
  dff output_o_reg_13_ ( .Q(output_o[13]), .D(s_output_o[13]), .CLK(clk_i) );
  dff output_o_reg_12_ ( .Q(output_o[12]), .D(s_output_o[12]), .CLK(clk_i) );
  dff output_o_reg_11_ ( .Q(output_o[11]), .D(s_output_o[11]), .CLK(clk_i) );
  dff output_o_reg_10_ ( .Q(output_o[10]), .D(s_output_o[10]), .CLK(clk_i) );
  dff output_o_reg_9_ ( .Q(output_o[9]), .D(s_output_o[9]), .CLK(clk_i) );
  dff output_o_reg_8_ ( .Q(output_o[8]), .D(s_output_o[8]), .CLK(clk_i) );
  dff output_o_reg_7_ ( .Q(output_o[7]), .D(s_output_o[7]), .CLK(clk_i) );
  dff output_o_reg_6_ ( .Q(output_o[6]), .D(s_output_o[6]), .CLK(clk_i) );
  dff output_o_reg_5_ ( .Q(output_o[5]), .D(s_output_o[5]), .CLK(clk_i) );
  dff output_o_reg_4_ ( .Q(output_o[4]), .D(s_output_o[4]), .CLK(clk_i) );
  dff output_o_reg_3_ ( .Q(output_o[3]), .D(s_output_o[3]), .CLK(clk_i) );
  dff output_o_reg_2_ ( .Q(output_o[2]), .D(s_output_o[2]), .CLK(clk_i) );
  dff output_o_reg_1_ ( .Q(output_o[1]), .D(s_output_o[1]), .CLK(clk_i) );
  dff output_o_reg_0_ ( .Q(output_o[0]), .D(s_output_o[0]), .CLK(clk_i) );
  dff ine_o_reg ( .Q(ine_o), .D(s_ine_o), .CLK(clk_i) );
  dff s_shr1_reg_0_ ( .Q(s_shr1_0_), .D(n4317), .CLK(clk_i) );
  xor2 U1308 ( .Y(n4246), .A0(n8048), .A1(exp_i[2]) );
  inv01 U1309 ( .Y(n4247), .A(n4246) );
  ao22 U1310 ( .Y(n4248), .A0(n7692), .A1(fract_28_i[1]), .B0(n7695), .B1(
        fract_28_i[4]) );
  inv01 U1311 ( .Y(n4249), .A(n4248) );
  ao21 U1312 ( .Y(n4250), .A0(n7810), .A1(n7811), .B0(n4261) );
  inv01 U1313 ( .Y(n4251), .A(n4250) );
  ao22 U1314 ( .Y(n4252), .A0(n7694), .A1(fract_28_i[2]), .B0(n7695), .B1(
        fract_28_i[5]) );
  inv01 U1315 ( .Y(n4253), .A(n4252) );
  inv01 U1316 ( .Y(n7851), .A(n4254) );
  nor02 U1317 ( .Y(n4255), .A0(n7988), .A1(n7900) );
  nor02 U1318 ( .Y(n4256), .A0(n7704), .A1(n7881) );
  nor02 U1319 ( .Y(n4254), .A0(n4255), .A1(n4256) );
  inv02 U1320 ( .Y(n7805), .A(s_shr1_0_) );
  inv01 U1321 ( .Y(n4257), .A(n4579) );
  ao22 U1322 ( .Y(n4258), .A0(n7693), .A1(fract_28_i[3]), .B0(n7695), .B1(
        fract_28_i[6]) );
  inv01 U1323 ( .Y(n4259), .A(n4258) );
  xor2 U1324 ( .Y(n4260), .A0(n7728), .A1(rmode_i[0]) );
  inv01 U1325 ( .Y(n4261), .A(n4260) );
  ao22 U1326 ( .Y(n4262), .A0(n7693), .A1(fract_28_i[0]), .B0(n7695), .B1(
        fract_28_i[3]) );
  inv01 U1327 ( .Y(n4263), .A(n4262) );
  ao22 U1328 ( .Y(n4264), .A0(n7806), .A1(n7788), .B0(n5953), .B1(n7787) );
  inv01 U1329 ( .Y(n4265), .A(n4264) );
  ao22 U1330 ( .Y(n4266), .A0(n7678), .A1(n7924), .B0(n7675), .B1(n7823) );
  inv01 U1331 ( .Y(n4267), .A(n4266) );
  ao22 U1332 ( .Y(n4268), .A0(n7672), .A1(n7827), .B0(n7670), .B1(n7823) );
  inv01 U1333 ( .Y(n4269), .A(n4268) );
  ao22 U1334 ( .Y(n4270), .A0(fract_28_i[24]), .A1(n7689), .B0(n7679), .B1(
        fract_28_i[25]) );
  inv01 U1335 ( .Y(n4271), .A(n4270) );
  nand02 U1336 ( .Y(n8010), .A0(n4272), .A1(n4273) );
  inv01 U1337 ( .Y(n4274), .A(fract_28_i[5]) );
  inv01 U1338 ( .Y(n4275), .A(fract_28_i[4]) );
  inv01 U1339 ( .Y(n4276), .A(n7690) );
  inv01 U1340 ( .Y(n4277), .A(n7679) );
  nand02 U1341 ( .Y(n4278), .A0(n4274), .A1(n4275) );
  nand02 U1342 ( .Y(n4279), .A0(n4274), .A1(n4276) );
  nand02 U1343 ( .Y(n4280), .A0(n4275), .A1(n4277) );
  nand02 U1344 ( .Y(n4281), .A0(n4276), .A1(n4277) );
  nand02 U1345 ( .Y(n4282), .A0(n4278), .A1(n4279) );
  inv01 U1346 ( .Y(n4272), .A(n4282) );
  nand02 U1347 ( .Y(n4283), .A0(n4280), .A1(n4281) );
  inv01 U1348 ( .Y(n4273), .A(n4283) );
  ao22 U1349 ( .Y(n4284), .A0(n7694), .A1(fract_28_i[4]), .B0(n7695), .B1(
        fract_28_i[7]) );
  inv01 U1350 ( .Y(n4285), .A(n4284) );
  nand02 U1351 ( .Y(n7994), .A0(n4286), .A1(n4287) );
  inv01 U1352 ( .Y(n4288), .A(fract_28_i[16]) );
  inv01 U1353 ( .Y(n4289), .A(fract_28_i[15]) );
  inv01 U1354 ( .Y(n4290), .A(n7689) );
  inv01 U1355 ( .Y(n4291), .A(n7679) );
  nand02 U1356 ( .Y(n4292), .A0(n4288), .A1(n4289) );
  nand02 U1357 ( .Y(n4293), .A0(n4288), .A1(n4290) );
  nand02 U1358 ( .Y(n4294), .A0(n4289), .A1(n4291) );
  nand02 U1359 ( .Y(n4295), .A0(n4290), .A1(n4291) );
  nand02 U1360 ( .Y(n4296), .A0(n4292), .A1(n4293) );
  inv01 U1361 ( .Y(n4286), .A(n4296) );
  nand02 U1362 ( .Y(n4297), .A0(n4294), .A1(n4295) );
  inv01 U1363 ( .Y(n4287), .A(n4297) );
  ao22 U1364 ( .Y(n4298), .A0(n7694), .A1(fract_28_i[15]), .B0(n7695), .B1(
        fract_28_i[18]) );
  inv01 U1365 ( .Y(n4299), .A(n4298) );
  nand02 U1366 ( .Y(n7877), .A0(n4300), .A1(n4301) );
  inv01 U1367 ( .Y(n4302), .A(fract_28_i[8]) );
  inv01 U1368 ( .Y(n4303), .A(fract_28_i[7]) );
  inv01 U1369 ( .Y(n4304), .A(n7689) );
  inv01 U1370 ( .Y(n4305), .A(n7679) );
  nand02 U1371 ( .Y(n4306), .A0(n4302), .A1(n4303) );
  nand02 U1372 ( .Y(n4307), .A0(n4302), .A1(n4304) );
  nand02 U1373 ( .Y(n4308), .A0(n4303), .A1(n4305) );
  nand02 U1374 ( .Y(n4309), .A0(n4304), .A1(n4305) );
  nand02 U1375 ( .Y(n4310), .A0(n4306), .A1(n4307) );
  inv01 U1376 ( .Y(n4300), .A(n4310) );
  nand02 U1377 ( .Y(n4311), .A0(n4308), .A1(n4309) );
  inv01 U1378 ( .Y(n4301), .A(n4311) );
  ao22 U1379 ( .Y(n4312), .A0(n7693), .A1(fract_28_i[7]), .B0(n7695), .B1(
        fract_28_i[10]) );
  inv01 U1380 ( .Y(n4313), .A(n4312) );
  ao22 U1381 ( .Y(n4314), .A0(n7689), .A1(fract_28_i[14]), .B0(n7679), .B1(
        fract_28_i[15]) );
  inv01 U1382 ( .Y(n4315), .A(n4314) );
  or02 U1383 ( .Y(n4316), .A0(n7704), .A1(n4707) );
  inv01 U1384 ( .Y(n4317), .A(n4316) );
  nand02 U1385 ( .Y(n8000), .A0(n4318), .A1(n4319) );
  inv01 U1386 ( .Y(n4320), .A(fract_28_i[23]) );
  inv01 U1387 ( .Y(n4321), .A(fract_28_i[22]) );
  inv01 U1388 ( .Y(n4322), .A(n7689) );
  inv01 U1389 ( .Y(n4323), .A(n7679) );
  nand02 U1390 ( .Y(n4324), .A0(n4320), .A1(n4321) );
  nand02 U1391 ( .Y(n4325), .A0(n4320), .A1(n4322) );
  nand02 U1392 ( .Y(n4326), .A0(n4321), .A1(n4323) );
  nand02 U1393 ( .Y(n4327), .A0(n4322), .A1(n4323) );
  nand02 U1394 ( .Y(n4328), .A0(n4324), .A1(n4325) );
  inv01 U1395 ( .Y(n4318), .A(n4328) );
  nand02 U1396 ( .Y(n4329), .A0(n4326), .A1(n4327) );
  inv01 U1397 ( .Y(n4319), .A(n4329) );
  ao22 U1398 ( .Y(n4330), .A0(n7692), .A1(fract_28_i[22]), .B0(n7695), .B1(
        fract_28_i[25]) );
  inv01 U1399 ( .Y(n4331), .A(n4330) );
  nand02 U1400 ( .Y(n7975), .A0(n4332), .A1(n4333) );
  inv01 U1401 ( .Y(n4334), .A(fract_28_i[16]) );
  inv01 U1402 ( .Y(n4335), .A(fract_28_i[13]) );
  inv01 U1403 ( .Y(n4336), .A(n7692) );
  inv01 U1404 ( .Y(n4337), .A(n7695) );
  nand02 U1405 ( .Y(n4338), .A0(n4334), .A1(n4335) );
  nand02 U1406 ( .Y(n4339), .A0(n4334), .A1(n4336) );
  nand02 U1407 ( .Y(n4340), .A0(n4335), .A1(n4337) );
  nand02 U1408 ( .Y(n4341), .A0(n4336), .A1(n4337) );
  nand02 U1409 ( .Y(n4342), .A0(n4338), .A1(n4339) );
  inv01 U1410 ( .Y(n4332), .A(n4342) );
  nand02 U1411 ( .Y(n4343), .A0(n4340), .A1(n4341) );
  inv01 U1412 ( .Y(n4333), .A(n4343) );
  ao22 U1413 ( .Y(n4344), .A0(n7690), .A1(fract_28_i[13]), .B0(n7679), .B1(
        fract_28_i[14]) );
  inv01 U1414 ( .Y(n4345), .A(n4344) );
  ao22 U1415 ( .Y(n4346), .A0(n7690), .A1(fract_28_i[18]), .B0(n7679), .B1(
        fract_28_i[19]) );
  inv01 U1416 ( .Y(n4347), .A(n4346) );
  ao22 U1417 ( .Y(n4348), .A0(n7694), .A1(fract_28_i[18]), .B0(n7695), .B1(
        fract_28_i[21]) );
  inv01 U1418 ( .Y(n4349), .A(n4348) );
  nand02 U1419 ( .Y(n7999), .A0(n4350), .A1(n4351) );
  inv01 U1420 ( .Y(n4352), .A(fract_28_i[11]) );
  inv01 U1421 ( .Y(n4353), .A(fract_28_i[10]) );
  inv01 U1422 ( .Y(n4354), .A(n7689) );
  inv01 U1423 ( .Y(n4355), .A(n7422) );
  nand02 U1424 ( .Y(n4356), .A0(n4352), .A1(n4353) );
  nand02 U1425 ( .Y(n4357), .A0(n4352), .A1(n4354) );
  nand02 U1426 ( .Y(n4358), .A0(n4353), .A1(n4355) );
  nand02 U1427 ( .Y(n4359), .A0(n4354), .A1(n4355) );
  nand02 U1428 ( .Y(n4360), .A0(n4356), .A1(n4357) );
  inv01 U1429 ( .Y(n4350), .A(n4360) );
  nand02 U1430 ( .Y(n4361), .A0(n4358), .A1(n4359) );
  inv01 U1431 ( .Y(n4351), .A(n4361) );
  ao22 U1432 ( .Y(n4362), .A0(n7693), .A1(fract_28_i[10]), .B0(n7695), .B1(
        fract_28_i[13]) );
  inv01 U1433 ( .Y(n4363), .A(n4362) );
  ao22 U1434 ( .Y(n4364), .A0(n7692), .A1(fract_28_i[8]), .B0(n7695), .B1(
        fract_28_i[11]) );
  inv01 U1435 ( .Y(n4365), .A(n4364) );
  ao22 U1436 ( .Y(n4366), .A0(n7690), .A1(fract_28_i[8]), .B0(n7679), .B1(
        fract_28_i[9]) );
  inv01 U1437 ( .Y(n4367), .A(n4366) );
  nand02 U1438 ( .Y(n7983), .A0(n4368), .A1(n4369) );
  inv01 U1439 ( .Y(n4370), .A(fract_28_i[14]) );
  inv01 U1440 ( .Y(n4371), .A(fract_28_i[11]) );
  inv01 U1441 ( .Y(n4372), .A(n7692) );
  inv01 U1442 ( .Y(n4373), .A(n7695) );
  nand02 U1443 ( .Y(n4374), .A0(n4370), .A1(n4371) );
  nand02 U1444 ( .Y(n4375), .A0(n4370), .A1(n4372) );
  nand02 U1445 ( .Y(n4376), .A0(n4371), .A1(n4373) );
  nand02 U1446 ( .Y(n4377), .A0(n4372), .A1(n4373) );
  nand02 U1447 ( .Y(n4378), .A0(n4374), .A1(n4375) );
  inv01 U1448 ( .Y(n4368), .A(n4378) );
  nand02 U1449 ( .Y(n4379), .A0(n4376), .A1(n4377) );
  inv01 U1450 ( .Y(n4369), .A(n4379) );
  ao22 U1451 ( .Y(n4380), .A0(n7689), .A1(fract_28_i[5]), .B0(n7679), .B1(
        fract_28_i[6]) );
  inv01 U1452 ( .Y(n4381), .A(n4380) );
  ao22 U1453 ( .Y(n4382), .A0(n7694), .A1(fract_28_i[14]), .B0(n7695), .B1(
        fract_28_i[17]) );
  inv01 U1454 ( .Y(n4383), .A(n4382) );
  ao22 U1455 ( .Y(n4384), .A0(n7690), .A1(fract_28_i[16]), .B0(n7679), .B1(
        fract_28_i[17]) );
  inv01 U1456 ( .Y(n4385), .A(n4384) );
  ao22 U1457 ( .Y(n4386), .A0(n7690), .A1(fract_28_i[11]), .B0(n7679), .B1(
        fract_28_i[12]) );
  inv01 U1458 ( .Y(n4387), .A(n4386) );
  ao22 U1459 ( .Y(n4388), .A0(n7694), .A1(fract_28_i[5]), .B0(n7695), .B1(
        fract_28_i[8]) );
  inv01 U1460 ( .Y(n4389), .A(n4388) );
  ao22 U1461 ( .Y(n4390), .A0(n7694), .A1(fract_28_i[16]), .B0(n7695), .B1(
        fract_28_i[19]) );
  inv01 U1462 ( .Y(n4391), .A(n4390) );
  inv01 U1463 ( .Y(n8050), .A(n4392) );
  nor02 U1464 ( .Y(n4393), .A0(n8034), .A1(n8033) );
  inv01 U1465 ( .Y(n4394), .A(n7191) );
  nor02 U1466 ( .Y(n4392), .A0(n4393), .A1(n4394) );
  ao22 U1467 ( .Y(n4395), .A0(n7690), .A1(fract_28_i[19]), .B0(n7679), .B1(
        fract_28_i[20]) );
  inv01 U1468 ( .Y(n4396), .A(n4395) );
  nand02 U1469 ( .Y(n7888), .A0(n4397), .A1(n4398) );
  inv01 U1470 ( .Y(n4399), .A(fract_28_i[7]) );
  inv01 U1471 ( .Y(n4400), .A(fract_28_i[6]) );
  inv01 U1472 ( .Y(n4401), .A(n7689) );
  inv01 U1473 ( .Y(n4402), .A(n7679) );
  nand02 U1474 ( .Y(n4403), .A0(n4399), .A1(n4400) );
  nand02 U1475 ( .Y(n4404), .A0(n4399), .A1(n4401) );
  nand02 U1476 ( .Y(n4405), .A0(n4400), .A1(n4402) );
  nand02 U1477 ( .Y(n4406), .A0(n4401), .A1(n4402) );
  nand02 U1478 ( .Y(n4407), .A0(n4403), .A1(n4404) );
  inv01 U1479 ( .Y(n4397), .A(n4407) );
  nand02 U1480 ( .Y(n4408), .A0(n4405), .A1(n4406) );
  inv01 U1481 ( .Y(n4398), .A(n4408) );
  ao22 U1482 ( .Y(n4409), .A0(n7692), .A1(fract_28_i[6]), .B0(n7695), .B1(
        fract_28_i[9]) );
  inv01 U1483 ( .Y(n4410), .A(n4409) );
  ao22 U1484 ( .Y(n4411), .A0(n7689), .A1(fract_28_i[12]), .B0(n7679), .B1(
        fract_28_i[13]) );
  inv01 U1485 ( .Y(n4412), .A(n4411) );
  ao22 U1486 ( .Y(n4413), .A0(n7689), .A1(fract_28_i[9]), .B0(n7679), .B1(
        fract_28_i[10]) );
  inv01 U1487 ( .Y(n4414), .A(n4413) );
  ao22 U1488 ( .Y(n4415), .A0(n7692), .A1(fract_28_i[19]), .B0(n7695), .B1(
        fract_28_i[22]) );
  inv01 U1489 ( .Y(n4416), .A(n4415) );
  ao22 U1490 ( .Y(n4417), .A0(n7694), .A1(fract_28_i[12]), .B0(n7695), .B1(
        fract_28_i[15]) );
  inv01 U1491 ( .Y(n4418), .A(n4417) );
  ao22 U1492 ( .Y(n4419), .A0(n7693), .A1(fract_28_i[9]), .B0(n7695), .B1(
        fract_28_i[12]) );
  inv01 U1493 ( .Y(n4420), .A(n4419) );
  nand02 U1494 ( .Y(n8013), .A0(n4421), .A1(n4422) );
  inv01 U1495 ( .Y(n4423), .A(fract_28_i[21]) );
  inv01 U1496 ( .Y(n4424), .A(fract_28_i[20]) );
  inv01 U1497 ( .Y(n4425), .A(n7690) );
  inv01 U1498 ( .Y(n4426), .A(n7679) );
  nand02 U1499 ( .Y(n4427), .A0(n4423), .A1(n4424) );
  nand02 U1500 ( .Y(n4428), .A0(n4423), .A1(n4425) );
  nand02 U1501 ( .Y(n4429), .A0(n4424), .A1(n4426) );
  nand02 U1502 ( .Y(n4430), .A0(n4425), .A1(n4426) );
  nand02 U1503 ( .Y(n4431), .A0(n4427), .A1(n4428) );
  inv01 U1504 ( .Y(n4421), .A(n4431) );
  nand02 U1505 ( .Y(n4432), .A0(n4429), .A1(n4430) );
  inv01 U1506 ( .Y(n4422), .A(n4432) );
  ao22 U1507 ( .Y(n4433), .A0(n7694), .A1(fract_28_i[20]), .B0(n7695), .B1(
        fract_28_i[23]) );
  inv01 U1508 ( .Y(n4434), .A(n4433) );
  ao22 U1509 ( .Y(n4435), .A0(fract_28_i[24]), .A1(n7693), .B0(n7695), .B1(
        fract_28_i[27]) );
  inv01 U1510 ( .Y(n4436), .A(n4435) );
  nand02 U1511 ( .Y(n7950), .A0(n4437), .A1(n4438) );
  inv01 U1512 ( .Y(n4439), .A(fract_28_i[20]) );
  inv01 U1513 ( .Y(n4440), .A(fract_28_i[17]) );
  inv01 U1514 ( .Y(n4441), .A(n7692) );
  inv01 U1515 ( .Y(n4442), .A(n7695) );
  nand02 U1516 ( .Y(n4443), .A0(n4439), .A1(n4440) );
  nand02 U1517 ( .Y(n4444), .A0(n4439), .A1(n4441) );
  nand02 U1518 ( .Y(n4445), .A0(n4440), .A1(n4442) );
  nand02 U1519 ( .Y(n4446), .A0(n4441), .A1(n4442) );
  nand02 U1520 ( .Y(n4447), .A0(n4443), .A1(n4444) );
  inv01 U1521 ( .Y(n4437), .A(n4447) );
  nand02 U1522 ( .Y(n4448), .A0(n4445), .A1(n4446) );
  inv01 U1523 ( .Y(n4438), .A(n4448) );
  ao22 U1524 ( .Y(n4449), .A0(n7690), .A1(fract_28_i[17]), .B0(n7679), .B1(
        fract_28_i[18]) );
  inv01 U1525 ( .Y(n4450), .A(n4449) );
  nand02 U1526 ( .Y(n7933), .A0(n4451), .A1(n4452) );
  inv01 U1527 ( .Y(n4453), .A(n7695) );
  inv01 U1528 ( .Y(n4454), .A(fract_28_i[21]) );
  inv01 U1529 ( .Y(n4455), .A(n7693) );
  inv01 U1530 ( .Y(n4456), .A(fract_28_i[24]) );
  nand02 U1531 ( .Y(n4457), .A0(n4453), .A1(n4454) );
  nand02 U1532 ( .Y(n4458), .A0(n4453), .A1(n4455) );
  nand02 U1533 ( .Y(n4459), .A0(n4454), .A1(n4456) );
  nand02 U1534 ( .Y(n4460), .A0(n4455), .A1(n4456) );
  nand02 U1535 ( .Y(n4461), .A0(n4457), .A1(n4458) );
  inv01 U1536 ( .Y(n4451), .A(n4461) );
  nand02 U1537 ( .Y(n4462), .A0(n4459), .A1(n4460) );
  inv01 U1538 ( .Y(n4452), .A(n4462) );
  ao22 U1539 ( .Y(n4463), .A0(n7690), .A1(fract_28_i[21]), .B0(n7679), .B1(
        fract_28_i[22]) );
  inv01 U1540 ( .Y(n4464), .A(n4463) );
  inv02 U1541 ( .Y(n7693), .A(n7691) );
  nand02 U1542 ( .Y(n7995), .A0(n4465), .A1(n4466) );
  inv01 U1543 ( .Y(n4467), .A(n7422) );
  inv01 U1544 ( .Y(n4468), .A(fract_28_i[23]) );
  inv01 U1545 ( .Y(n4469), .A(n7689) );
  inv01 U1546 ( .Y(n4470), .A(fract_28_i[24]) );
  nand02 U1547 ( .Y(n4471), .A0(n4467), .A1(n4468) );
  nand02 U1548 ( .Y(n4472), .A0(n4467), .A1(n4469) );
  nand02 U1549 ( .Y(n4473), .A0(n4468), .A1(n4470) );
  nand02 U1550 ( .Y(n4474), .A0(n4469), .A1(n4470) );
  nand02 U1551 ( .Y(n4475), .A0(n4471), .A1(n4472) );
  inv01 U1552 ( .Y(n4465), .A(n4475) );
  nand02 U1553 ( .Y(n4476), .A0(n4473), .A1(n4474) );
  inv01 U1554 ( .Y(n4466), .A(n4476) );
  ao22 U1555 ( .Y(n4477), .A0(n7693), .A1(fract_28_i[23]), .B0(n7695), .B1(
        fract_28_i[26]) );
  inv01 U1556 ( .Y(n4478), .A(n4477) );
  buf04 U1557 ( .Y(n7674), .A(n7893) );
  inv08 U1558 ( .Y(n5873), .A(n7674) );
  nand02 U1559 ( .Y(n8015), .A0(n4479), .A1(n4480) );
  inv01 U1560 ( .Y(n4481), .A(n2550_8_) );
  inv01 U1561 ( .Y(n4482), .A(s_expo9_1[8]) );
  inv01 U1562 ( .Y(n4483), .A(n7667) );
  nand02 U1563 ( .Y(n4479), .A0(n7667), .A1(n4481) );
  nand02 U1564 ( .Y(n4480), .A0(n4482), .A1(n4483) );
  buf04 U1565 ( .Y(n7667), .A(n8016) );
  ao22 U1566 ( .Y(n4484), .A0(n7676), .A1(n7934), .B0(n7674), .B1(n7931) );
  inv01 U1567 ( .Y(n4485), .A(n4484) );
  ao22 U1568 ( .Y(n4486), .A0(n7676), .A1(n7931), .B0(n7675), .B1(n7834) );
  inv01 U1569 ( .Y(n4487), .A(n4486) );
  or02 U1570 ( .Y(n4488), .A0(n8090), .A1(n8091) );
  inv01 U1571 ( .Y(n4489), .A(n4488) );
  buf02 U1572 ( .Y(n4490), .A(s_fracto28_12090_6_) );
  buf02 U1573 ( .Y(n4491), .A(s_fracto28_12090_22_) );
  buf02 U1574 ( .Y(n4492), .A(s_fracto28_12090_14_) );
  ao22 U1575 ( .Y(n4493), .A0(n7615), .A1(n7842), .B0(n7678), .B1(n7899) );
  inv01 U1576 ( .Y(n4494), .A(n4493) );
  buf02 U1577 ( .Y(n4495), .A(s_fracto28_12090_21_) );
  ao22 U1578 ( .Y(n4496), .A0(n7623), .A1(n7835), .B0(n7675), .B1(n7868) );
  inv01 U1579 ( .Y(n4497), .A(n4496) );
  nand02 U1580 ( .Y(n7836), .A0(n4498), .A1(n4499) );
  inv01 U1581 ( .Y(n4500), .A(n7849) );
  inv01 U1582 ( .Y(n4501), .A(n7848) );
  inv01 U1583 ( .Y(n4502), .A(n7676) );
  inv01 U1584 ( .Y(n4503), .A(n7677) );
  nand02 U1585 ( .Y(n4504), .A0(n4500), .A1(n4501) );
  nand02 U1586 ( .Y(n4505), .A0(n4500), .A1(n4502) );
  nand02 U1587 ( .Y(n4506), .A0(n4501), .A1(n4503) );
  nand02 U1588 ( .Y(n4507), .A0(n4502), .A1(n4503) );
  nand02 U1589 ( .Y(n4508), .A0(n4504), .A1(n4505) );
  inv01 U1590 ( .Y(n4498), .A(n4508) );
  nand02 U1591 ( .Y(n4509), .A0(n4506), .A1(n4507) );
  inv01 U1592 ( .Y(n4499), .A(n4509) );
  ao22 U1593 ( .Y(n4510), .A0(n7674), .A1(n7848), .B0(n7669), .B1(n7842) );
  inv01 U1594 ( .Y(n4511), .A(n4510) );
  nand02 U1595 ( .Y(n4512), .A0(n8102), .A1(n7887) );
  inv02 U1596 ( .Y(n4513), .A(n4512) );
  inv01 U1597 ( .Y(n7797), .A(n4514) );
  inv01 U1598 ( .Y(n4515), .A(opb_i[23]) );
  inv01 U1599 ( .Y(n4516), .A(opb_i[24]) );
  inv01 U1600 ( .Y(n4517), .A(opb_i[25]) );
  inv01 U1601 ( .Y(n4518), .A(opb_i[26]) );
  nor02 U1602 ( .Y(n4514), .A0(n4519), .A1(n4520) );
  nor02 U1603 ( .Y(n4521), .A0(n4515), .A1(n4516) );
  inv01 U1604 ( .Y(n4519), .A(n4521) );
  nor02 U1605 ( .Y(n4522), .A0(n4517), .A1(n4518) );
  inv01 U1606 ( .Y(n4520), .A(n4522) );
  or02 U1607 ( .Y(n4523), .A0(opa_i[10]), .A1(opa_i[0]) );
  inv01 U1608 ( .Y(n4524), .A(n4523) );
  inv01 U1609 ( .Y(s_fracto28_12090_13_), .A(n4525) );
  inv01 U1610 ( .Y(n4526), .A(n7985) );
  inv01 U1611 ( .Y(n4527), .A(n7984) );
  inv01 U1612 ( .Y(n4528), .A(n4605) );
  inv01 U1613 ( .Y(n4529), .A(n4267) );
  nor02 U1614 ( .Y(n4525), .A0(n4530), .A1(n4531) );
  nor02 U1615 ( .Y(n4532), .A0(n4526), .A1(n4527) );
  inv01 U1616 ( .Y(n4530), .A(n4532) );
  nor02 U1617 ( .Y(n4533), .A0(n4528), .A1(n4529) );
  inv01 U1618 ( .Y(n4531), .A(n4533) );
  inv01 U1619 ( .Y(s_fracto28_12090_5_), .A(n4534) );
  inv01 U1620 ( .Y(n4535), .A(n7859) );
  inv01 U1621 ( .Y(n4536), .A(n4622) );
  inv01 U1622 ( .Y(n4537), .A(n4614) );
  inv01 U1623 ( .Y(n4538), .A(n4269) );
  nor02 U1624 ( .Y(n4534), .A0(n4539), .A1(n4540) );
  nor02 U1625 ( .Y(n4541), .A0(n4535), .A1(n4536) );
  inv01 U1626 ( .Y(n4539), .A(n4541) );
  nor02 U1627 ( .Y(n4542), .A0(n4537), .A1(n4538) );
  inv01 U1628 ( .Y(n4540), .A(n4542) );
  nand02 U1629 ( .Y(n7724), .A0(n4543), .A1(n4544) );
  inv01 U1630 ( .Y(n4545), .A(n7731) );
  inv01 U1631 ( .Y(n4546), .A(n7730) );
  inv01 U1632 ( .Y(n4547), .A(opa_i[31]) );
  inv01 U1633 ( .Y(n4548), .A(opb_i[31]) );
  nand02 U1634 ( .Y(n4549), .A0(n4545), .A1(n4546) );
  nand02 U1635 ( .Y(n4550), .A0(n4545), .A1(n4547) );
  nand02 U1636 ( .Y(n4551), .A0(n4546), .A1(n4548) );
  nand02 U1637 ( .Y(n4552), .A0(n4547), .A1(n4548) );
  nand02 U1638 ( .Y(n4553), .A0(n4549), .A1(n4550) );
  inv01 U1639 ( .Y(n4543), .A(n4553) );
  nand02 U1640 ( .Y(n4554), .A0(n4551), .A1(n4552) );
  inv01 U1641 ( .Y(n4544), .A(n4554) );
  nand02 U1642 ( .Y(n7982), .A0(n4555), .A1(n4556) );
  inv01 U1643 ( .Y(n4557), .A(n7603) );
  inv01 U1644 ( .Y(n4558), .A(n7852) );
  inv01 U1645 ( .Y(n4559), .A(n7670) );
  inv01 U1646 ( .Y(n4560), .A(n7673) );
  nand02 U1647 ( .Y(n4561), .A0(n4557), .A1(n4558) );
  nand02 U1648 ( .Y(n4562), .A0(n4557), .A1(n4559) );
  nand02 U1649 ( .Y(n4563), .A0(n4558), .A1(n4560) );
  nand02 U1650 ( .Y(n4564), .A0(n4559), .A1(n4560) );
  nand02 U1651 ( .Y(n4565), .A0(n4561), .A1(n4562) );
  inv01 U1652 ( .Y(n4555), .A(n4565) );
  nand02 U1653 ( .Y(n4566), .A0(n4563), .A1(n4564) );
  inv01 U1654 ( .Y(n4556), .A(n4566) );
  ao22 U1655 ( .Y(n4567), .A0(n7675), .A1(n7852), .B0(n7677), .B1(n7602) );
  inv01 U1656 ( .Y(n4568), .A(n4567) );
  or03 U1657 ( .Y(n4569), .A0(n8076), .A1(n4610), .A2(n7316) );
  inv01 U1658 ( .Y(n4570), .A(n4569) );
  nor02 U1659 ( .Y(n7710), .A0(exp_i[1]), .A1(n4571) );
  nor02 U1660 ( .Y(n4572), .A0(exp_i[0]), .A1(exp_i[2]) );
  inv01 U1661 ( .Y(n4571), .A(n4572) );
  ao22 U1662 ( .Y(n4573), .A0(n7678), .A1(n7857), .B0(n7671), .B1(n7858) );
  inv01 U1663 ( .Y(n4574), .A(n4573) );
  ao22 U1664 ( .Y(n4575), .A0(n7677), .A1(n7819), .B0(n7675), .B1(n7825) );
  inv01 U1665 ( .Y(n4576), .A(n4575) );
  inv01 U1666 ( .Y(n7789), .A(n4577) );
  inv01 U1667 ( .Y(n4578), .A(n7795) );
  inv01 U1668 ( .Y(n4579), .A(n7794) );
  inv01 U1669 ( .Y(n4580), .A(n7793) );
  nand02 U1670 ( .Y(n4577), .A0(n4580), .A1(n4581) );
  nand02 U1671 ( .Y(n4582), .A0(n4578), .A1(n4579) );
  inv01 U1672 ( .Y(n4581), .A(n4582) );
  inv02 U1673 ( .Y(n4871), .A(n7940) );
  ao22 U1674 ( .Y(n4583), .A0(n7677), .A1(n7855), .B0(n7670), .B1(n7856) );
  inv01 U1675 ( .Y(n4584), .A(n4583) );
  inv01 U1676 ( .Y(n7796), .A(n4585) );
  inv01 U1677 ( .Y(n4586), .A(n7792) );
  inv01 U1678 ( .Y(n4587), .A(n7801) );
  inv01 U1679 ( .Y(n4588), .A(n4265) );
  nand02 U1680 ( .Y(n4585), .A0(n4588), .A1(n4589) );
  nand02 U1681 ( .Y(n4590), .A0(n4586), .A1(n4587) );
  inv01 U1682 ( .Y(n4589), .A(n4590) );
  inv02 U1683 ( .Y(n4675), .A(n7850) );
  ao22 U1684 ( .Y(n4591), .A0(n7675), .A1(n7856), .B0(n7677), .B1(n7858) );
  inv01 U1685 ( .Y(n4592), .A(n4591) );
  nand02 U1686 ( .Y(n7945), .A0(n4593), .A1(n4594) );
  inv01 U1687 ( .Y(n4595), .A(n7924) );
  inv01 U1688 ( .Y(n4596), .A(n7920) );
  inv01 U1689 ( .Y(n4597), .A(n7669) );
  nand02 U1690 ( .Y(n4598), .A0(n4595), .A1(n4596) );
  nand02 U1691 ( .Y(n4599), .A0(n4595), .A1(n5873) );
  nand02 U1692 ( .Y(n4600), .A0(n4596), .A1(n4597) );
  nand02 U1693 ( .Y(n4601), .A0(n5873), .A1(n4597) );
  nand02 U1694 ( .Y(n4602), .A0(n4598), .A1(n4599) );
  inv01 U1695 ( .Y(n4593), .A(n4602) );
  nand02 U1696 ( .Y(n4603), .A0(n4600), .A1(n4601) );
  inv01 U1697 ( .Y(n4594), .A(n4603) );
  ao22 U1698 ( .Y(n4604), .A0(n7676), .A1(n7920), .B0(n7677), .B1(n7827) );
  inv01 U1699 ( .Y(n4605), .A(n4604) );
  ao22 U1700 ( .Y(n4606), .A0(n7669), .A1(n7913), .B0(n7674), .B1(n7944) );
  inv01 U1701 ( .Y(n4607), .A(n4606) );
  buf02 U1702 ( .Y(n4608), .A(n7977) );
  nand03 U1703 ( .Y(n4609), .A0(n8104), .A1(n7879), .A2(fract_28_i[4]) );
  inv02 U1704 ( .Y(n4610), .A(n4609) );
  ao22 U1705 ( .Y(n4611), .A0(n7669), .A1(n7857), .B0(n7676), .B1(n7944) );
  inv01 U1706 ( .Y(n4612), .A(n4611) );
  ao22 U1707 ( .Y(n4613), .A0(n7676), .A1(n7861), .B0(n7678), .B1(n7862) );
  inv01 U1708 ( .Y(n4614), .A(n4613) );
  ao22 U1709 ( .Y(n4615), .A0(n7678), .A1(n7910), .B0(n7676), .B1(n7908) );
  inv01 U1710 ( .Y(n4616), .A(n4615) );
  ao22 U1711 ( .Y(n4617), .A0(n7678), .A1(n7916), .B0(n7676), .B1(n7923) );
  inv01 U1712 ( .Y(n4618), .A(n4617) );
  nand03 U1713 ( .Y(n4619), .A0(n4732), .A1(n7986), .A2(fract_28_i[0]) );
  inv02 U1714 ( .Y(n4620), .A(n4619) );
  ao22 U1715 ( .Y(n4621), .A0(n7675), .A1(n7860), .B0(n7677), .B1(n7818) );
  inv01 U1716 ( .Y(n4622), .A(n4621) );
  ao22 U1717 ( .Y(n4623), .A0(n7675), .A1(n7853), .B0(n7676), .B1(n7854) );
  inv01 U1718 ( .Y(n4624), .A(n4623) );
  inv01 U1719 ( .Y(n7798), .A(n4625) );
  inv01 U1720 ( .Y(n4626), .A(opb_i[27]) );
  inv01 U1721 ( .Y(n4627), .A(opb_i[28]) );
  inv01 U1722 ( .Y(n4628), .A(opb_i[29]) );
  inv01 U1723 ( .Y(n4629), .A(opb_i[30]) );
  nor02 U1724 ( .Y(n4625), .A0(n4630), .A1(n4631) );
  nor02 U1725 ( .Y(n4632), .A0(n4626), .A1(n4627) );
  inv01 U1726 ( .Y(n4630), .A(n4632) );
  nor02 U1727 ( .Y(n4633), .A0(n4628), .A1(n4629) );
  inv01 U1728 ( .Y(n4631), .A(n4633) );
  nand02 U1729 ( .Y(n7984), .A0(n4634), .A1(n4635) );
  inv01 U1730 ( .Y(n4636), .A(n7825) );
  inv01 U1731 ( .Y(n4637), .A(n7819) );
  inv01 U1732 ( .Y(n4638), .A(n7673) );
  inv01 U1733 ( .Y(n4639), .A(n7670) );
  nand02 U1734 ( .Y(n4640), .A0(n4636), .A1(n4637) );
  nand02 U1735 ( .Y(n4641), .A0(n4636), .A1(n4638) );
  nand02 U1736 ( .Y(n4642), .A0(n4637), .A1(n4639) );
  nand02 U1737 ( .Y(n4643), .A0(n4638), .A1(n4639) );
  nand02 U1738 ( .Y(n4644), .A0(n4640), .A1(n4641) );
  inv01 U1739 ( .Y(n4634), .A(n4644) );
  nand02 U1740 ( .Y(n4645), .A0(n4642), .A1(n4643) );
  inv01 U1741 ( .Y(n4635), .A(n4645) );
  ao22 U1742 ( .Y(n4646), .A0(n7678), .A1(n7913), .B0(n7674), .B1(n7854) );
  inv01 U1743 ( .Y(n4647), .A(n4646) );
  or02 U1744 ( .Y(n4648), .A0(n8047), .A1(n8048) );
  inv01 U1745 ( .Y(n4649), .A(n4648) );
  xor2 U1746 ( .Y(n4650), .A0(opa_i[31]), .A1(n4806) );
  inv01 U1747 ( .Y(n4651), .A(n4650) );
  inv01 U1748 ( .Y(n7809), .A(n4652) );
  inv01 U1749 ( .Y(n4653), .A(n7813) );
  inv01 U1750 ( .Y(n4654), .A(rmode_i[0]) );
  inv01 U1751 ( .Y(n4655), .A(n7811) );
  nand02 U1752 ( .Y(n4652), .A0(n4655), .A1(n4656) );
  nand02 U1753 ( .Y(n4657), .A0(n4653), .A1(n4654) );
  inv01 U1754 ( .Y(n4656), .A(n4657) );
  ao22 U1755 ( .Y(n4658), .A0(n7850), .A1(n7601), .B0(n7623), .B1(n7852) );
  inv01 U1756 ( .Y(n4659), .A(n4658) );
  nand02 U1757 ( .Y(n7985), .A0(n4660), .A1(n4661) );
  inv01 U1758 ( .Y(n4662), .A(n7862) );
  inv01 U1759 ( .Y(n4663), .A(n7861) );
  inv01 U1760 ( .Y(n4664), .A(n7669) );
  nand02 U1761 ( .Y(n4665), .A0(n4662), .A1(n4663) );
  nand02 U1762 ( .Y(n4666), .A0(n4662), .A1(n5873) );
  nand02 U1763 ( .Y(n4667), .A0(n4663), .A1(n4664) );
  nand02 U1764 ( .Y(n4668), .A0(n5873), .A1(n4664) );
  nand02 U1765 ( .Y(n4669), .A0(n4665), .A1(n4666) );
  inv01 U1766 ( .Y(n4660), .A(n4669) );
  nand02 U1767 ( .Y(n4670), .A0(n4667), .A1(n4668) );
  inv01 U1768 ( .Y(n4661), .A(n4670) );
  nand02 U1769 ( .Y(n7859), .A0(n4671), .A1(n4672) );
  inv02 U1770 ( .Y(n4673), .A(n7825) );
  inv01 U1771 ( .Y(n4674), .A(n7819) );
  inv01 U1772 ( .Y(n4676), .A(n7623) );
  nand02 U1773 ( .Y(n4677), .A0(n4673), .A1(n4674) );
  nand02 U1774 ( .Y(n4678), .A0(n4673), .A1(n4675) );
  nand02 U1775 ( .Y(n4679), .A0(n4674), .A1(n4676) );
  nand02 U1776 ( .Y(n4680), .A0(n4675), .A1(n4676) );
  nand02 U1777 ( .Y(n4681), .A0(n4677), .A1(n4678) );
  inv01 U1778 ( .Y(n4671), .A(n4681) );
  nand02 U1779 ( .Y(n4682), .A0(n4679), .A1(n4680) );
  inv01 U1780 ( .Y(n4672), .A(n4682) );
  nand02 U1781 ( .Y(n7942), .A0(n4683), .A1(n4684) );
  inv02 U1782 ( .Y(n4685), .A(n7857) );
  inv01 U1783 ( .Y(n4686), .A(n7854) );
  inv01 U1784 ( .Y(n4687), .A(n7615) );
  nand02 U1785 ( .Y(n4688), .A0(n4685), .A1(n4686) );
  nand02 U1786 ( .Y(n4689), .A0(n4685), .A1(n4871) );
  nand02 U1787 ( .Y(n4690), .A0(n4686), .A1(n4687) );
  nand02 U1788 ( .Y(n4691), .A0(n4871), .A1(n4687) );
  nand02 U1789 ( .Y(n4692), .A0(n4688), .A1(n4689) );
  inv01 U1790 ( .Y(n4683), .A(n4692) );
  nand02 U1791 ( .Y(n4693), .A0(n4690), .A1(n4691) );
  inv01 U1792 ( .Y(n4684), .A(n4693) );
  nand02 U1793 ( .Y(n7946), .A0(n4694), .A1(n4695) );
  inv01 U1794 ( .Y(n4696), .A(n7862) );
  inv01 U1795 ( .Y(n4697), .A(n7861) );
  inv01 U1796 ( .Y(n4698), .A(n7615) );
  nand02 U1797 ( .Y(n4699), .A0(n4696), .A1(n4697) );
  nand02 U1798 ( .Y(n4700), .A0(n4696), .A1(n4871) );
  nand02 U1799 ( .Y(n4701), .A0(n4697), .A1(n4698) );
  nand02 U1800 ( .Y(n4702), .A0(n4871), .A1(n4698) );
  nand02 U1801 ( .Y(n4703), .A0(n4699), .A1(n4700) );
  inv01 U1802 ( .Y(n4694), .A(n4703) );
  nand02 U1803 ( .Y(n4704), .A0(n4701), .A1(n4702) );
  inv01 U1804 ( .Y(n4695), .A(n4704) );
  nor02 U1805 ( .Y(n7711), .A0(exp_i[4]), .A1(n4705) );
  nor02 U1806 ( .Y(n4706), .A0(exp_i[3]), .A1(exp_i[5]) );
  inv01 U1807 ( .Y(n4705), .A(n4706) );
  inv02 U1808 ( .Y(n4707), .A(n7706) );
  inv04 U1809 ( .Y(n5608), .A(n7938) );
  inv02 U1810 ( .Y(n7938), .A(n7501) );
  buf02 U1811 ( .Y(n4708), .A(n7729) );
  or03 U1812 ( .Y(n4709), .A0(n7739), .A1(n7734), .A2(s_expo9_2[8]) );
  inv01 U1813 ( .Y(n4710), .A(n4709) );
  xor2 U1814 ( .Y(n4711), .A0(n8043), .A1(exp_i[5]) );
  inv01 U1815 ( .Y(n4712), .A(n4711) );
  or03 U1816 ( .Y(n4713), .A0(n7750), .A1(n2866_8_), .A2(n7570) );
  inv01 U1817 ( .Y(n4714), .A(n4713) );
  xor2 U1818 ( .Y(n4715), .A0(n7191), .A1(n7708) );
  inv01 U1819 ( .Y(n4716), .A(n4715) );
  inv01 U1820 ( .Y(n8028), .A(n4717) );
  nor02 U1821 ( .Y(n4718), .A0(n7542), .A1(n8038) );
  inv01 U1822 ( .Y(n4719), .A(n8046) );
  nor02 U1823 ( .Y(n4717), .A0(n4718), .A1(n4719) );
  buf02 U1824 ( .Y(n4720), .A(n8037) );
  inv01 U1825 ( .Y(n7800), .A(n4721) );
  inv01 U1826 ( .Y(n4722), .A(opa_i[27]) );
  inv01 U1827 ( .Y(n4723), .A(opa_i[28]) );
  inv01 U1828 ( .Y(n4724), .A(opa_i[29]) );
  inv01 U1829 ( .Y(n4725), .A(opa_i[30]) );
  nor02 U1830 ( .Y(n4721), .A0(n4726), .A1(n4727) );
  nor02 U1831 ( .Y(n4728), .A0(n4722), .A1(n4723) );
  inv01 U1832 ( .Y(n4726), .A(n4728) );
  nor02 U1833 ( .Y(n4729), .A0(n4724), .A1(n4725) );
  inv01 U1834 ( .Y(n4727), .A(n4729) );
  inv01 U1835 ( .Y(n4730), .A(n6554) );
  nand03 U1836 ( .Y(n4731), .A0(n7955), .A1(n7889), .A2(n6966) );
  inv02 U1837 ( .Y(n4732), .A(n4731) );
  nand02 U1838 ( .Y(n8027), .A0(n4733), .A1(n4734) );
  inv01 U1839 ( .Y(n4735), .A(n7793) );
  inv01 U1840 ( .Y(n4736), .A(n7707) );
  inv01 U1841 ( .Y(n4737), .A(n8028) );
  inv01 U1842 ( .Y(n4738), .A(n8029) );
  nand02 U1843 ( .Y(n4739), .A0(n4735), .A1(n4736) );
  nand02 U1844 ( .Y(n4740), .A0(n4735), .A1(n4737) );
  nand02 U1845 ( .Y(n4741), .A0(n4736), .A1(n4738) );
  nand02 U1846 ( .Y(n4742), .A0(n4737), .A1(n4738) );
  nand02 U1847 ( .Y(n4743), .A0(n4739), .A1(n4740) );
  inv01 U1848 ( .Y(n4733), .A(n4743) );
  nand02 U1849 ( .Y(n4744), .A0(n4741), .A1(n4742) );
  inv01 U1850 ( .Y(n4734), .A(n4744) );
  nand03 U1851 ( .Y(n4745), .A0(n7245), .A1(n7947), .A2(n8072) );
  inv02 U1852 ( .Y(n4746), .A(n4745) );
  xor2 U1853 ( .Y(n4747), .A0(n7188), .A1(n7190) );
  inv01 U1854 ( .Y(n4748), .A(n4747) );
  xor2 U1855 ( .Y(n4749), .A0(n7704), .A1(exp_i[0]) );
  inv01 U1856 ( .Y(n4750), .A(n4749) );
  inv01 U1857 ( .Y(n8095), .A(n4751) );
  inv01 U1858 ( .Y(n4752), .A(n8075) );
  inv01 U1859 ( .Y(n4753), .A(n8079) );
  inv01 U1860 ( .Y(n4754), .A(n8078) );
  nand02 U1861 ( .Y(n4751), .A0(n4754), .A1(n4755) );
  nand02 U1862 ( .Y(n4756), .A0(n4752), .A1(n4753) );
  inv01 U1863 ( .Y(n4755), .A(n4756) );
  or03 U1864 ( .Y(n4757), .A0(n8081), .A1(n8082), .A2(n8077) );
  inv01 U1865 ( .Y(n4758), .A(n4757) );
  inv01 U1866 ( .Y(n7799), .A(n4759) );
  inv01 U1867 ( .Y(n4760), .A(opa_i[23]) );
  inv01 U1868 ( .Y(n4761), .A(opa_i[24]) );
  inv01 U1869 ( .Y(n4762), .A(opa_i[25]) );
  inv01 U1870 ( .Y(n4763), .A(opa_i[26]) );
  nor02 U1871 ( .Y(n4759), .A0(n4764), .A1(n4765) );
  nor02 U1872 ( .Y(n4766), .A0(n4760), .A1(n4761) );
  inv01 U1873 ( .Y(n4764), .A(n4766) );
  nor02 U1874 ( .Y(n4767), .A0(n4762), .A1(n4763) );
  inv01 U1875 ( .Y(n4765), .A(n4767) );
  or03 U1876 ( .Y(n4768), .A0(n8066), .A1(n8064), .A2(n8065) );
  inv01 U1877 ( .Y(n4769), .A(n4768) );
  xor2 U1878 ( .Y(n4770), .A0(n8038), .A1(n8039) );
  inv01 U1879 ( .Y(n4771), .A(n4770) );
  inv01 U1880 ( .Y(n8111), .A(n4772) );
  inv01 U1881 ( .Y(n4773), .A(n8060) );
  inv01 U1882 ( .Y(n4774), .A(n8058) );
  inv01 U1883 ( .Y(n4775), .A(n8080) );
  nand02 U1884 ( .Y(n4772), .A0(n4775), .A1(n4776) );
  nand02 U1885 ( .Y(n4777), .A0(n4773), .A1(n4774) );
  inv01 U1886 ( .Y(n4776), .A(n4777) );
  inv01 U1887 ( .Y(n4778), .A(n8017) );
  ao21 U1888 ( .Y(n4779), .A0(n8040), .A1(exp_i[6]), .B0(exp_i[7]) );
  inv01 U1889 ( .Y(n4780), .A(n4779) );
  inv01 U1890 ( .Y(n7886), .A(n4781) );
  nor02 U1891 ( .Y(n4782), .A0(n7879), .A1(n7700) );
  nor02 U1892 ( .Y(n4783), .A0(n7889), .A1(n7881) );
  nor02 U1893 ( .Y(n4784), .A0(n7880), .A1(n7701) );
  nor02 U1894 ( .Y(n4781), .A0(n4784), .A1(n4785) );
  nor02 U1895 ( .Y(n4786), .A0(n4782), .A1(n4783) );
  inv01 U1896 ( .Y(n4785), .A(n4786) );
  inv01 U1897 ( .Y(n7872), .A(n4787) );
  nor02 U1898 ( .Y(n4788), .A0(n7882), .A1(n7698) );
  nor02 U1899 ( .Y(n4789), .A0(n7880), .A1(n7881) );
  nor02 U1900 ( .Y(n4790), .A0(n7879), .A1(n7701) );
  nor02 U1901 ( .Y(n4787), .A0(n4790), .A1(n4791) );
  nor02 U1902 ( .Y(n4792), .A0(n4788), .A1(n4789) );
  inv01 U1903 ( .Y(n4791), .A(n4792) );
  inv02 U1904 ( .Y(n7889), .A(fract_28_i[3]) );
  buf02 U1905 ( .Y(n7700), .A(n7697) );
  inv02 U1906 ( .Y(n7879), .A(fract_28_i[5]) );
  inv01 U1907 ( .Y(n7953), .A(n4793) );
  nor02 U1908 ( .Y(n4794), .A0(n7880), .A1(n7699) );
  nor02 U1909 ( .Y(n4795), .A0(n7955), .A1(n7881) );
  nor02 U1910 ( .Y(n4796), .A0(n7889), .A1(n7701) );
  nor02 U1911 ( .Y(n4793), .A0(n4796), .A1(n4797) );
  nor02 U1912 ( .Y(n4798), .A0(n4794), .A1(n4795) );
  inv01 U1913 ( .Y(n4797), .A(n4798) );
  inv02 U1914 ( .Y(n7880), .A(fract_28_i[4]) );
  buf02 U1915 ( .Y(n7699), .A(n7696) );
  inv01 U1916 ( .Y(n8006), .A(n4799) );
  nor02 U1917 ( .Y(n4800), .A0(n7889), .A1(n7698) );
  nor02 U1918 ( .Y(n4801), .A0(n7986), .A1(n7881) );
  nor02 U1919 ( .Y(n4802), .A0(n7955), .A1(n7701) );
  nor02 U1920 ( .Y(n4799), .A0(n4802), .A1(n4803) );
  nor02 U1921 ( .Y(n4804), .A0(n4800), .A1(n4801) );
  inv01 U1922 ( .Y(n4803), .A(n4804) );
  xor2 U1923 ( .Y(n4805), .A0(opb_i[31]), .A1(fpu_op_i) );
  inv01 U1924 ( .Y(n4806), .A(n4805) );
  nand02 U1925 ( .Y(n7989), .A0(n4807), .A1(n4808) );
  inv01 U1926 ( .Y(n4809), .A(n7935) );
  inv01 U1927 ( .Y(n4810), .A(n7658) );
  inv01 U1928 ( .Y(n4811), .A(n7865) );
  inv01 U1929 ( .Y(n4812), .A(s_shl1_3_) );
  inv02 U1930 ( .Y(n4813), .A(n7678) );
  nand02 U1931 ( .Y(n4814), .A0(n4809), .A1(n4810) );
  nand02 U1932 ( .Y(n4815), .A0(n4809), .A1(n4811) );
  nand02 U1933 ( .Y(n4816), .A0(n4809), .A1(n4812) );
  nand02 U1934 ( .Y(n4817), .A0(n4810), .A1(n4813) );
  nand02 U1935 ( .Y(n4818), .A0(n4811), .A1(n4813) );
  nand02 U1936 ( .Y(n4819), .A0(n4812), .A1(n4813) );
  nand02 U1937 ( .Y(n4820), .A0(n4814), .A1(n4815) );
  inv01 U1938 ( .Y(n4821), .A(n4820) );
  nand02 U1939 ( .Y(n4822), .A0(n4816), .A1(n4821) );
  inv01 U1940 ( .Y(n4807), .A(n4822) );
  nand02 U1941 ( .Y(n4823), .A0(n4817), .A1(n4818) );
  inv01 U1942 ( .Y(n4824), .A(n4823) );
  nand02 U1943 ( .Y(n4825), .A0(n4819), .A1(n4824) );
  inv01 U1944 ( .Y(n4808), .A(n4825) );
  nand02 U1945 ( .Y(n7837), .A0(n4826), .A1(n4827) );
  inv01 U1946 ( .Y(n4828), .A(n7846) );
  inv01 U1947 ( .Y(n4829), .A(n7625) );
  inv01 U1948 ( .Y(n4830), .A(n7844) );
  inv01 U1949 ( .Y(n4831), .A(n7843) );
  inv02 U1950 ( .Y(n4832), .A(n7675) );
  nand02 U1951 ( .Y(n4833), .A0(n4828), .A1(n4829) );
  nand02 U1952 ( .Y(n4834), .A0(n4828), .A1(n4830) );
  nand02 U1953 ( .Y(n4835), .A0(n4828), .A1(n4831) );
  nand02 U1954 ( .Y(n4836), .A0(n4829), .A1(n4832) );
  nand02 U1955 ( .Y(n4837), .A0(n4830), .A1(n4832) );
  nand02 U1956 ( .Y(n4838), .A0(n4831), .A1(n4832) );
  nand02 U1957 ( .Y(n4839), .A0(n4833), .A1(n4834) );
  inv01 U1958 ( .Y(n4840), .A(n4839) );
  nand02 U1959 ( .Y(n4841), .A0(n4835), .A1(n4840) );
  inv01 U1960 ( .Y(n4826), .A(n4841) );
  nand02 U1961 ( .Y(n4842), .A0(n4836), .A1(n4837) );
  inv01 U1962 ( .Y(n4843), .A(n4842) );
  nand02 U1963 ( .Y(n4844), .A0(n4838), .A1(n4843) );
  inv01 U1964 ( .Y(n4827), .A(n4844) );
  inv01 U1965 ( .Y(n7865), .A(n7991) );
  inv01 U1966 ( .Y(n7843), .A(n7981) );
  nand02 U1967 ( .Y(n7863), .A0(n4845), .A1(n4846) );
  inv01 U1968 ( .Y(n4847), .A(n7831) );
  inv01 U1969 ( .Y(n4848), .A(n7660) );
  inv01 U1970 ( .Y(n4849), .A(n7866) );
  inv01 U1971 ( .Y(n4850), .A(n7865) );
  nand02 U1972 ( .Y(n4851), .A0(n4847), .A1(n4848) );
  nand02 U1973 ( .Y(n4852), .A0(n4847), .A1(n4849) );
  nand02 U1974 ( .Y(n4853), .A0(n4847), .A1(n4850) );
  nand02 U1975 ( .Y(n4854), .A0(n4848), .A1(n4675) );
  nand02 U1976 ( .Y(n4855), .A0(n4849), .A1(n4675) );
  nand02 U1977 ( .Y(n4856), .A0(n4850), .A1(n4675) );
  nand02 U1978 ( .Y(n4857), .A0(n4851), .A1(n4852) );
  inv01 U1979 ( .Y(n4858), .A(n4857) );
  nand02 U1980 ( .Y(n4859), .A0(n4853), .A1(n4858) );
  inv01 U1981 ( .Y(n4845), .A(n4859) );
  nand02 U1982 ( .Y(n4860), .A0(n4854), .A1(n4855) );
  inv01 U1983 ( .Y(n4861), .A(n4860) );
  nand02 U1984 ( .Y(n4862), .A0(n4856), .A1(n4861) );
  inv01 U1985 ( .Y(n4846), .A(n4862) );
  ao32 U1986 ( .Y(n4863), .A0(n7865), .A1(n7866), .A2(n7647), .B0(n7678), .B1(
        n7927) );
  inv01 U1987 ( .Y(n4864), .A(n4863) );
  nand02 U1988 ( .Y(n7936), .A0(n4865), .A1(n4866) );
  inv01 U1989 ( .Y(n4867), .A(n7848) );
  inv01 U1990 ( .Y(n4868), .A(n7654) );
  inv01 U1991 ( .Y(n4869), .A(n7844) );
  inv01 U1992 ( .Y(n4870), .A(n7843) );
  nand02 U1993 ( .Y(n4872), .A0(n4867), .A1(n4868) );
  nand02 U1994 ( .Y(n4873), .A0(n4867), .A1(n4869) );
  nand02 U1995 ( .Y(n4874), .A0(n4867), .A1(n4870) );
  nand02 U1996 ( .Y(n4875), .A0(n4868), .A1(n4871) );
  nand02 U1997 ( .Y(n4876), .A0(n4869), .A1(n4871) );
  nand02 U1998 ( .Y(n4877), .A0(n4870), .A1(n4871) );
  nand02 U1999 ( .Y(n4878), .A0(n4872), .A1(n4873) );
  inv01 U2000 ( .Y(n4879), .A(n4878) );
  nand02 U2001 ( .Y(n4880), .A0(n4874), .A1(n4879) );
  inv01 U2002 ( .Y(n4865), .A(n4880) );
  nand02 U2003 ( .Y(n4881), .A0(n4875), .A1(n4876) );
  inv01 U2004 ( .Y(n4882), .A(n4881) );
  nand02 U2005 ( .Y(n4883), .A0(n4877), .A1(n4882) );
  inv01 U2006 ( .Y(n4866), .A(n4883) );
  inv02 U2007 ( .Y(n7831), .A(n7616) );
  ao32 U2008 ( .Y(n4884), .A0(n7843), .A1(n7654), .A2(s_shr1_3_), .B0(n7678), 
        .B1(n7892) );
  inv01 U2009 ( .Y(n4885), .A(n4884) );
  inv01 U2010 ( .Y(s_ine_o), .A(n4886) );
  inv01 U2011 ( .Y(n4887), .A(n7427) );
  inv01 U2012 ( .Y(n4888), .A(n7413) );
  inv01 U2013 ( .Y(n4889), .A(n7796) );
  nand02 U2014 ( .Y(n4886), .A0(n4889), .A1(n4890) );
  nand02 U2015 ( .Y(n4891), .A0(n4887), .A1(n4888) );
  inv01 U2016 ( .Y(n4890), .A(n4891) );
  nand02 U2017 ( .Y(n4892), .A0(n8106), .A1(n7974) );
  inv04 U2018 ( .Y(n4893), .A(n4892) );
  nand02 U2019 ( .Y(n4894), .A0(n8113), .A1(n7956) );
  inv02 U2020 ( .Y(n4895), .A(n4894) );
  inv02 U2021 ( .Y(s_expo9_2[8]), .A(n8015) );
  inv01 U2022 ( .Y(s_output_o[26]), .A(n4896) );
  nor02 U2023 ( .Y(n4897), .A0(n7745), .A1(n7651) );
  nor02 U2024 ( .Y(n4898), .A0(n7744), .A1(n7650) );
  inv01 U2025 ( .Y(n4899), .A(n7736) );
  nor02 U2026 ( .Y(n4896), .A0(n4899), .A1(n4900) );
  nor02 U2027 ( .Y(n4901), .A0(n4897), .A1(n4898) );
  inv01 U2028 ( .Y(n4900), .A(n4901) );
  inv01 U2029 ( .Y(s_output_o[29]), .A(n4902) );
  nor02 U2030 ( .Y(n4903), .A0(n7739), .A1(n7651) );
  nor02 U2031 ( .Y(n4904), .A0(n7738), .A1(n7650) );
  inv01 U2032 ( .Y(n4905), .A(n7736) );
  nor02 U2033 ( .Y(n4902), .A0(n4905), .A1(n4906) );
  nor02 U2034 ( .Y(n4907), .A0(n4903), .A1(n4904) );
  inv01 U2035 ( .Y(n4906), .A(n4907) );
  inv01 U2036 ( .Y(s_output_o[23]), .A(n4908) );
  nor02 U2037 ( .Y(n4909), .A0(n7324), .A1(n7651) );
  nor02 U2038 ( .Y(n4910), .A0(n7750), .A1(n7650) );
  inv01 U2039 ( .Y(n4911), .A(n7736) );
  nor02 U2040 ( .Y(n4908), .A0(n4911), .A1(n4912) );
  nor02 U2041 ( .Y(n4913), .A0(n4909), .A1(n4910) );
  inv01 U2042 ( .Y(n4912), .A(n4913) );
  inv02 U2043 ( .Y(n7736), .A(n7661) );
  inv01 U2044 ( .Y(n7909), .A(n4914) );
  nor02 U2045 ( .Y(n4915), .A0(n7703), .A1(n7911) );
  nor02 U2046 ( .Y(n4916), .A0(n7902), .A1(n7702) );
  inv01 U2047 ( .Y(n4917), .A(n4478) );
  nor02 U2048 ( .Y(n4914), .A0(n4917), .A1(n4918) );
  nor02 U2049 ( .Y(n4919), .A0(n4915), .A1(n4916) );
  inv01 U2050 ( .Y(n4918), .A(n4919) );
  inv01 U2051 ( .Y(n7928), .A(n4920) );
  nor02 U2052 ( .Y(n4921), .A0(n7932), .A1(n7703) );
  nor02 U2053 ( .Y(n4922), .A0(n7922), .A1(n7702) );
  inv01 U2054 ( .Y(n4923), .A(n7933) );
  nor02 U2055 ( .Y(n4920), .A0(n4923), .A1(n4924) );
  nor02 U2056 ( .Y(n4925), .A0(n4921), .A1(n4922) );
  inv01 U2057 ( .Y(n4924), .A(n4925) );
  inv01 U2058 ( .Y(n7898), .A(n4926) );
  nor02 U2059 ( .Y(n4927), .A0(n7902), .A1(n7703) );
  nor02 U2060 ( .Y(n4928), .A0(n7900), .A1(n7702) );
  inv01 U2061 ( .Y(n4929), .A(n4436) );
  nor02 U2062 ( .Y(n4926), .A0(n4929), .A1(n4930) );
  nor02 U2063 ( .Y(n4931), .A0(n4927), .A1(n4928) );
  inv01 U2064 ( .Y(n4930), .A(n4931) );
  inv01 U2065 ( .Y(s_output_o[28]), .A(n4932) );
  nor02 U2066 ( .Y(n4933), .A0(n7741), .A1(n7651) );
  nor02 U2067 ( .Y(n4934), .A0(n7740), .A1(n7650) );
  inv01 U2068 ( .Y(n4935), .A(n7736) );
  nor02 U2069 ( .Y(n4932), .A0(n4935), .A1(n4936) );
  nor02 U2070 ( .Y(n4937), .A0(n4933), .A1(n4934) );
  inv01 U2071 ( .Y(n4936), .A(n4937) );
  nand02 U2072 ( .Y(n8004), .A0(n4938), .A1(n4939) );
  inv02 U2073 ( .Y(n4940), .A(n7830) );
  inv02 U2074 ( .Y(n4941), .A(n7834) );
  inv02 U2075 ( .Y(n4942), .A(n7978) );
  inv02 U2076 ( .Y(n4943), .A(n7626) );
  inv02 U2077 ( .Y(n4944), .A(n7672) );
  inv02 U2078 ( .Y(n4945), .A(n7670) );
  nand02 U2079 ( .Y(n4946), .A0(n4942), .A1(n4947) );
  nand02 U2080 ( .Y(n4948), .A0(n4943), .A1(n4949) );
  nand02 U2081 ( .Y(n4950), .A0(n4944), .A1(n4951) );
  nand02 U2082 ( .Y(n4952), .A0(n4944), .A1(n4953) );
  nand02 U2083 ( .Y(n4954), .A0(n4945), .A1(n4955) );
  nand02 U2084 ( .Y(n4956), .A0(n4945), .A1(n4957) );
  nand02 U2085 ( .Y(n4958), .A0(n4945), .A1(n4959) );
  nand02 U2086 ( .Y(n4960), .A0(n4945), .A1(n4961) );
  nand02 U2087 ( .Y(n4962), .A0(n4940), .A1(n4941) );
  inv01 U2088 ( .Y(n4947), .A(n4962) );
  nand02 U2089 ( .Y(n4963), .A0(n4940), .A1(n4941) );
  inv01 U2090 ( .Y(n4949), .A(n4963) );
  nand02 U2091 ( .Y(n4964), .A0(n4940), .A1(n4942) );
  inv01 U2092 ( .Y(n4951), .A(n4964) );
  nand02 U2093 ( .Y(n4965), .A0(n4940), .A1(n4943) );
  inv01 U2094 ( .Y(n4953), .A(n4965) );
  nand02 U2095 ( .Y(n4966), .A0(n4941), .A1(n4942) );
  inv01 U2096 ( .Y(n4955), .A(n4966) );
  nand02 U2097 ( .Y(n4967), .A0(n4941), .A1(n4943) );
  inv01 U2098 ( .Y(n4957), .A(n4967) );
  nand02 U2099 ( .Y(n4968), .A0(n4942), .A1(n4944) );
  inv01 U2100 ( .Y(n4959), .A(n4968) );
  nand02 U2101 ( .Y(n4969), .A0(n4943), .A1(n4944) );
  inv01 U2102 ( .Y(n4961), .A(n4969) );
  nand02 U2103 ( .Y(n4970), .A0(n4946), .A1(n4948) );
  inv01 U2104 ( .Y(n4971), .A(n4970) );
  nand02 U2105 ( .Y(n4972), .A0(n4950), .A1(n4952) );
  inv01 U2106 ( .Y(n4973), .A(n4972) );
  nand02 U2107 ( .Y(n4974), .A0(n4971), .A1(n4973) );
  inv01 U2108 ( .Y(n4938), .A(n4974) );
  nand02 U2109 ( .Y(n4975), .A0(n4954), .A1(n4956) );
  inv01 U2110 ( .Y(n4976), .A(n4975) );
  nand02 U2111 ( .Y(n4977), .A0(n4958), .A1(n4960) );
  inv01 U2112 ( .Y(n4978), .A(n4977) );
  nand02 U2113 ( .Y(n4979), .A0(n4976), .A1(n4978) );
  inv01 U2114 ( .Y(n4939), .A(n4979) );
  inv01 U2115 ( .Y(n7917), .A(n4980) );
  nor02 U2116 ( .Y(n4981), .A0(n7922), .A1(n7703) );
  nor02 U2117 ( .Y(n4982), .A0(n7702), .A1(n7911) );
  inv01 U2118 ( .Y(n4983), .A(n4331) );
  nor02 U2119 ( .Y(n4980), .A0(n4983), .A1(n4984) );
  nor02 U2120 ( .Y(n4985), .A0(n4981), .A1(n4982) );
  inv01 U2121 ( .Y(n4984), .A(n4985) );
  inv01 U2122 ( .Y(s_output_o[25]), .A(n4986) );
  nor02 U2123 ( .Y(n4987), .A0(n7747), .A1(n7651) );
  nor02 U2124 ( .Y(n4988), .A0(n7746), .A1(n7650) );
  inv01 U2125 ( .Y(n4989), .A(n7736) );
  nor02 U2126 ( .Y(n4986), .A0(n4989), .A1(n4990) );
  nor02 U2127 ( .Y(n4991), .A0(n4987), .A1(n4988) );
  inv01 U2128 ( .Y(n4990), .A(n4991) );
  nand02 U2129 ( .Y(n7895), .A0(n4992), .A1(n4993) );
  inv02 U2130 ( .Y(n4994), .A(n7899) );
  inv02 U2131 ( .Y(n4995), .A(n7898) );
  inv02 U2132 ( .Y(n4996), .A(n7897) );
  inv02 U2133 ( .Y(n4997), .A(n7669) );
  inv02 U2134 ( .Y(n4998), .A(n7678) );
  inv02 U2135 ( .Y(n4999), .A(n7676) );
  nand02 U2136 ( .Y(n5000), .A0(n4996), .A1(n5001) );
  nand02 U2137 ( .Y(n5002), .A0(n4997), .A1(n5003) );
  nand02 U2138 ( .Y(n5004), .A0(n4998), .A1(n5005) );
  nand02 U2139 ( .Y(n5006), .A0(n4998), .A1(n5007) );
  nand02 U2140 ( .Y(n5008), .A0(n4999), .A1(n5009) );
  nand02 U2141 ( .Y(n5010), .A0(n4999), .A1(n5011) );
  nand02 U2142 ( .Y(n5012), .A0(n4999), .A1(n5013) );
  nand02 U2143 ( .Y(n5014), .A0(n4999), .A1(n5015) );
  nand02 U2144 ( .Y(n5016), .A0(n4994), .A1(n4995) );
  inv01 U2145 ( .Y(n5001), .A(n5016) );
  nand02 U2146 ( .Y(n5017), .A0(n4994), .A1(n4995) );
  inv01 U2147 ( .Y(n5003), .A(n5017) );
  nand02 U2148 ( .Y(n5018), .A0(n4994), .A1(n4996) );
  inv01 U2149 ( .Y(n5005), .A(n5018) );
  nand02 U2150 ( .Y(n5019), .A0(n4994), .A1(n4997) );
  inv01 U2151 ( .Y(n5007), .A(n5019) );
  nand02 U2152 ( .Y(n5020), .A0(n4995), .A1(n4996) );
  inv01 U2153 ( .Y(n5009), .A(n5020) );
  nand02 U2154 ( .Y(n5021), .A0(n4995), .A1(n4997) );
  inv01 U2155 ( .Y(n5011), .A(n5021) );
  nand02 U2156 ( .Y(n5022), .A0(n4996), .A1(n4998) );
  inv01 U2157 ( .Y(n5013), .A(n5022) );
  nand02 U2158 ( .Y(n5023), .A0(n4997), .A1(n4998) );
  inv01 U2159 ( .Y(n5015), .A(n5023) );
  nand02 U2160 ( .Y(n5024), .A0(n5000), .A1(n5002) );
  inv01 U2161 ( .Y(n5025), .A(n5024) );
  nand02 U2162 ( .Y(n5026), .A0(n5004), .A1(n5006) );
  inv01 U2163 ( .Y(n5027), .A(n5026) );
  nand02 U2164 ( .Y(n5028), .A0(n5025), .A1(n5027) );
  inv01 U2165 ( .Y(n4992), .A(n5028) );
  nand02 U2166 ( .Y(n5029), .A0(n5008), .A1(n5010) );
  inv01 U2167 ( .Y(n5030), .A(n5029) );
  nand02 U2168 ( .Y(n5031), .A0(n5012), .A1(n5014) );
  inv01 U2169 ( .Y(n5032), .A(n5031) );
  nand02 U2170 ( .Y(n5033), .A0(n5030), .A1(n5032) );
  inv01 U2171 ( .Y(n4993), .A(n5033) );
  nand02 U2172 ( .Y(n7965), .A0(n5034), .A1(n5035) );
  inv02 U2173 ( .Y(n5036), .A(n7857) );
  inv02 U2174 ( .Y(n5037), .A(n7913) );
  inv02 U2175 ( .Y(n5038), .A(n7944) );
  inv02 U2176 ( .Y(n5039), .A(n7669) );
  inv02 U2177 ( .Y(n5040), .A(n7676) );
  nand02 U2178 ( .Y(n5041), .A0(n5038), .A1(n5042) );
  nand02 U2179 ( .Y(n5043), .A0(n5039), .A1(n5044) );
  nand02 U2180 ( .Y(n5045), .A0(n5040), .A1(n5046) );
  nand02 U2181 ( .Y(n5047), .A0(n5040), .A1(n5048) );
  nand02 U2182 ( .Y(n5049), .A0(n5873), .A1(n5050) );
  nand02 U2183 ( .Y(n5051), .A0(n5873), .A1(n5052) );
  nand02 U2184 ( .Y(n5053), .A0(n5873), .A1(n5054) );
  nand02 U2185 ( .Y(n5055), .A0(n5873), .A1(n5056) );
  nand02 U2186 ( .Y(n5057), .A0(n5036), .A1(n5037) );
  inv01 U2187 ( .Y(n5042), .A(n5057) );
  nand02 U2188 ( .Y(n5058), .A0(n5036), .A1(n5037) );
  inv01 U2189 ( .Y(n5044), .A(n5058) );
  nand02 U2190 ( .Y(n5059), .A0(n5036), .A1(n5038) );
  inv01 U2191 ( .Y(n5046), .A(n5059) );
  nand02 U2192 ( .Y(n5060), .A0(n5036), .A1(n5039) );
  inv01 U2193 ( .Y(n5048), .A(n5060) );
  nand02 U2194 ( .Y(n5061), .A0(n5037), .A1(n5038) );
  inv01 U2195 ( .Y(n5050), .A(n5061) );
  nand02 U2196 ( .Y(n5062), .A0(n5037), .A1(n5039) );
  inv01 U2197 ( .Y(n5052), .A(n5062) );
  nand02 U2198 ( .Y(n5063), .A0(n5038), .A1(n5040) );
  inv01 U2199 ( .Y(n5054), .A(n5063) );
  nand02 U2200 ( .Y(n5064), .A0(n5039), .A1(n5040) );
  inv01 U2201 ( .Y(n5056), .A(n5064) );
  nand02 U2202 ( .Y(n5065), .A0(n5041), .A1(n5043) );
  inv01 U2203 ( .Y(n5066), .A(n5065) );
  nand02 U2204 ( .Y(n5067), .A0(n5045), .A1(n5047) );
  inv01 U2205 ( .Y(n5068), .A(n5067) );
  nand02 U2206 ( .Y(n5069), .A0(n5066), .A1(n5068) );
  inv01 U2207 ( .Y(n5034), .A(n5069) );
  nand02 U2208 ( .Y(n5070), .A0(n5049), .A1(n5051) );
  inv01 U2209 ( .Y(n5071), .A(n5070) );
  nand02 U2210 ( .Y(n5072), .A0(n5053), .A1(n5055) );
  inv01 U2211 ( .Y(n5073), .A(n5072) );
  nand02 U2212 ( .Y(n5074), .A0(n5071), .A1(n5073) );
  inv01 U2213 ( .Y(n5035), .A(n5074) );
  inv01 U2214 ( .Y(n7758), .A(n5075) );
  inv01 U2215 ( .Y(n5076), .A(opa_i[12]) );
  inv01 U2216 ( .Y(n5077), .A(opa_i[13]) );
  inv01 U2217 ( .Y(n5078), .A(opa_i[11]) );
  nand02 U2218 ( .Y(n5075), .A0(n5078), .A1(n5079) );
  nand02 U2219 ( .Y(n5080), .A0(n5076), .A1(n5077) );
  inv01 U2220 ( .Y(n5079), .A(n5080) );
  inv01 U2221 ( .Y(s_output_o[27]), .A(n5081) );
  nor02 U2222 ( .Y(n5082), .A0(n7743), .A1(n7651) );
  nor02 U2223 ( .Y(n5083), .A0(n7742), .A1(n7650) );
  inv01 U2224 ( .Y(n5084), .A(n7736) );
  nor02 U2225 ( .Y(n5081), .A0(n5084), .A1(n5085) );
  nor02 U2226 ( .Y(n5086), .A0(n5082), .A1(n5083) );
  inv01 U2227 ( .Y(n5085), .A(n5086) );
  inv01 U2228 ( .Y(s_output_o[24]), .A(n5087) );
  nor02 U2229 ( .Y(n5088), .A0(n7749), .A1(n7651) );
  nor02 U2230 ( .Y(n5089), .A0(n7748), .A1(n7650) );
  inv01 U2231 ( .Y(n5090), .A(n7736) );
  nor02 U2232 ( .Y(n5087), .A0(n5090), .A1(n5091) );
  nor02 U2233 ( .Y(n5092), .A0(n5088), .A1(n5089) );
  inv01 U2234 ( .Y(n5091), .A(n5092) );
  inv01 U2235 ( .Y(s_output_o[30]), .A(n5093) );
  nor02 U2236 ( .Y(n5094), .A0(n7734), .A1(n7651) );
  nor02 U2237 ( .Y(n5095), .A0(n7732), .A1(n7650) );
  inv01 U2238 ( .Y(n5096), .A(n7736) );
  nor02 U2239 ( .Y(n5093), .A0(n5096), .A1(n5097) );
  nor02 U2240 ( .Y(n5098), .A0(n5094), .A1(n5095) );
  inv01 U2241 ( .Y(n5097), .A(n5098) );
  buf04 U2242 ( .Y(n7651), .A(n7735) );
  nand02 U2243 ( .Y(n7828), .A0(n5099), .A1(n5100) );
  inv02 U2244 ( .Y(n5101), .A(n7835) );
  inv02 U2245 ( .Y(n5102), .A(n7834) );
  inv02 U2246 ( .Y(n5103), .A(n7833) );
  inv02 U2247 ( .Y(n5104), .A(n7670) );
  inv02 U2248 ( .Y(n5105), .A(n7677) );
  inv02 U2249 ( .Y(n5106), .A(n7673) );
  nand02 U2250 ( .Y(n5107), .A0(n5103), .A1(n5108) );
  nand02 U2251 ( .Y(n5109), .A0(n5104), .A1(n5110) );
  nand02 U2252 ( .Y(n5111), .A0(n5105), .A1(n5112) );
  nand02 U2253 ( .Y(n5113), .A0(n5105), .A1(n5114) );
  nand02 U2254 ( .Y(n5115), .A0(n5106), .A1(n5116) );
  nand02 U2255 ( .Y(n5117), .A0(n5106), .A1(n5118) );
  nand02 U2256 ( .Y(n5119), .A0(n5106), .A1(n5120) );
  nand02 U2257 ( .Y(n5121), .A0(n5106), .A1(n5122) );
  nand02 U2258 ( .Y(n5123), .A0(n5101), .A1(n5102) );
  inv01 U2259 ( .Y(n5108), .A(n5123) );
  nand02 U2260 ( .Y(n5124), .A0(n5101), .A1(n5102) );
  inv01 U2261 ( .Y(n5110), .A(n5124) );
  nand02 U2262 ( .Y(n5125), .A0(n5101), .A1(n5103) );
  inv01 U2263 ( .Y(n5112), .A(n5125) );
  nand02 U2264 ( .Y(n5126), .A0(n5101), .A1(n5104) );
  inv01 U2265 ( .Y(n5114), .A(n5126) );
  nand02 U2266 ( .Y(n5127), .A0(n5102), .A1(n5103) );
  inv01 U2267 ( .Y(n5116), .A(n5127) );
  nand02 U2268 ( .Y(n5128), .A0(n5102), .A1(n5104) );
  inv01 U2269 ( .Y(n5118), .A(n5128) );
  nand02 U2270 ( .Y(n5129), .A0(n5103), .A1(n5105) );
  inv01 U2271 ( .Y(n5120), .A(n5129) );
  nand02 U2272 ( .Y(n5130), .A0(n5104), .A1(n5105) );
  inv01 U2273 ( .Y(n5122), .A(n5130) );
  nand02 U2274 ( .Y(n5131), .A0(n5107), .A1(n5109) );
  inv01 U2275 ( .Y(n5132), .A(n5131) );
  nand02 U2276 ( .Y(n5133), .A0(n5111), .A1(n5113) );
  inv01 U2277 ( .Y(n5134), .A(n5133) );
  nand02 U2278 ( .Y(n5135), .A0(n5132), .A1(n5134) );
  inv01 U2279 ( .Y(n5099), .A(n5135) );
  nand02 U2280 ( .Y(n5136), .A0(n5115), .A1(n5117) );
  inv01 U2281 ( .Y(n5137), .A(n5136) );
  nand02 U2282 ( .Y(n5138), .A0(n5119), .A1(n5121) );
  inv01 U2283 ( .Y(n5139), .A(n5138) );
  nand02 U2284 ( .Y(n5140), .A0(n5137), .A1(n5139) );
  inv01 U2285 ( .Y(n5100), .A(n5140) );
  nand02 U2286 ( .Y(n7997), .A0(n5141), .A1(n5142) );
  inv02 U2287 ( .Y(n5143), .A(n7852) );
  inv02 U2288 ( .Y(n5144), .A(n7912) );
  inv02 U2289 ( .Y(n5145), .A(n7858) );
  inv02 U2290 ( .Y(n5146), .A(n7670) );
  inv02 U2291 ( .Y(n5147), .A(n7657) );
  inv02 U2292 ( .Y(n5148), .A(n7673) );
  nand02 U2293 ( .Y(n5149), .A0(n5145), .A1(n5150) );
  nand02 U2294 ( .Y(n5151), .A0(n5146), .A1(n5152) );
  nand02 U2295 ( .Y(n5153), .A0(n5147), .A1(n5154) );
  nand02 U2296 ( .Y(n5155), .A0(n5147), .A1(n5156) );
  nand02 U2297 ( .Y(n5157), .A0(n5148), .A1(n5158) );
  nand02 U2298 ( .Y(n5159), .A0(n5148), .A1(n5160) );
  nand02 U2299 ( .Y(n5161), .A0(n5148), .A1(n5162) );
  nand02 U2300 ( .Y(n5163), .A0(n5148), .A1(n5164) );
  nand02 U2301 ( .Y(n5165), .A0(n5143), .A1(n5144) );
  inv01 U2302 ( .Y(n5150), .A(n5165) );
  nand02 U2303 ( .Y(n5166), .A0(n5143), .A1(n5144) );
  inv01 U2304 ( .Y(n5152), .A(n5166) );
  nand02 U2305 ( .Y(n5167), .A0(n5143), .A1(n5145) );
  inv01 U2306 ( .Y(n5154), .A(n5167) );
  nand02 U2307 ( .Y(n5168), .A0(n5143), .A1(n5146) );
  inv01 U2308 ( .Y(n5156), .A(n5168) );
  nand02 U2309 ( .Y(n5169), .A0(n5144), .A1(n5145) );
  inv01 U2310 ( .Y(n5158), .A(n5169) );
  nand02 U2311 ( .Y(n5170), .A0(n5144), .A1(n5146) );
  inv01 U2312 ( .Y(n5160), .A(n5170) );
  nand02 U2313 ( .Y(n5171), .A0(n5145), .A1(n5147) );
  inv01 U2314 ( .Y(n5162), .A(n5171) );
  nand02 U2315 ( .Y(n5172), .A0(n5146), .A1(n5147) );
  inv01 U2316 ( .Y(n5164), .A(n5172) );
  nand02 U2317 ( .Y(n5173), .A0(n5149), .A1(n5151) );
  inv01 U2318 ( .Y(n5174), .A(n5173) );
  nand02 U2319 ( .Y(n5175), .A0(n5153), .A1(n5155) );
  inv01 U2320 ( .Y(n5176), .A(n5175) );
  nand02 U2321 ( .Y(n5177), .A0(n5174), .A1(n5176) );
  inv01 U2322 ( .Y(n5141), .A(n5177) );
  nand02 U2323 ( .Y(n5178), .A0(n5157), .A1(n5159) );
  inv01 U2324 ( .Y(n5179), .A(n5178) );
  nand02 U2325 ( .Y(n5180), .A0(n5161), .A1(n5163) );
  inv01 U2326 ( .Y(n5181), .A(n5180) );
  nand02 U2327 ( .Y(n5182), .A0(n5179), .A1(n5181) );
  inv01 U2328 ( .Y(n5142), .A(n5182) );
  nand02 U2329 ( .Y(n7992), .A0(n5183), .A1(n5184) );
  inv02 U2330 ( .Y(n5185), .A(n7963) );
  inv02 U2331 ( .Y(n5186), .A(n7890) );
  inv02 U2332 ( .Y(n5187), .A(n7839) );
  inv02 U2333 ( .Y(n5188), .A(n7670) );
  inv02 U2334 ( .Y(n5189), .A(n7659) );
  inv02 U2335 ( .Y(n5190), .A(n7671) );
  nand02 U2336 ( .Y(n5191), .A0(n5187), .A1(n5192) );
  nand02 U2337 ( .Y(n5193), .A0(n5188), .A1(n5194) );
  nand02 U2338 ( .Y(n5195), .A0(n5189), .A1(n5196) );
  nand02 U2339 ( .Y(n5197), .A0(n5189), .A1(n5198) );
  nand02 U2340 ( .Y(n5199), .A0(n5190), .A1(n5200) );
  nand02 U2341 ( .Y(n5201), .A0(n5190), .A1(n5202) );
  nand02 U2342 ( .Y(n5203), .A0(n5190), .A1(n5204) );
  nand02 U2343 ( .Y(n5205), .A0(n5190), .A1(n5206) );
  nand02 U2344 ( .Y(n5207), .A0(n5185), .A1(n5186) );
  inv01 U2345 ( .Y(n5192), .A(n5207) );
  nand02 U2346 ( .Y(n5208), .A0(n5185), .A1(n5186) );
  inv01 U2347 ( .Y(n5194), .A(n5208) );
  nand02 U2348 ( .Y(n5209), .A0(n5185), .A1(n5187) );
  inv01 U2349 ( .Y(n5196), .A(n5209) );
  nand02 U2350 ( .Y(n5210), .A0(n5185), .A1(n5188) );
  inv01 U2351 ( .Y(n5198), .A(n5210) );
  nand02 U2352 ( .Y(n5211), .A0(n5186), .A1(n5187) );
  inv01 U2353 ( .Y(n5200), .A(n5211) );
  nand02 U2354 ( .Y(n5212), .A0(n5186), .A1(n5188) );
  inv01 U2355 ( .Y(n5202), .A(n5212) );
  nand02 U2356 ( .Y(n5213), .A0(n5187), .A1(n5189) );
  inv01 U2357 ( .Y(n5204), .A(n5213) );
  nand02 U2358 ( .Y(n5214), .A0(n5188), .A1(n5189) );
  inv01 U2359 ( .Y(n5206), .A(n5214) );
  nand02 U2360 ( .Y(n5215), .A0(n5191), .A1(n5193) );
  inv01 U2361 ( .Y(n5216), .A(n5215) );
  nand02 U2362 ( .Y(n5217), .A0(n5195), .A1(n5197) );
  inv01 U2363 ( .Y(n5218), .A(n5217) );
  nand02 U2364 ( .Y(n5219), .A0(n5216), .A1(n5218) );
  inv01 U2365 ( .Y(n5183), .A(n5219) );
  nand02 U2366 ( .Y(n5220), .A0(n5199), .A1(n5201) );
  inv01 U2367 ( .Y(n5221), .A(n5220) );
  nand02 U2368 ( .Y(n5222), .A0(n5203), .A1(n5205) );
  inv01 U2369 ( .Y(n5223), .A(n5222) );
  nand02 U2370 ( .Y(n5224), .A0(n5221), .A1(n5223) );
  inv01 U2371 ( .Y(n5184), .A(n5224) );
  nand02 U2372 ( .Y(n7883), .A0(n5225), .A1(n5226) );
  inv02 U2373 ( .Y(n5227), .A(n7856) );
  inv02 U2374 ( .Y(n5228), .A(n7855) );
  inv02 U2375 ( .Y(n5229), .A(n7854) );
  inv02 U2376 ( .Y(n5230), .A(n7678) );
  inv02 U2377 ( .Y(n5231), .A(n7670) );
  inv02 U2378 ( .Y(n5232), .A(n7671) );
  nand02 U2379 ( .Y(n5233), .A0(n5229), .A1(n5234) );
  nand02 U2380 ( .Y(n5235), .A0(n5230), .A1(n5236) );
  nand02 U2381 ( .Y(n5237), .A0(n5231), .A1(n5238) );
  nand02 U2382 ( .Y(n5239), .A0(n5231), .A1(n5240) );
  nand02 U2383 ( .Y(n5241), .A0(n5232), .A1(n5242) );
  nand02 U2384 ( .Y(n5243), .A0(n5232), .A1(n5244) );
  nand02 U2385 ( .Y(n5245), .A0(n5232), .A1(n5246) );
  nand02 U2386 ( .Y(n5247), .A0(n5232), .A1(n5248) );
  nand02 U2387 ( .Y(n5249), .A0(n5227), .A1(n5228) );
  inv01 U2388 ( .Y(n5234), .A(n5249) );
  nand02 U2389 ( .Y(n5250), .A0(n5227), .A1(n5228) );
  inv01 U2390 ( .Y(n5236), .A(n5250) );
  nand02 U2391 ( .Y(n5251), .A0(n5227), .A1(n5229) );
  inv01 U2392 ( .Y(n5238), .A(n5251) );
  nand02 U2393 ( .Y(n5252), .A0(n5227), .A1(n5230) );
  inv01 U2394 ( .Y(n5240), .A(n5252) );
  nand02 U2395 ( .Y(n5253), .A0(n5228), .A1(n5229) );
  inv01 U2396 ( .Y(n5242), .A(n5253) );
  nand02 U2397 ( .Y(n5254), .A0(n5228), .A1(n5230) );
  inv01 U2398 ( .Y(n5244), .A(n5254) );
  nand02 U2399 ( .Y(n5255), .A0(n5229), .A1(n5231) );
  inv01 U2400 ( .Y(n5246), .A(n5255) );
  nand02 U2401 ( .Y(n5256), .A0(n5230), .A1(n5231) );
  inv01 U2402 ( .Y(n5248), .A(n5256) );
  nand02 U2403 ( .Y(n5257), .A0(n5233), .A1(n5235) );
  inv01 U2404 ( .Y(n5258), .A(n5257) );
  nand02 U2405 ( .Y(n5259), .A0(n5237), .A1(n5239) );
  inv01 U2406 ( .Y(n5260), .A(n5259) );
  nand02 U2407 ( .Y(n5261), .A0(n5258), .A1(n5260) );
  inv01 U2408 ( .Y(n5225), .A(n5261) );
  nand02 U2409 ( .Y(n5262), .A0(n5241), .A1(n5243) );
  inv01 U2410 ( .Y(n5263), .A(n5262) );
  nand02 U2411 ( .Y(n5264), .A0(n5245), .A1(n5247) );
  inv01 U2412 ( .Y(n5265), .A(n5264) );
  nand02 U2413 ( .Y(n5266), .A0(n5263), .A1(n5265) );
  inv01 U2414 ( .Y(n5226), .A(n5266) );
  nand02 U2415 ( .Y(n8012), .A0(n5267), .A1(n5268) );
  inv02 U2416 ( .Y(n5269), .A(n7578) );
  inv02 U2417 ( .Y(n5270), .A(n7649) );
  inv02 U2418 ( .Y(n5271), .A(n7833) );
  inv02 U2419 ( .Y(n5272), .A(n7831) );
  inv02 U2420 ( .Y(n5273), .A(n7835) );
  nand02 U2421 ( .Y(n5274), .A0(n5270), .A1(n5275) );
  nand02 U2422 ( .Y(n5276), .A0(n5271), .A1(n5277) );
  nand02 U2423 ( .Y(n5278), .A0(n5272), .A1(n5279) );
  nand02 U2424 ( .Y(n5280), .A0(n5272), .A1(n5281) );
  nand02 U2425 ( .Y(n5282), .A0(n5273), .A1(n5283) );
  nand02 U2426 ( .Y(n5284), .A0(n5273), .A1(n5285) );
  nand02 U2427 ( .Y(n5286), .A0(n5273), .A1(n5287) );
  nand02 U2428 ( .Y(n5288), .A0(n5273), .A1(n5289) );
  nand02 U2429 ( .Y(n5290), .A0(n6051), .A1(n5269) );
  inv01 U2430 ( .Y(n5275), .A(n5290) );
  nand02 U2431 ( .Y(n5291), .A0(n6219), .A1(n5269) );
  inv01 U2432 ( .Y(n5277), .A(n5291) );
  nand02 U2433 ( .Y(n5292), .A0(n6092), .A1(n5270) );
  inv01 U2434 ( .Y(n5279), .A(n5292) );
  nand02 U2435 ( .Y(n5293), .A0(n6092), .A1(n5271) );
  inv01 U2436 ( .Y(n5281), .A(n5293) );
  nand02 U2437 ( .Y(n5294), .A0(n5269), .A1(n5270) );
  inv01 U2438 ( .Y(n5283), .A(n5294) );
  nand02 U2439 ( .Y(n5295), .A0(n5269), .A1(n5271) );
  inv01 U2440 ( .Y(n5285), .A(n5295) );
  nand02 U2441 ( .Y(n5296), .A0(n5270), .A1(n5272) );
  inv01 U2442 ( .Y(n5287), .A(n5296) );
  nand02 U2443 ( .Y(n5297), .A0(n5271), .A1(n5272) );
  inv01 U2444 ( .Y(n5289), .A(n5297) );
  nand02 U2445 ( .Y(n5298), .A0(n5274), .A1(n5276) );
  inv01 U2446 ( .Y(n5299), .A(n5298) );
  nand02 U2447 ( .Y(n5300), .A0(n5278), .A1(n5280) );
  inv01 U2448 ( .Y(n5301), .A(n5300) );
  nand02 U2449 ( .Y(n5302), .A0(n5299), .A1(n5301) );
  inv01 U2450 ( .Y(n5267), .A(n5302) );
  nand02 U2451 ( .Y(n5303), .A0(n5282), .A1(n5284) );
  inv01 U2452 ( .Y(n5304), .A(n5303) );
  nand02 U2453 ( .Y(n5305), .A0(n5286), .A1(n5288) );
  inv01 U2454 ( .Y(n5306), .A(n5305) );
  nand02 U2455 ( .Y(n5307), .A0(n5304), .A1(n5306) );
  inv01 U2456 ( .Y(n5268), .A(n5307) );
  nand02 U2457 ( .Y(n8001), .A0(n5308), .A1(n5309) );
  inv02 U2458 ( .Y(n5310), .A(n7586) );
  inv02 U2459 ( .Y(n5311), .A(n7639) );
  inv02 U2460 ( .Y(n5312), .A(n7944) );
  inv02 U2461 ( .Y(n5313), .A(n7854) );
  inv02 U2462 ( .Y(n5314), .A(n7857) );
  nand02 U2463 ( .Y(n5315), .A0(n5311), .A1(n5316) );
  nand02 U2464 ( .Y(n5317), .A0(n5312), .A1(n5318) );
  nand02 U2465 ( .Y(n5319), .A0(n5313), .A1(n5320) );
  nand02 U2466 ( .Y(n5321), .A0(n5313), .A1(n5322) );
  nand02 U2467 ( .Y(n5323), .A0(n5314), .A1(n5324) );
  nand02 U2468 ( .Y(n5325), .A0(n5314), .A1(n5326) );
  nand02 U2469 ( .Y(n5327), .A0(n5314), .A1(n5328) );
  nand02 U2470 ( .Y(n5329), .A0(n5314), .A1(n5330) );
  nand02 U2471 ( .Y(n5331), .A0(n6471), .A1(n5310) );
  inv01 U2472 ( .Y(n5316), .A(n5331) );
  nand02 U2473 ( .Y(n5332), .A0(n6429), .A1(n5310) );
  inv01 U2474 ( .Y(n5318), .A(n5332) );
  nand02 U2475 ( .Y(n5333), .A0(n5736), .A1(n5311) );
  inv01 U2476 ( .Y(n5320), .A(n5333) );
  nand02 U2477 ( .Y(n5334), .A0(n5736), .A1(n5312) );
  inv01 U2478 ( .Y(n5322), .A(n5334) );
  nand02 U2479 ( .Y(n5335), .A0(n5310), .A1(n5311) );
  inv01 U2480 ( .Y(n5324), .A(n5335) );
  nand02 U2481 ( .Y(n5336), .A0(n5310), .A1(n5312) );
  inv01 U2482 ( .Y(n5326), .A(n5336) );
  nand02 U2483 ( .Y(n5337), .A0(n5311), .A1(n5313) );
  inv01 U2484 ( .Y(n5328), .A(n5337) );
  nand02 U2485 ( .Y(n5338), .A0(n5312), .A1(n5313) );
  inv01 U2486 ( .Y(n5330), .A(n5338) );
  nand02 U2487 ( .Y(n5339), .A0(n5315), .A1(n5317) );
  inv01 U2488 ( .Y(n5340), .A(n5339) );
  nand02 U2489 ( .Y(n5341), .A0(n5319), .A1(n5321) );
  inv01 U2490 ( .Y(n5342), .A(n5341) );
  nand02 U2491 ( .Y(n5343), .A0(n5340), .A1(n5342) );
  inv01 U2492 ( .Y(n5308), .A(n5343) );
  nand02 U2493 ( .Y(n5344), .A0(n5323), .A1(n5325) );
  inv01 U2494 ( .Y(n5345), .A(n5344) );
  nand02 U2495 ( .Y(n5346), .A0(n5327), .A1(n5329) );
  inv01 U2496 ( .Y(n5347), .A(n5346) );
  nand02 U2497 ( .Y(n5348), .A0(n5345), .A1(n5347) );
  inv01 U2498 ( .Y(n5309), .A(n5348) );
  inv01 U2499 ( .Y(n7762), .A(n5349) );
  inv01 U2500 ( .Y(n5350), .A(opa_i[2]) );
  inv01 U2501 ( .Y(n5351), .A(opa_i[3]) );
  inv01 U2502 ( .Y(n5352), .A(opa_i[22]) );
  nand02 U2503 ( .Y(n5349), .A0(n5352), .A1(n5353) );
  nand02 U2504 ( .Y(n5354), .A0(n5350), .A1(n5351) );
  inv01 U2505 ( .Y(n5353), .A(n5354) );
  inv02 U2506 ( .Y(n7944), .A(n7432) );
  inv02 U2507 ( .Y(n7857), .A(n7551) );
  nand02 U2508 ( .Y(n7906), .A0(n5355), .A1(n5356) );
  inv02 U2509 ( .Y(n5357), .A(n7913) );
  inv02 U2510 ( .Y(n5358), .A(n7912) );
  inv02 U2511 ( .Y(n5359), .A(n7601) );
  inv02 U2512 ( .Y(n5360), .A(n7675) );
  inv02 U2513 ( .Y(n5361), .A(n7647) );
  nand02 U2514 ( .Y(n5362), .A0(n5359), .A1(n5363) );
  nand02 U2515 ( .Y(n5364), .A0(n5360), .A1(n5365) );
  nand02 U2516 ( .Y(n5366), .A0(n5361), .A1(n5367) );
  nand02 U2517 ( .Y(n5368), .A0(n5361), .A1(n5369) );
  nand02 U2518 ( .Y(n5370), .A0(n5873), .A1(n5371) );
  nand02 U2519 ( .Y(n5372), .A0(n5873), .A1(n5373) );
  nand02 U2520 ( .Y(n5374), .A0(n5873), .A1(n5375) );
  nand02 U2521 ( .Y(n5376), .A0(n5873), .A1(n5377) );
  nand02 U2522 ( .Y(n5378), .A0(n5357), .A1(n5358) );
  inv01 U2523 ( .Y(n5363), .A(n5378) );
  nand02 U2524 ( .Y(n5379), .A0(n5357), .A1(n5358) );
  inv01 U2525 ( .Y(n5365), .A(n5379) );
  nand02 U2526 ( .Y(n5380), .A0(n5357), .A1(n5359) );
  inv01 U2527 ( .Y(n5367), .A(n5380) );
  nand02 U2528 ( .Y(n5381), .A0(n5357), .A1(n5360) );
  inv01 U2529 ( .Y(n5369), .A(n5381) );
  nand02 U2530 ( .Y(n5382), .A0(n5358), .A1(n5359) );
  inv01 U2531 ( .Y(n5371), .A(n5382) );
  nand02 U2532 ( .Y(n5383), .A0(n5358), .A1(n5360) );
  inv01 U2533 ( .Y(n5373), .A(n5383) );
  nand02 U2534 ( .Y(n5384), .A0(n5359), .A1(n5361) );
  inv01 U2535 ( .Y(n5375), .A(n5384) );
  nand02 U2536 ( .Y(n5385), .A0(n5360), .A1(n5361) );
  inv01 U2537 ( .Y(n5377), .A(n5385) );
  nand02 U2538 ( .Y(n5386), .A0(n5362), .A1(n5364) );
  inv01 U2539 ( .Y(n5387), .A(n5386) );
  nand02 U2540 ( .Y(n5388), .A0(n5366), .A1(n5368) );
  inv01 U2541 ( .Y(n5389), .A(n5388) );
  nand02 U2542 ( .Y(n5390), .A0(n5387), .A1(n5389) );
  inv01 U2543 ( .Y(n5355), .A(n5390) );
  nand02 U2544 ( .Y(n5391), .A0(n5370), .A1(n5372) );
  inv01 U2545 ( .Y(n5392), .A(n5391) );
  nand02 U2546 ( .Y(n5393), .A0(n5374), .A1(n5376) );
  inv01 U2547 ( .Y(n5394), .A(n5393) );
  nand02 U2548 ( .Y(n5395), .A0(n5392), .A1(n5394) );
  inv01 U2549 ( .Y(n5356), .A(n5395) );
  nand02 U2550 ( .Y(n7972), .A0(n5396), .A1(n5397) );
  inv02 U2551 ( .Y(n5398), .A(n7935) );
  inv02 U2552 ( .Y(n5399), .A(n7931) );
  inv02 U2553 ( .Y(n5400), .A(n7978) );
  inv02 U2554 ( .Y(n5401), .A(n7653) );
  inv02 U2555 ( .Y(n5402), .A(n7668) );
  inv02 U2556 ( .Y(n5403), .A(n7676) );
  nand02 U2557 ( .Y(n5404), .A0(n5400), .A1(n5405) );
  nand02 U2558 ( .Y(n5406), .A0(n5401), .A1(n5407) );
  nand02 U2559 ( .Y(n5408), .A0(n5402), .A1(n5409) );
  nand02 U2560 ( .Y(n5410), .A0(n5402), .A1(n5411) );
  nand02 U2561 ( .Y(n5412), .A0(n5403), .A1(n5413) );
  nand02 U2562 ( .Y(n5414), .A0(n5403), .A1(n5415) );
  nand02 U2563 ( .Y(n5416), .A0(n5403), .A1(n5417) );
  nand02 U2564 ( .Y(n5418), .A0(n5403), .A1(n5419) );
  nand02 U2565 ( .Y(n5420), .A0(n5398), .A1(n5399) );
  inv01 U2566 ( .Y(n5405), .A(n5420) );
  nand02 U2567 ( .Y(n5421), .A0(n5398), .A1(n5399) );
  inv01 U2568 ( .Y(n5407), .A(n5421) );
  nand02 U2569 ( .Y(n5422), .A0(n5398), .A1(n5400) );
  inv01 U2570 ( .Y(n5409), .A(n5422) );
  nand02 U2571 ( .Y(n5423), .A0(n5398), .A1(n5401) );
  inv01 U2572 ( .Y(n5411), .A(n5423) );
  nand02 U2573 ( .Y(n5424), .A0(n5399), .A1(n5400) );
  inv01 U2574 ( .Y(n5413), .A(n5424) );
  nand02 U2575 ( .Y(n5425), .A0(n5399), .A1(n5401) );
  inv01 U2576 ( .Y(n5415), .A(n5425) );
  nand02 U2577 ( .Y(n5426), .A0(n5400), .A1(n5402) );
  inv01 U2578 ( .Y(n5417), .A(n5426) );
  nand02 U2579 ( .Y(n5427), .A0(n5401), .A1(n5402) );
  inv01 U2580 ( .Y(n5419), .A(n5427) );
  nand02 U2581 ( .Y(n5428), .A0(n5404), .A1(n5406) );
  inv01 U2582 ( .Y(n5429), .A(n5428) );
  nand02 U2583 ( .Y(n5430), .A0(n5408), .A1(n5410) );
  inv01 U2584 ( .Y(n5431), .A(n5430) );
  nand02 U2585 ( .Y(n5432), .A0(n5429), .A1(n5431) );
  inv01 U2586 ( .Y(n5396), .A(n5432) );
  nand02 U2587 ( .Y(n5433), .A0(n5412), .A1(n5414) );
  inv01 U2588 ( .Y(n5434), .A(n5433) );
  nand02 U2589 ( .Y(n5435), .A0(n5416), .A1(n5418) );
  inv01 U2590 ( .Y(n5436), .A(n5435) );
  nand02 U2591 ( .Y(n5437), .A0(n5434), .A1(n5436) );
  inv01 U2592 ( .Y(n5397), .A(n5437) );
  inv02 U2593 ( .Y(n7912), .A(n8001) );
  inv02 U2594 ( .Y(n7978), .A(n8012) );
  nand02 U2595 ( .Y(n7951), .A0(n5438), .A1(n5439) );
  inv02 U2596 ( .Y(n5440), .A(n7861) );
  inv02 U2597 ( .Y(n5441), .A(n7958) );
  inv02 U2598 ( .Y(n5442), .A(n7823) );
  inv02 U2599 ( .Y(n5443), .A(n7672) );
  inv02 U2600 ( .Y(n5444), .A(n7625) );
  inv02 U2601 ( .Y(n5445), .A(n7678) );
  nand02 U2602 ( .Y(n5446), .A0(n5442), .A1(n5447) );
  nand02 U2603 ( .Y(n5448), .A0(n5443), .A1(n5449) );
  nand02 U2604 ( .Y(n5450), .A0(n5444), .A1(n5451) );
  nand02 U2605 ( .Y(n5452), .A0(n5444), .A1(n5453) );
  nand02 U2606 ( .Y(n5454), .A0(n5445), .A1(n5455) );
  nand02 U2607 ( .Y(n5456), .A0(n5445), .A1(n5457) );
  nand02 U2608 ( .Y(n5458), .A0(n5445), .A1(n5459) );
  nand02 U2609 ( .Y(n5460), .A0(n5445), .A1(n5461) );
  nand02 U2610 ( .Y(n5462), .A0(n5440), .A1(n5441) );
  inv01 U2611 ( .Y(n5447), .A(n5462) );
  nand02 U2612 ( .Y(n5463), .A0(n5440), .A1(n5441) );
  inv01 U2613 ( .Y(n5449), .A(n5463) );
  nand02 U2614 ( .Y(n5464), .A0(n5440), .A1(n5442) );
  inv01 U2615 ( .Y(n5451), .A(n5464) );
  nand02 U2616 ( .Y(n5465), .A0(n5440), .A1(n5443) );
  inv01 U2617 ( .Y(n5453), .A(n5465) );
  nand02 U2618 ( .Y(n5466), .A0(n5441), .A1(n5442) );
  inv01 U2619 ( .Y(n5455), .A(n5466) );
  nand02 U2620 ( .Y(n5467), .A0(n5441), .A1(n5443) );
  inv01 U2621 ( .Y(n5457), .A(n5467) );
  nand02 U2622 ( .Y(n5468), .A0(n5442), .A1(n5444) );
  inv01 U2623 ( .Y(n5459), .A(n5468) );
  nand02 U2624 ( .Y(n5469), .A0(n5443), .A1(n5444) );
  inv01 U2625 ( .Y(n5461), .A(n5469) );
  nand02 U2626 ( .Y(n5470), .A0(n5446), .A1(n5448) );
  inv01 U2627 ( .Y(n5471), .A(n5470) );
  nand02 U2628 ( .Y(n5472), .A0(n5450), .A1(n5452) );
  inv01 U2629 ( .Y(n5473), .A(n5472) );
  nand02 U2630 ( .Y(n5474), .A0(n5471), .A1(n5473) );
  inv01 U2631 ( .Y(n5438), .A(n5474) );
  nand02 U2632 ( .Y(n5475), .A0(n5454), .A1(n5456) );
  inv01 U2633 ( .Y(n5476), .A(n5475) );
  nand02 U2634 ( .Y(n5477), .A0(n5458), .A1(n5460) );
  inv01 U2635 ( .Y(n5478), .A(n5477) );
  nand02 U2636 ( .Y(n5479), .A0(n5476), .A1(n5478) );
  inv01 U2637 ( .Y(n5439), .A(n5479) );
  nand02 U2638 ( .Y(n7914), .A0(n5480), .A1(n5481) );
  inv02 U2639 ( .Y(n5482), .A(n7924) );
  inv02 U2640 ( .Y(n5483), .A(n7923) );
  inv02 U2641 ( .Y(n5484), .A(n7819) );
  inv02 U2642 ( .Y(n5485), .A(n7675) );
  inv02 U2643 ( .Y(n5486), .A(n7668) );
  nand02 U2644 ( .Y(n5487), .A0(n5484), .A1(n5488) );
  nand02 U2645 ( .Y(n5489), .A0(n5485), .A1(n5490) );
  nand02 U2646 ( .Y(n5491), .A0(n5486), .A1(n5492) );
  nand02 U2647 ( .Y(n5493), .A0(n5486), .A1(n5494) );
  nand02 U2648 ( .Y(n5495), .A0(n5873), .A1(n5496) );
  nand02 U2649 ( .Y(n5497), .A0(n5873), .A1(n5498) );
  nand02 U2650 ( .Y(n5499), .A0(n5873), .A1(n5500) );
  nand02 U2651 ( .Y(n5501), .A0(n5873), .A1(n5502) );
  nand02 U2652 ( .Y(n5503), .A0(n5482), .A1(n5483) );
  inv01 U2653 ( .Y(n5488), .A(n5503) );
  nand02 U2654 ( .Y(n5504), .A0(n5482), .A1(n5483) );
  inv01 U2655 ( .Y(n5490), .A(n5504) );
  nand02 U2656 ( .Y(n5505), .A0(n5482), .A1(n5484) );
  inv01 U2657 ( .Y(n5492), .A(n5505) );
  nand02 U2658 ( .Y(n5506), .A0(n5482), .A1(n5485) );
  inv01 U2659 ( .Y(n5494), .A(n5506) );
  nand02 U2660 ( .Y(n5507), .A0(n5483), .A1(n5484) );
  inv01 U2661 ( .Y(n5496), .A(n5507) );
  nand02 U2662 ( .Y(n5508), .A0(n5483), .A1(n5485) );
  inv01 U2663 ( .Y(n5498), .A(n5508) );
  nand02 U2664 ( .Y(n5509), .A0(n5484), .A1(n5486) );
  inv01 U2665 ( .Y(n5500), .A(n5509) );
  nand02 U2666 ( .Y(n5510), .A0(n5485), .A1(n5486) );
  inv01 U2667 ( .Y(n5502), .A(n5510) );
  nand02 U2668 ( .Y(n5511), .A0(n5487), .A1(n5489) );
  inv01 U2669 ( .Y(n5512), .A(n5511) );
  nand02 U2670 ( .Y(n5513), .A0(n5491), .A1(n5493) );
  inv01 U2671 ( .Y(n5514), .A(n5513) );
  nand02 U2672 ( .Y(n5515), .A0(n5512), .A1(n5514) );
  inv01 U2673 ( .Y(n5480), .A(n5515) );
  nand02 U2674 ( .Y(n5516), .A0(n5495), .A1(n5497) );
  inv01 U2675 ( .Y(n5517), .A(n5516) );
  nand02 U2676 ( .Y(n5518), .A0(n5499), .A1(n5501) );
  inv01 U2677 ( .Y(n5519), .A(n5518) );
  nand02 U2678 ( .Y(n5520), .A0(n5517), .A1(n5519) );
  inv01 U2679 ( .Y(n5481), .A(n5520) );
  nand02 U2680 ( .Y(n7869), .A0(n5521), .A1(n5522) );
  inv02 U2681 ( .Y(n5523), .A(n7840) );
  inv02 U2682 ( .Y(n5524), .A(n7849) );
  inv02 U2683 ( .Y(n5525), .A(n7848) );
  inv02 U2684 ( .Y(n5526), .A(n7678) );
  inv02 U2685 ( .Y(n5527), .A(n7670) );
  inv02 U2686 ( .Y(n5528), .A(n7672) );
  nand02 U2687 ( .Y(n5529), .A0(n5525), .A1(n5530) );
  nand02 U2688 ( .Y(n5531), .A0(n5526), .A1(n5532) );
  nand02 U2689 ( .Y(n5533), .A0(n5527), .A1(n5534) );
  nand02 U2690 ( .Y(n5535), .A0(n5527), .A1(n5536) );
  nand02 U2691 ( .Y(n5537), .A0(n5528), .A1(n5538) );
  nand02 U2692 ( .Y(n5539), .A0(n5528), .A1(n5540) );
  nand02 U2693 ( .Y(n5541), .A0(n5528), .A1(n5542) );
  nand02 U2694 ( .Y(n5543), .A0(n5528), .A1(n5544) );
  nand02 U2695 ( .Y(n5545), .A0(n5523), .A1(n5524) );
  inv01 U2696 ( .Y(n5530), .A(n5545) );
  nand02 U2697 ( .Y(n5546), .A0(n5523), .A1(n5524) );
  inv01 U2698 ( .Y(n5532), .A(n5546) );
  nand02 U2699 ( .Y(n5547), .A0(n5523), .A1(n5525) );
  inv01 U2700 ( .Y(n5534), .A(n5547) );
  nand02 U2701 ( .Y(n5548), .A0(n5523), .A1(n5526) );
  inv01 U2702 ( .Y(n5536), .A(n5548) );
  nand02 U2703 ( .Y(n5549), .A0(n5524), .A1(n5525) );
  inv01 U2704 ( .Y(n5538), .A(n5549) );
  nand02 U2705 ( .Y(n5550), .A0(n5524), .A1(n5526) );
  inv01 U2706 ( .Y(n5540), .A(n5550) );
  nand02 U2707 ( .Y(n5551), .A0(n5525), .A1(n5527) );
  inv01 U2708 ( .Y(n5542), .A(n5551) );
  nand02 U2709 ( .Y(n5552), .A0(n5526), .A1(n5527) );
  inv01 U2710 ( .Y(n5544), .A(n5552) );
  nand02 U2711 ( .Y(n5553), .A0(n5529), .A1(n5531) );
  inv01 U2712 ( .Y(n5554), .A(n5553) );
  nand02 U2713 ( .Y(n5555), .A0(n5533), .A1(n5535) );
  inv01 U2714 ( .Y(n5556), .A(n5555) );
  nand02 U2715 ( .Y(n5557), .A0(n5554), .A1(n5556) );
  inv01 U2716 ( .Y(n5521), .A(n5557) );
  nand02 U2717 ( .Y(n5558), .A0(n5537), .A1(n5539) );
  inv01 U2718 ( .Y(n5559), .A(n5558) );
  nand02 U2719 ( .Y(n5560), .A0(n5541), .A1(n5543) );
  inv01 U2720 ( .Y(n5561), .A(n5560) );
  nand02 U2721 ( .Y(n5562), .A0(n5559), .A1(n5561) );
  inv01 U2722 ( .Y(n5522), .A(n5562) );
  nand02 U2723 ( .Y(n7925), .A0(n5563), .A1(n5564) );
  inv02 U2724 ( .Y(n5565), .A(n7935) );
  inv02 U2725 ( .Y(n5566), .A(n7934) );
  inv02 U2726 ( .Y(n5567), .A(n7831) );
  inv02 U2727 ( .Y(n5568), .A(n7675) );
  inv02 U2728 ( .Y(n5569), .A(n7668) );
  nand02 U2729 ( .Y(n5570), .A0(n5567), .A1(n5571) );
  nand02 U2730 ( .Y(n5572), .A0(n5568), .A1(n5573) );
  nand02 U2731 ( .Y(n5574), .A0(n5569), .A1(n5575) );
  nand02 U2732 ( .Y(n5576), .A0(n5569), .A1(n5577) );
  nand02 U2733 ( .Y(n5578), .A0(n5873), .A1(n5579) );
  nand02 U2734 ( .Y(n5580), .A0(n5873), .A1(n5581) );
  nand02 U2735 ( .Y(n5582), .A0(n5873), .A1(n5583) );
  nand02 U2736 ( .Y(n5584), .A0(n5873), .A1(n5585) );
  nand02 U2737 ( .Y(n5586), .A0(n5565), .A1(n5566) );
  inv01 U2738 ( .Y(n5571), .A(n5586) );
  nand02 U2739 ( .Y(n5587), .A0(n5565), .A1(n5566) );
  inv01 U2740 ( .Y(n5573), .A(n5587) );
  nand02 U2741 ( .Y(n5588), .A0(n5565), .A1(n5567) );
  inv01 U2742 ( .Y(n5575), .A(n5588) );
  nand02 U2743 ( .Y(n5589), .A0(n5565), .A1(n5568) );
  inv01 U2744 ( .Y(n5577), .A(n5589) );
  nand02 U2745 ( .Y(n5590), .A0(n5566), .A1(n5567) );
  inv01 U2746 ( .Y(n5579), .A(n5590) );
  nand02 U2747 ( .Y(n5591), .A0(n5566), .A1(n5568) );
  inv01 U2748 ( .Y(n5581), .A(n5591) );
  nand02 U2749 ( .Y(n5592), .A0(n5567), .A1(n5569) );
  inv01 U2750 ( .Y(n5583), .A(n5592) );
  nand02 U2751 ( .Y(n5593), .A0(n5568), .A1(n5569) );
  inv01 U2752 ( .Y(n5585), .A(n5593) );
  nand02 U2753 ( .Y(n5594), .A0(n5570), .A1(n5572) );
  inv01 U2754 ( .Y(n5595), .A(n5594) );
  nand02 U2755 ( .Y(n5596), .A0(n5574), .A1(n5576) );
  inv01 U2756 ( .Y(n5597), .A(n5596) );
  nand02 U2757 ( .Y(n5598), .A0(n5595), .A1(n5597) );
  inv01 U2758 ( .Y(n5563), .A(n5598) );
  nand02 U2759 ( .Y(n5599), .A0(n5578), .A1(n5580) );
  inv01 U2760 ( .Y(n5600), .A(n5599) );
  nand02 U2761 ( .Y(n5601), .A0(n5582), .A1(n5584) );
  inv01 U2762 ( .Y(n5602), .A(n5601) );
  nand02 U2763 ( .Y(n5603), .A0(n5600), .A1(n5602) );
  inv01 U2764 ( .Y(n5564), .A(n5603) );
  nand02 U2765 ( .Y(n7959), .A0(n5604), .A1(n5605) );
  inv02 U2766 ( .Y(n5606), .A(n7842) );
  inv02 U2767 ( .Y(n5607), .A(n7892) );
  inv02 U2768 ( .Y(n5609), .A(n7668) );
  inv02 U2769 ( .Y(n5610), .A(n7676) );
  nand02 U2770 ( .Y(n5611), .A0(n5608), .A1(n5612) );
  nand02 U2771 ( .Y(n5613), .A0(n5609), .A1(n5614) );
  nand02 U2772 ( .Y(n5615), .A0(n5610), .A1(n5616) );
  nand02 U2773 ( .Y(n5617), .A0(n5610), .A1(n5618) );
  nand02 U2774 ( .Y(n5619), .A0(n5873), .A1(n5620) );
  nand02 U2775 ( .Y(n5621), .A0(n5873), .A1(n5622) );
  nand02 U2776 ( .Y(n5623), .A0(n5873), .A1(n5624) );
  nand02 U2777 ( .Y(n5625), .A0(n5873), .A1(n5626) );
  nand02 U2778 ( .Y(n5627), .A0(n5606), .A1(n5607) );
  inv01 U2779 ( .Y(n5612), .A(n5627) );
  nand02 U2780 ( .Y(n5628), .A0(n5606), .A1(n5607) );
  inv01 U2781 ( .Y(n5614), .A(n5628) );
  nand02 U2782 ( .Y(n5629), .A0(n5606), .A1(n5608) );
  inv01 U2783 ( .Y(n5616), .A(n5629) );
  nand02 U2784 ( .Y(n5630), .A0(n5606), .A1(n5609) );
  inv01 U2785 ( .Y(n5618), .A(n5630) );
  nand02 U2786 ( .Y(n5631), .A0(n5607), .A1(n5608) );
  inv01 U2787 ( .Y(n5620), .A(n5631) );
  nand02 U2788 ( .Y(n5632), .A0(n5607), .A1(n5609) );
  inv01 U2789 ( .Y(n5622), .A(n5632) );
  nand02 U2790 ( .Y(n5633), .A0(n5608), .A1(n5610) );
  inv01 U2791 ( .Y(n5624), .A(n5633) );
  nand02 U2792 ( .Y(n5634), .A0(n5609), .A1(n5610) );
  inv01 U2793 ( .Y(n5626), .A(n5634) );
  nand02 U2794 ( .Y(n5635), .A0(n5611), .A1(n5613) );
  inv01 U2795 ( .Y(n5636), .A(n5635) );
  nand02 U2796 ( .Y(n5637), .A0(n5615), .A1(n5617) );
  inv01 U2797 ( .Y(n5638), .A(n5637) );
  nand02 U2798 ( .Y(n5639), .A0(n5636), .A1(n5638) );
  inv01 U2799 ( .Y(n5604), .A(n5639) );
  nand02 U2800 ( .Y(n5640), .A0(n5619), .A1(n5621) );
  inv01 U2801 ( .Y(n5641), .A(n5640) );
  nand02 U2802 ( .Y(n5642), .A0(n5623), .A1(n5625) );
  inv01 U2803 ( .Y(n5643), .A(n5642) );
  nand02 U2804 ( .Y(n5644), .A0(n5641), .A1(n5643) );
  inv01 U2805 ( .Y(n5605), .A(n5644) );
  nand02 U2806 ( .Y(n7969), .A0(n5645), .A1(n5646) );
  inv02 U2807 ( .Y(n5647), .A(n7920) );
  inv02 U2808 ( .Y(n5648), .A(n7862) );
  inv02 U2809 ( .Y(n5649), .A(n7924) );
  inv02 U2810 ( .Y(n5650), .A(n7676) );
  inv02 U2811 ( .Y(n5651), .A(n7668) );
  nand02 U2812 ( .Y(n5652), .A0(n5649), .A1(n5653) );
  nand02 U2813 ( .Y(n5654), .A0(n5650), .A1(n5655) );
  nand02 U2814 ( .Y(n5656), .A0(n5873), .A1(n5657) );
  nand02 U2815 ( .Y(n5658), .A0(n5873), .A1(n5659) );
  nand02 U2816 ( .Y(n5660), .A0(n5651), .A1(n5661) );
  nand02 U2817 ( .Y(n5662), .A0(n5651), .A1(n5663) );
  nand02 U2818 ( .Y(n5664), .A0(n5651), .A1(n5665) );
  nand02 U2819 ( .Y(n5666), .A0(n5651), .A1(n5667) );
  nand02 U2820 ( .Y(n5668), .A0(n5647), .A1(n5648) );
  inv01 U2821 ( .Y(n5653), .A(n5668) );
  nand02 U2822 ( .Y(n5669), .A0(n5647), .A1(n5648) );
  inv01 U2823 ( .Y(n5655), .A(n5669) );
  nand02 U2824 ( .Y(n5670), .A0(n5647), .A1(n5649) );
  inv01 U2825 ( .Y(n5657), .A(n5670) );
  nand02 U2826 ( .Y(n5671), .A0(n5647), .A1(n5650) );
  inv01 U2827 ( .Y(n5659), .A(n5671) );
  nand02 U2828 ( .Y(n5672), .A0(n5648), .A1(n5649) );
  inv01 U2829 ( .Y(n5661), .A(n5672) );
  nand02 U2830 ( .Y(n5673), .A0(n5648), .A1(n5650) );
  inv01 U2831 ( .Y(n5663), .A(n5673) );
  nand02 U2832 ( .Y(n5674), .A0(n5649), .A1(n5873) );
  inv01 U2833 ( .Y(n5665), .A(n5674) );
  nand02 U2834 ( .Y(n5675), .A0(n5650), .A1(n5873) );
  inv01 U2835 ( .Y(n5667), .A(n5675) );
  nand02 U2836 ( .Y(n5676), .A0(n5652), .A1(n5654) );
  inv01 U2837 ( .Y(n5677), .A(n5676) );
  nand02 U2838 ( .Y(n5678), .A0(n5656), .A1(n5658) );
  inv01 U2839 ( .Y(n5679), .A(n5678) );
  nand02 U2840 ( .Y(n5680), .A0(n5677), .A1(n5679) );
  inv01 U2841 ( .Y(n5645), .A(n5680) );
  nand02 U2842 ( .Y(n5681), .A0(n5660), .A1(n5662) );
  inv01 U2843 ( .Y(n5682), .A(n5681) );
  nand02 U2844 ( .Y(n5683), .A0(n5664), .A1(n5666) );
  inv01 U2845 ( .Y(n5684), .A(n5683) );
  nand02 U2846 ( .Y(n5685), .A0(n5682), .A1(n5684) );
  inv01 U2847 ( .Y(n5646), .A(n5685) );
  inv02 U2848 ( .Y(n7924), .A(n7471) );
  inv01 U2849 ( .Y(n7761), .A(n5686) );
  inv01 U2850 ( .Y(n5687), .A(opa_i[20]) );
  inv01 U2851 ( .Y(n5688), .A(opa_i[21]) );
  inv01 U2852 ( .Y(n5689), .A(opa_i[1]) );
  nand02 U2853 ( .Y(n5686), .A0(n5689), .A1(n5690) );
  nand02 U2854 ( .Y(n5691), .A0(n5687), .A1(n5688) );
  inv01 U2855 ( .Y(n5690), .A(n5691) );
  nand02 U2856 ( .Y(n7815), .A0(n5692), .A1(n5693) );
  inv02 U2857 ( .Y(n5694), .A(n7827) );
  inv02 U2858 ( .Y(n5695), .A(n7825) );
  inv02 U2859 ( .Y(n5696), .A(n7823) );
  inv02 U2860 ( .Y(n5697), .A(n7677) );
  inv02 U2861 ( .Y(n5698), .A(n7671) );
  inv02 U2862 ( .Y(n5699), .A(n7670) );
  nand02 U2863 ( .Y(n5700), .A0(n5696), .A1(n5701) );
  nand02 U2864 ( .Y(n5702), .A0(n5697), .A1(n5703) );
  nand02 U2865 ( .Y(n5704), .A0(n5698), .A1(n5705) );
  nand02 U2866 ( .Y(n5706), .A0(n5698), .A1(n5707) );
  nand02 U2867 ( .Y(n5708), .A0(n5699), .A1(n5709) );
  nand02 U2868 ( .Y(n5710), .A0(n5699), .A1(n5711) );
  nand02 U2869 ( .Y(n5712), .A0(n5699), .A1(n5713) );
  nand02 U2870 ( .Y(n5714), .A0(n5699), .A1(n5715) );
  nand02 U2871 ( .Y(n5716), .A0(n5694), .A1(n5695) );
  inv01 U2872 ( .Y(n5701), .A(n5716) );
  nand02 U2873 ( .Y(n5717), .A0(n5694), .A1(n5695) );
  inv01 U2874 ( .Y(n5703), .A(n5717) );
  nand02 U2875 ( .Y(n5718), .A0(n5694), .A1(n5696) );
  inv01 U2876 ( .Y(n5705), .A(n5718) );
  nand02 U2877 ( .Y(n5719), .A0(n5694), .A1(n5697) );
  inv01 U2878 ( .Y(n5707), .A(n5719) );
  nand02 U2879 ( .Y(n5720), .A0(n5695), .A1(n5696) );
  inv01 U2880 ( .Y(n5709), .A(n5720) );
  nand02 U2881 ( .Y(n5721), .A0(n5695), .A1(n5697) );
  inv01 U2882 ( .Y(n5711), .A(n5721) );
  nand02 U2883 ( .Y(n5722), .A0(n5696), .A1(n5698) );
  inv01 U2884 ( .Y(n5713), .A(n5722) );
  nand02 U2885 ( .Y(n5723), .A0(n5697), .A1(n5698) );
  inv01 U2886 ( .Y(n5715), .A(n5723) );
  nand02 U2887 ( .Y(n5724), .A0(n5700), .A1(n5702) );
  inv01 U2888 ( .Y(n5725), .A(n5724) );
  nand02 U2889 ( .Y(n5726), .A0(n5704), .A1(n5706) );
  inv01 U2890 ( .Y(n5727), .A(n5726) );
  nand02 U2891 ( .Y(n5728), .A0(n5725), .A1(n5727) );
  inv01 U2892 ( .Y(n5692), .A(n5728) );
  nand02 U2893 ( .Y(n5729), .A0(n5708), .A1(n5710) );
  inv01 U2894 ( .Y(n5730), .A(n5729) );
  nand02 U2895 ( .Y(n5731), .A0(n5712), .A1(n5714) );
  inv01 U2896 ( .Y(n5732), .A(n5731) );
  nand02 U2897 ( .Y(n5733), .A0(n5730), .A1(n5732) );
  inv01 U2898 ( .Y(n5693), .A(n5733) );
  nand02 U2899 ( .Y(n7996), .A0(n5734), .A1(n5735) );
  inv02 U2900 ( .Y(n5736), .A(n7595) );
  inv02 U2901 ( .Y(n5737), .A(n7586) );
  inv02 U2902 ( .Y(n5738), .A(n7640) );
  inv02 U2903 ( .Y(n5739), .A(n7848) );
  inv02 U2904 ( .Y(n5740), .A(n7842) );
  nand02 U2905 ( .Y(n5741), .A0(n5738), .A1(n5742) );
  nand02 U2906 ( .Y(n5743), .A0(n5608), .A1(n5744) );
  nand02 U2907 ( .Y(n5745), .A0(n5739), .A1(n5746) );
  nand02 U2908 ( .Y(n5747), .A0(n5739), .A1(n5748) );
  nand02 U2909 ( .Y(n5749), .A0(n5740), .A1(n5750) );
  nand02 U2910 ( .Y(n5751), .A0(n5740), .A1(n5752) );
  nand02 U2911 ( .Y(n5753), .A0(n5740), .A1(n5754) );
  nand02 U2912 ( .Y(n5755), .A0(n5740), .A1(n5756) );
  nand02 U2913 ( .Y(n5757), .A0(n5736), .A1(n5737) );
  inv01 U2914 ( .Y(n5742), .A(n5757) );
  nand02 U2915 ( .Y(n5758), .A0(n5736), .A1(n5737) );
  inv01 U2916 ( .Y(n5744), .A(n5758) );
  nand02 U2917 ( .Y(n5759), .A0(n5736), .A1(n5738) );
  inv01 U2918 ( .Y(n5746), .A(n5759) );
  nand02 U2919 ( .Y(n5760), .A0(n5736), .A1(n5608) );
  inv01 U2920 ( .Y(n5748), .A(n5760) );
  nand02 U2921 ( .Y(n5761), .A0(n5737), .A1(n5738) );
  inv01 U2922 ( .Y(n5750), .A(n5761) );
  nand02 U2923 ( .Y(n5762), .A0(n5737), .A1(n5608) );
  inv01 U2924 ( .Y(n5752), .A(n5762) );
  nand02 U2925 ( .Y(n5763), .A0(n5738), .A1(n5739) );
  inv01 U2926 ( .Y(n5754), .A(n5763) );
  nand02 U2927 ( .Y(n5764), .A0(n5608), .A1(n5739) );
  inv01 U2928 ( .Y(n5756), .A(n5764) );
  nand02 U2929 ( .Y(n5765), .A0(n5741), .A1(n5743) );
  inv01 U2930 ( .Y(n5766), .A(n5765) );
  nand02 U2931 ( .Y(n5767), .A0(n5745), .A1(n5747) );
  inv01 U2932 ( .Y(n5768), .A(n5767) );
  nand02 U2933 ( .Y(n5769), .A0(n5766), .A1(n5768) );
  inv01 U2934 ( .Y(n5734), .A(n5769) );
  nand02 U2935 ( .Y(n5770), .A0(n5749), .A1(n5751) );
  inv01 U2936 ( .Y(n5771), .A(n5770) );
  nand02 U2937 ( .Y(n5772), .A0(n5753), .A1(n5755) );
  inv01 U2938 ( .Y(n5773), .A(n5772) );
  nand02 U2939 ( .Y(n5774), .A0(n5771), .A1(n5773) );
  inv01 U2940 ( .Y(n5735), .A(n5774) );
  nand02 U2941 ( .Y(n7731), .A0(n5775), .A1(n7413) );
  inv01 U2942 ( .Y(n5776), .A(n7757) );
  inv01 U2943 ( .Y(n5777), .A(n7756) );
  nand02 U2944 ( .Y(n5775), .A0(n5776), .A1(n5777) );
  inv01 U2945 ( .Y(n7763), .A(n5778) );
  inv01 U2946 ( .Y(n5779), .A(opa_i[5]) );
  inv01 U2947 ( .Y(n5780), .A(opa_i[6]) );
  inv01 U2948 ( .Y(n5781), .A(opa_i[4]) );
  nand02 U2949 ( .Y(n5778), .A0(n5781), .A1(n5782) );
  nand02 U2950 ( .Y(n5783), .A0(n5779), .A1(n5780) );
  inv01 U2951 ( .Y(n5782), .A(n5783) );
  nand02 U2952 ( .Y(n7966), .A0(n5784), .A1(n5785) );
  inv02 U2953 ( .Y(n5786), .A(n7908) );
  inv02 U2954 ( .Y(n5787), .A(n7854) );
  inv02 U2955 ( .Y(n5788), .A(n7885) );
  inv02 U2956 ( .Y(n5789), .A(n7655) );
  inv02 U2957 ( .Y(n5790), .A(n7615) );
  inv02 U2958 ( .Y(n5791), .A(n7678) );
  nand02 U2959 ( .Y(n5792), .A0(n5788), .A1(n5793) );
  nand02 U2960 ( .Y(n5794), .A0(n5789), .A1(n5795) );
  nand02 U2961 ( .Y(n5796), .A0(n5790), .A1(n5797) );
  nand02 U2962 ( .Y(n5798), .A0(n5790), .A1(n5799) );
  nand02 U2963 ( .Y(n5800), .A0(n5791), .A1(n5801) );
  nand02 U2964 ( .Y(n5802), .A0(n5791), .A1(n5803) );
  nand02 U2965 ( .Y(n5804), .A0(n5791), .A1(n5805) );
  nand02 U2966 ( .Y(n5806), .A0(n5791), .A1(n5807) );
  nand02 U2967 ( .Y(n5808), .A0(n5786), .A1(n5787) );
  inv01 U2968 ( .Y(n5793), .A(n5808) );
  nand02 U2969 ( .Y(n5809), .A0(n5786), .A1(n5787) );
  inv01 U2970 ( .Y(n5795), .A(n5809) );
  nand02 U2971 ( .Y(n5810), .A0(n5786), .A1(n5788) );
  inv01 U2972 ( .Y(n5797), .A(n5810) );
  nand02 U2973 ( .Y(n5811), .A0(n5786), .A1(n5789) );
  inv01 U2974 ( .Y(n5799), .A(n5811) );
  nand02 U2975 ( .Y(n5812), .A0(n5787), .A1(n5788) );
  inv01 U2976 ( .Y(n5801), .A(n5812) );
  nand02 U2977 ( .Y(n5813), .A0(n5787), .A1(n5789) );
  inv01 U2978 ( .Y(n5803), .A(n5813) );
  nand02 U2979 ( .Y(n5814), .A0(n5788), .A1(n5790) );
  inv01 U2980 ( .Y(n5805), .A(n5814) );
  nand02 U2981 ( .Y(n5815), .A0(n5789), .A1(n5790) );
  inv01 U2982 ( .Y(n5807), .A(n5815) );
  nand02 U2983 ( .Y(n5816), .A0(n5792), .A1(n5794) );
  inv01 U2984 ( .Y(n5817), .A(n5816) );
  nand02 U2985 ( .Y(n5818), .A0(n5796), .A1(n5798) );
  inv01 U2986 ( .Y(n5819), .A(n5818) );
  nand02 U2987 ( .Y(n5820), .A0(n5817), .A1(n5819) );
  inv01 U2988 ( .Y(n5784), .A(n5820) );
  nand02 U2989 ( .Y(n5821), .A0(n5800), .A1(n5802) );
  inv01 U2990 ( .Y(n5822), .A(n5821) );
  nand02 U2991 ( .Y(n5823), .A0(n5804), .A1(n5806) );
  inv01 U2992 ( .Y(n5824), .A(n5823) );
  nand02 U2993 ( .Y(n5825), .A0(n5822), .A1(n5824) );
  inv01 U2994 ( .Y(n5785), .A(n5825) );
  nand02 U2995 ( .Y(n7952), .A0(n5826), .A1(n5827) );
  inv02 U2996 ( .Y(n5828), .A(n7860) );
  inv02 U2997 ( .Y(n5829), .A(n7953) );
  inv02 U2998 ( .Y(n5830), .A(n7818) );
  inv02 U2999 ( .Y(n5831), .A(n7670) );
  inv02 U3000 ( .Y(n5832), .A(n7283) );
  inv02 U3001 ( .Y(n5833), .A(n7677) );
  nand02 U3002 ( .Y(n5834), .A0(n5830), .A1(n5835) );
  nand02 U3003 ( .Y(n5836), .A0(n5831), .A1(n5837) );
  nand02 U3004 ( .Y(n5838), .A0(n5832), .A1(n5839) );
  nand02 U3005 ( .Y(n5840), .A0(n5832), .A1(n5841) );
  nand02 U3006 ( .Y(n5842), .A0(n5833), .A1(n5843) );
  nand02 U3007 ( .Y(n5844), .A0(n5833), .A1(n5845) );
  nand02 U3008 ( .Y(n5846), .A0(n5833), .A1(n5847) );
  nand02 U3009 ( .Y(n5848), .A0(n5833), .A1(n5849) );
  nand02 U3010 ( .Y(n5850), .A0(n5828), .A1(n5829) );
  inv01 U3011 ( .Y(n5835), .A(n5850) );
  nand02 U3012 ( .Y(n5851), .A0(n5828), .A1(n5829) );
  inv01 U3013 ( .Y(n5837), .A(n5851) );
  nand02 U3014 ( .Y(n5852), .A0(n5828), .A1(n5830) );
  inv01 U3015 ( .Y(n5839), .A(n5852) );
  nand02 U3016 ( .Y(n5853), .A0(n5828), .A1(n5831) );
  inv01 U3017 ( .Y(n5841), .A(n5853) );
  nand02 U3018 ( .Y(n5854), .A0(n5829), .A1(n5830) );
  inv01 U3019 ( .Y(n5843), .A(n5854) );
  nand02 U3020 ( .Y(n5855), .A0(n5829), .A1(n5831) );
  inv01 U3021 ( .Y(n5845), .A(n5855) );
  nand02 U3022 ( .Y(n5856), .A0(n5830), .A1(n5832) );
  inv01 U3023 ( .Y(n5847), .A(n5856) );
  nand02 U3024 ( .Y(n5857), .A0(n5831), .A1(n5832) );
  inv01 U3025 ( .Y(n5849), .A(n5857) );
  nand02 U3026 ( .Y(n5858), .A0(n5834), .A1(n5836) );
  inv01 U3027 ( .Y(n5859), .A(n5858) );
  nand02 U3028 ( .Y(n5860), .A0(n5838), .A1(n5840) );
  inv01 U3029 ( .Y(n5861), .A(n5860) );
  nand02 U3030 ( .Y(n5862), .A0(n5859), .A1(n5861) );
  inv01 U3031 ( .Y(n5826), .A(n5862) );
  nand02 U3032 ( .Y(n5863), .A0(n5842), .A1(n5844) );
  inv01 U3033 ( .Y(n5864), .A(n5863) );
  nand02 U3034 ( .Y(n5865), .A0(n5846), .A1(n5848) );
  inv01 U3035 ( .Y(n5866), .A(n5865) );
  nand02 U3036 ( .Y(n5867), .A0(n5864), .A1(n5866) );
  inv01 U3037 ( .Y(n5827), .A(n5867) );
  nand02 U3038 ( .Y(n7973), .A0(n5868), .A1(n5869) );
  inv02 U3039 ( .Y(n5870), .A(n7934) );
  inv02 U3040 ( .Y(n5871), .A(n7431) );
  inv02 U3041 ( .Y(n5872), .A(n7930) );
  inv02 U3042 ( .Y(n5874), .A(n7615) );
  inv02 U3043 ( .Y(n5875), .A(n7678) );
  nand02 U3044 ( .Y(n5876), .A0(n5872), .A1(n5877) );
  nand02 U3045 ( .Y(n5878), .A0(n5873), .A1(n5879) );
  nand02 U3046 ( .Y(n5880), .A0(n5874), .A1(n5881) );
  nand02 U3047 ( .Y(n5882), .A0(n5874), .A1(n5883) );
  nand02 U3048 ( .Y(n5884), .A0(n5875), .A1(n5885) );
  nand02 U3049 ( .Y(n5886), .A0(n5875), .A1(n5887) );
  nand02 U3050 ( .Y(n5888), .A0(n5875), .A1(n5889) );
  nand02 U3051 ( .Y(n5890), .A0(n5875), .A1(n5891) );
  nand02 U3052 ( .Y(n5892), .A0(n5870), .A1(n5871) );
  inv01 U3053 ( .Y(n5877), .A(n5892) );
  nand02 U3054 ( .Y(n5893), .A0(n5870), .A1(n5871) );
  inv01 U3055 ( .Y(n5879), .A(n5893) );
  nand02 U3056 ( .Y(n5894), .A0(n5870), .A1(n5872) );
  inv01 U3057 ( .Y(n5881), .A(n5894) );
  nand02 U3058 ( .Y(n5895), .A0(n5870), .A1(n5873) );
  inv01 U3059 ( .Y(n5883), .A(n5895) );
  nand02 U3060 ( .Y(n5896), .A0(n5871), .A1(n5872) );
  inv01 U3061 ( .Y(n5885), .A(n5896) );
  nand02 U3062 ( .Y(n5897), .A0(n5871), .A1(n5873) );
  inv01 U3063 ( .Y(n5887), .A(n5897) );
  nand02 U3064 ( .Y(n5898), .A0(n5872), .A1(n5874) );
  inv01 U3065 ( .Y(n5889), .A(n5898) );
  nand02 U3066 ( .Y(n5899), .A0(n5873), .A1(n5874) );
  inv01 U3067 ( .Y(n5891), .A(n5899) );
  nand02 U3068 ( .Y(n5900), .A0(n5876), .A1(n5878) );
  inv01 U3069 ( .Y(n5901), .A(n5900) );
  nand02 U3070 ( .Y(n5902), .A0(n5880), .A1(n5882) );
  inv01 U3071 ( .Y(n5903), .A(n5902) );
  nand02 U3072 ( .Y(n5904), .A0(n5901), .A1(n5903) );
  inv01 U3073 ( .Y(n5868), .A(n5904) );
  nand02 U3074 ( .Y(n5905), .A0(n5884), .A1(n5886) );
  inv01 U3075 ( .Y(n5906), .A(n5905) );
  nand02 U3076 ( .Y(n5907), .A0(n5888), .A1(n5890) );
  inv01 U3077 ( .Y(n5908), .A(n5907) );
  nand02 U3078 ( .Y(n5909), .A0(n5906), .A1(n5908) );
  inv01 U3079 ( .Y(n5869), .A(n5909) );
  inv04 U3080 ( .Y(n7615), .A(n7614) );
  nand02 U3081 ( .Y(n7829), .A0(n5910), .A1(n5911) );
  inv02 U3082 ( .Y(n5912), .A(n7832) );
  inv02 U3083 ( .Y(n5913), .A(n7831) );
  inv02 U3084 ( .Y(n5914), .A(n7830) );
  inv02 U3085 ( .Y(n5915), .A(n7675) );
  inv02 U3086 ( .Y(n5916), .A(n7623) );
  inv02 U3087 ( .Y(n5917), .A(n7660) );
  nand02 U3088 ( .Y(n5918), .A0(n5914), .A1(n5919) );
  nand02 U3089 ( .Y(n5920), .A0(n5915), .A1(n5921) );
  nand02 U3090 ( .Y(n5922), .A0(n5916), .A1(n5923) );
  nand02 U3091 ( .Y(n5924), .A0(n5916), .A1(n5925) );
  nand02 U3092 ( .Y(n5926), .A0(n5917), .A1(n5927) );
  nand02 U3093 ( .Y(n5928), .A0(n5917), .A1(n5929) );
  nand02 U3094 ( .Y(n5930), .A0(n5917), .A1(n5931) );
  nand02 U3095 ( .Y(n5932), .A0(n5917), .A1(n5933) );
  nand02 U3096 ( .Y(n5934), .A0(n5912), .A1(n5913) );
  inv01 U3097 ( .Y(n5919), .A(n5934) );
  nand02 U3098 ( .Y(n5935), .A0(n5912), .A1(n5913) );
  inv01 U3099 ( .Y(n5921), .A(n5935) );
  nand02 U3100 ( .Y(n5936), .A0(n5912), .A1(n5914) );
  inv01 U3101 ( .Y(n5923), .A(n5936) );
  nand02 U3102 ( .Y(n5937), .A0(n5912), .A1(n5915) );
  inv01 U3103 ( .Y(n5925), .A(n5937) );
  nand02 U3104 ( .Y(n5938), .A0(n5913), .A1(n5914) );
  inv01 U3105 ( .Y(n5927), .A(n5938) );
  nand02 U3106 ( .Y(n5939), .A0(n5913), .A1(n5915) );
  inv01 U3107 ( .Y(n5929), .A(n5939) );
  nand02 U3108 ( .Y(n5940), .A0(n5914), .A1(n5916) );
  inv01 U3109 ( .Y(n5931), .A(n5940) );
  nand02 U3110 ( .Y(n5941), .A0(n5915), .A1(n5916) );
  inv01 U3111 ( .Y(n5933), .A(n5941) );
  nand02 U3112 ( .Y(n5942), .A0(n5918), .A1(n5920) );
  inv01 U3113 ( .Y(n5943), .A(n5942) );
  nand02 U3114 ( .Y(n5944), .A0(n5922), .A1(n5924) );
  inv01 U3115 ( .Y(n5945), .A(n5944) );
  nand02 U3116 ( .Y(n5946), .A0(n5943), .A1(n5945) );
  inv01 U3117 ( .Y(n5910), .A(n5946) );
  nand02 U3118 ( .Y(n5947), .A0(n5926), .A1(n5928) );
  inv01 U3119 ( .Y(n5948), .A(n5947) );
  nand02 U3120 ( .Y(n5949), .A0(n5930), .A1(n5932) );
  inv01 U3121 ( .Y(n5950), .A(n5949) );
  nand02 U3122 ( .Y(n5951), .A0(n5948), .A1(n5950) );
  inv01 U3123 ( .Y(n5911), .A(n5951) );
  or04 U3124 ( .Y(n5952), .A0(s_fracto28_1[2]), .A1(s_fracto28_1[1]), .A2(
        s_fracto28_1[0]), .A3(n7807) );
  inv01 U3125 ( .Y(n5953), .A(n5952) );
  nand02 U3126 ( .Y(n7816), .A0(n5954), .A1(n5955) );
  inv02 U3127 ( .Y(n5956), .A(n7821) );
  inv02 U3128 ( .Y(n5957), .A(n7819) );
  inv02 U3129 ( .Y(n5958), .A(n7818) );
  inv02 U3130 ( .Y(n5959), .A(n7675) );
  inv02 U3131 ( .Y(n5960), .A(n7623) );
  inv02 U3132 ( .Y(n5961), .A(n7657) );
  nand02 U3133 ( .Y(n5962), .A0(n5958), .A1(n5963) );
  nand02 U3134 ( .Y(n5964), .A0(n5959), .A1(n5965) );
  nand02 U3135 ( .Y(n5966), .A0(n5960), .A1(n5967) );
  nand02 U3136 ( .Y(n5968), .A0(n5960), .A1(n5969) );
  nand02 U3137 ( .Y(n5970), .A0(n5961), .A1(n5971) );
  nand02 U3138 ( .Y(n5972), .A0(n5961), .A1(n5973) );
  nand02 U3139 ( .Y(n5974), .A0(n5961), .A1(n5975) );
  nand02 U3140 ( .Y(n5976), .A0(n5961), .A1(n5977) );
  nand02 U3141 ( .Y(n5978), .A0(n5956), .A1(n5957) );
  inv01 U3142 ( .Y(n5963), .A(n5978) );
  nand02 U3143 ( .Y(n5979), .A0(n5956), .A1(n5957) );
  inv01 U3144 ( .Y(n5965), .A(n5979) );
  nand02 U3145 ( .Y(n5980), .A0(n5956), .A1(n5958) );
  inv01 U3146 ( .Y(n5967), .A(n5980) );
  nand02 U3147 ( .Y(n5981), .A0(n5956), .A1(n5959) );
  inv01 U3148 ( .Y(n5969), .A(n5981) );
  nand02 U3149 ( .Y(n5982), .A0(n5957), .A1(n5958) );
  inv01 U3150 ( .Y(n5971), .A(n5982) );
  nand02 U3151 ( .Y(n5983), .A0(n5957), .A1(n5959) );
  inv01 U3152 ( .Y(n5973), .A(n5983) );
  nand02 U3153 ( .Y(n5984), .A0(n5958), .A1(n5960) );
  inv01 U3154 ( .Y(n5975), .A(n5984) );
  nand02 U3155 ( .Y(n5985), .A0(n5959), .A1(n5960) );
  inv01 U3156 ( .Y(n5977), .A(n5985) );
  nand02 U3157 ( .Y(n5986), .A0(n5962), .A1(n5964) );
  inv01 U3158 ( .Y(n5987), .A(n5986) );
  nand02 U3159 ( .Y(n5988), .A0(n5966), .A1(n5968) );
  inv01 U3160 ( .Y(n5989), .A(n5988) );
  nand02 U3161 ( .Y(n5990), .A0(n5987), .A1(n5989) );
  inv01 U3162 ( .Y(n5954), .A(n5990) );
  nand02 U3163 ( .Y(n5991), .A0(n5970), .A1(n5972) );
  inv01 U3164 ( .Y(n5992), .A(n5991) );
  nand02 U3165 ( .Y(n5993), .A0(n5974), .A1(n5976) );
  inv01 U3166 ( .Y(n5994), .A(n5993) );
  nand02 U3167 ( .Y(n5995), .A0(n5992), .A1(n5994) );
  inv01 U3168 ( .Y(n5955), .A(n5995) );
  inv04 U3169 ( .Y(n7623), .A(n7622) );
  nand02 U3170 ( .Y(n7998), .A0(n5996), .A1(n5997) );
  inv02 U3171 ( .Y(n5998), .A(n7855) );
  inv02 U3172 ( .Y(n5999), .A(n7602) );
  inv02 U3173 ( .Y(n6000), .A(n7856) );
  inv02 U3174 ( .Y(n6001), .A(n7677) );
  inv02 U3175 ( .Y(n6002), .A(n7623) );
  inv02 U3176 ( .Y(n6003), .A(n7675) );
  nand02 U3177 ( .Y(n6004), .A0(n6000), .A1(n6005) );
  nand02 U3178 ( .Y(n6006), .A0(n6001), .A1(n6007) );
  nand02 U3179 ( .Y(n6008), .A0(n6002), .A1(n6009) );
  nand02 U3180 ( .Y(n6010), .A0(n6002), .A1(n6011) );
  nand02 U3181 ( .Y(n6012), .A0(n6003), .A1(n6013) );
  nand02 U3182 ( .Y(n6014), .A0(n6003), .A1(n6015) );
  nand02 U3183 ( .Y(n6016), .A0(n6003), .A1(n6017) );
  nand02 U3184 ( .Y(n6018), .A0(n6003), .A1(n6019) );
  nand02 U3185 ( .Y(n6020), .A0(n5998), .A1(n5999) );
  inv01 U3186 ( .Y(n6005), .A(n6020) );
  nand02 U3187 ( .Y(n6021), .A0(n5998), .A1(n5999) );
  inv01 U3188 ( .Y(n6007), .A(n6021) );
  nand02 U3189 ( .Y(n6022), .A0(n5998), .A1(n6000) );
  inv01 U3190 ( .Y(n6009), .A(n6022) );
  nand02 U3191 ( .Y(n6023), .A0(n5998), .A1(n6001) );
  inv01 U3192 ( .Y(n6011), .A(n6023) );
  nand02 U3193 ( .Y(n6024), .A0(n5999), .A1(n6000) );
  inv01 U3194 ( .Y(n6013), .A(n6024) );
  nand02 U3195 ( .Y(n6025), .A0(n5999), .A1(n6001) );
  inv01 U3196 ( .Y(n6015), .A(n6025) );
  nand02 U3197 ( .Y(n6026), .A0(n6000), .A1(n6002) );
  inv01 U3198 ( .Y(n6017), .A(n6026) );
  nand02 U3199 ( .Y(n6027), .A0(n6001), .A1(n6002) );
  inv01 U3200 ( .Y(n6019), .A(n6027) );
  nand02 U3201 ( .Y(n6028), .A0(n6004), .A1(n6006) );
  inv01 U3202 ( .Y(n6029), .A(n6028) );
  nand02 U3203 ( .Y(n6030), .A0(n6008), .A1(n6010) );
  inv01 U3204 ( .Y(n6031), .A(n6030) );
  nand02 U3205 ( .Y(n6032), .A0(n6029), .A1(n6031) );
  inv01 U3206 ( .Y(n5996), .A(n6032) );
  nand02 U3207 ( .Y(n6033), .A0(n6012), .A1(n6014) );
  inv01 U3208 ( .Y(n6034), .A(n6033) );
  nand02 U3209 ( .Y(n6035), .A0(n6016), .A1(n6018) );
  inv01 U3210 ( .Y(n6036), .A(n6035) );
  nand02 U3211 ( .Y(n6037), .A0(n6034), .A1(n6036) );
  inv01 U3212 ( .Y(n5997), .A(n6037) );
  inv01 U3213 ( .Y(n7806), .A(n6038) );
  inv01 U3214 ( .Y(n6039), .A(n7808) );
  inv01 U3215 ( .Y(n6040), .A(n____return2766_0_) );
  inv01 U3216 ( .Y(n6041), .A(n____return2766_1_) );
  inv01 U3217 ( .Y(n6042), .A(n____return2766_2_) );
  nand02 U3218 ( .Y(n6038), .A0(n6043), .A1(n6044) );
  nand02 U3219 ( .Y(n6045), .A0(n6039), .A1(n6040) );
  inv01 U3220 ( .Y(n6043), .A(n6045) );
  nand02 U3221 ( .Y(n6046), .A0(n6041), .A1(n6042) );
  inv01 U3222 ( .Y(n6044), .A(n6046) );
  inv02 U3223 ( .Y(n7856), .A(n7483) );
  nand02 U3224 ( .Y(n7962), .A0(n6047), .A1(n6048) );
  inv02 U3225 ( .Y(n6049), .A(n7649) );
  inv02 U3226 ( .Y(n6050), .A(n7297) );
  inv02 U3227 ( .Y(n6051), .A(n7867) );
  inv02 U3228 ( .Y(n6052), .A(n7963) );
  inv02 U3229 ( .Y(n6053), .A(n7578) );
  inv02 U3230 ( .Y(n6054), .A(n7839) );
  nand02 U3231 ( .Y(n6055), .A0(n6051), .A1(n6056) );
  nand02 U3232 ( .Y(n6057), .A0(n6052), .A1(n6058) );
  nand02 U3233 ( .Y(n6059), .A0(n6053), .A1(n6060) );
  nand02 U3234 ( .Y(n6061), .A0(n6053), .A1(n6062) );
  nand02 U3235 ( .Y(n6063), .A0(n6054), .A1(n6064) );
  nand02 U3236 ( .Y(n6065), .A0(n6054), .A1(n6066) );
  nand02 U3237 ( .Y(n6067), .A0(n6054), .A1(n6068) );
  nand02 U3238 ( .Y(n6069), .A0(n6054), .A1(n6070) );
  nand02 U3239 ( .Y(n6071), .A0(n6049), .A1(n6050) );
  inv01 U3240 ( .Y(n6056), .A(n6071) );
  nand02 U3241 ( .Y(n6072), .A0(n6049), .A1(n6050) );
  inv01 U3242 ( .Y(n6058), .A(n6072) );
  nand02 U3243 ( .Y(n6073), .A0(n6049), .A1(n6051) );
  inv01 U3244 ( .Y(n6060), .A(n6073) );
  nand02 U3245 ( .Y(n6074), .A0(n6049), .A1(n6052) );
  inv01 U3246 ( .Y(n6062), .A(n6074) );
  nand02 U3247 ( .Y(n6075), .A0(n6050), .A1(n6051) );
  inv01 U3248 ( .Y(n6064), .A(n6075) );
  nand02 U3249 ( .Y(n6076), .A0(n6050), .A1(n6052) );
  inv01 U3250 ( .Y(n6066), .A(n6076) );
  nand02 U3251 ( .Y(n6077), .A0(n6051), .A1(n6053) );
  inv01 U3252 ( .Y(n6068), .A(n6077) );
  nand02 U3253 ( .Y(n6078), .A0(n6052), .A1(n6053) );
  inv01 U3254 ( .Y(n6070), .A(n6078) );
  nand02 U3255 ( .Y(n6079), .A0(n6055), .A1(n6057) );
  inv01 U3256 ( .Y(n6080), .A(n6079) );
  nand02 U3257 ( .Y(n6081), .A0(n6059), .A1(n6061) );
  inv01 U3258 ( .Y(n6082), .A(n6081) );
  nand02 U3259 ( .Y(n6083), .A0(n6080), .A1(n6082) );
  inv01 U3260 ( .Y(n6047), .A(n6083) );
  nand02 U3261 ( .Y(n6084), .A0(n6063), .A1(n6065) );
  inv01 U3262 ( .Y(n6085), .A(n6084) );
  nand02 U3263 ( .Y(n6086), .A0(n6067), .A1(n6069) );
  inv01 U3264 ( .Y(n6087), .A(n6086) );
  nand02 U3265 ( .Y(n6088), .A0(n6085), .A1(n6087) );
  inv01 U3266 ( .Y(n6048), .A(n6088) );
  nand02 U3267 ( .Y(n7968), .A0(n6089), .A1(n6090) );
  inv02 U3268 ( .Y(n6091), .A(n7578) );
  inv02 U3269 ( .Y(n6092), .A(n7593) );
  inv02 U3270 ( .Y(n6093), .A(n7649) );
  inv02 U3271 ( .Y(n6094), .A(n7858) );
  inv02 U3272 ( .Y(n6095), .A(n7852) );
  inv02 U3273 ( .Y(n6096), .A(n7603) );
  nand02 U3274 ( .Y(n6097), .A0(n6093), .A1(n6098) );
  nand02 U3275 ( .Y(n6099), .A0(n6094), .A1(n6100) );
  nand02 U3276 ( .Y(n6101), .A0(n6095), .A1(n6102) );
  nand02 U3277 ( .Y(n6103), .A0(n6095), .A1(n6104) );
  nand02 U3278 ( .Y(n6105), .A0(n6096), .A1(n6106) );
  nand02 U3279 ( .Y(n6107), .A0(n6096), .A1(n6108) );
  nand02 U3280 ( .Y(n6109), .A0(n6096), .A1(n6110) );
  nand02 U3281 ( .Y(n6111), .A0(n6096), .A1(n6112) );
  nand02 U3282 ( .Y(n6113), .A0(n6091), .A1(n6092) );
  inv01 U3283 ( .Y(n6098), .A(n6113) );
  nand02 U3284 ( .Y(n6114), .A0(n6091), .A1(n6092) );
  inv01 U3285 ( .Y(n6100), .A(n6114) );
  nand02 U3286 ( .Y(n6115), .A0(n6091), .A1(n6093) );
  inv01 U3287 ( .Y(n6102), .A(n6115) );
  nand02 U3288 ( .Y(n6116), .A0(n6091), .A1(n6094) );
  inv01 U3289 ( .Y(n6104), .A(n6116) );
  nand02 U3290 ( .Y(n6117), .A0(n6092), .A1(n6093) );
  inv01 U3291 ( .Y(n6106), .A(n6117) );
  nand02 U3292 ( .Y(n6118), .A0(n6092), .A1(n6094) );
  inv01 U3293 ( .Y(n6108), .A(n6118) );
  nand02 U3294 ( .Y(n6119), .A0(n6093), .A1(n6095) );
  inv01 U3295 ( .Y(n6110), .A(n6119) );
  nand02 U3296 ( .Y(n6120), .A0(n6094), .A1(n6095) );
  inv01 U3297 ( .Y(n6112), .A(n6120) );
  nand02 U3298 ( .Y(n6121), .A0(n6097), .A1(n6099) );
  inv01 U3299 ( .Y(n6122), .A(n6121) );
  nand02 U3300 ( .Y(n6123), .A0(n6101), .A1(n6103) );
  inv01 U3301 ( .Y(n6124), .A(n6123) );
  nand02 U3302 ( .Y(n6125), .A0(n6122), .A1(n6124) );
  inv01 U3303 ( .Y(n6089), .A(n6125) );
  nand02 U3304 ( .Y(n6126), .A0(n6105), .A1(n6107) );
  inv01 U3305 ( .Y(n6127), .A(n6126) );
  nand02 U3306 ( .Y(n6128), .A0(n6109), .A1(n6111) );
  inv01 U3307 ( .Y(n6129), .A(n6128) );
  nand02 U3308 ( .Y(n6130), .A0(n6127), .A1(n6129) );
  inv01 U3309 ( .Y(n6090), .A(n6130) );
  nand02 U3310 ( .Y(n7993), .A0(n6131), .A1(n6132) );
  inv02 U3311 ( .Y(n6133), .A(n7849) );
  inv02 U3312 ( .Y(n6134), .A(n7623) );
  inv02 U3313 ( .Y(n6135), .A(n7840) );
  inv02 U3314 ( .Y(n6136), .A(n7677) );
  inv02 U3315 ( .Y(n6137), .A(n7297) );
  inv02 U3316 ( .Y(n6138), .A(n7675) );
  nand02 U3317 ( .Y(n6139), .A0(n6135), .A1(n6140) );
  nand02 U3318 ( .Y(n6141), .A0(n6136), .A1(n6142) );
  nand02 U3319 ( .Y(n6143), .A0(n6137), .A1(n6144) );
  nand02 U3320 ( .Y(n6145), .A0(n6137), .A1(n6146) );
  nand02 U3321 ( .Y(n6147), .A0(n6138), .A1(n6148) );
  nand02 U3322 ( .Y(n6149), .A0(n6138), .A1(n6150) );
  nand02 U3323 ( .Y(n6151), .A0(n6138), .A1(n6152) );
  nand02 U3324 ( .Y(n6153), .A0(n6138), .A1(n6154) );
  nand02 U3325 ( .Y(n6155), .A0(n6133), .A1(n6134) );
  inv01 U3326 ( .Y(n6140), .A(n6155) );
  nand02 U3327 ( .Y(n6156), .A0(n6133), .A1(n6134) );
  inv01 U3328 ( .Y(n6142), .A(n6156) );
  nand02 U3329 ( .Y(n6157), .A0(n6133), .A1(n6135) );
  inv01 U3330 ( .Y(n6144), .A(n6157) );
  nand02 U3331 ( .Y(n6158), .A0(n6133), .A1(n6136) );
  inv01 U3332 ( .Y(n6146), .A(n6158) );
  nand02 U3333 ( .Y(n6159), .A0(n6134), .A1(n6135) );
  inv01 U3334 ( .Y(n6148), .A(n6159) );
  nand02 U3335 ( .Y(n6160), .A0(n6134), .A1(n6136) );
  inv01 U3336 ( .Y(n6150), .A(n6160) );
  nand02 U3337 ( .Y(n6161), .A0(n6135), .A1(n6137) );
  inv01 U3338 ( .Y(n6152), .A(n6161) );
  nand02 U3339 ( .Y(n6162), .A0(n6136), .A1(n6137) );
  inv01 U3340 ( .Y(n6154), .A(n6162) );
  nand02 U3341 ( .Y(n6163), .A0(n6139), .A1(n6141) );
  inv01 U3342 ( .Y(n6164), .A(n6163) );
  nand02 U3343 ( .Y(n6165), .A0(n6143), .A1(n6145) );
  inv01 U3344 ( .Y(n6166), .A(n6165) );
  nand02 U3345 ( .Y(n6167), .A0(n6164), .A1(n6166) );
  inv01 U3346 ( .Y(n6131), .A(n6167) );
  nand02 U3347 ( .Y(n6168), .A0(n6147), .A1(n6149) );
  inv01 U3348 ( .Y(n6169), .A(n6168) );
  nand02 U3349 ( .Y(n6170), .A0(n6151), .A1(n6153) );
  inv01 U3350 ( .Y(n6171), .A(n6170) );
  nand02 U3351 ( .Y(n6172), .A0(n6169), .A1(n6171) );
  inv01 U3352 ( .Y(n6132), .A(n6172) );
  nand02 U3353 ( .Y(n8005), .A0(n6173), .A1(n6174) );
  inv02 U3354 ( .Y(n6175), .A(n8006) );
  inv02 U3355 ( .Y(n6176), .A(n7431) );
  inv02 U3356 ( .Y(n6177), .A(n7868) );
  inv02 U3357 ( .Y(n6178), .A(n7677) );
  inv02 U3358 ( .Y(n6179), .A(n7678) );
  inv02 U3359 ( .Y(n6180), .A(n7283) );
  nand02 U3360 ( .Y(n6181), .A0(n6177), .A1(n6182) );
  nand02 U3361 ( .Y(n6183), .A0(n6178), .A1(n6184) );
  nand02 U3362 ( .Y(n6185), .A0(n6179), .A1(n6186) );
  nand02 U3363 ( .Y(n6187), .A0(n6179), .A1(n6188) );
  nand02 U3364 ( .Y(n6189), .A0(n6180), .A1(n6190) );
  nand02 U3365 ( .Y(n6191), .A0(n6180), .A1(n6192) );
  nand02 U3366 ( .Y(n6193), .A0(n6180), .A1(n6194) );
  nand02 U3367 ( .Y(n6195), .A0(n6180), .A1(n6196) );
  nand02 U3368 ( .Y(n6197), .A0(n6175), .A1(n6176) );
  inv01 U3369 ( .Y(n6182), .A(n6197) );
  nand02 U3370 ( .Y(n6198), .A0(n6175), .A1(n6176) );
  inv01 U3371 ( .Y(n6184), .A(n6198) );
  nand02 U3372 ( .Y(n6199), .A0(n6175), .A1(n6177) );
  inv01 U3373 ( .Y(n6186), .A(n6199) );
  nand02 U3374 ( .Y(n6200), .A0(n6175), .A1(n6178) );
  inv01 U3375 ( .Y(n6188), .A(n6200) );
  nand02 U3376 ( .Y(n6201), .A0(n6176), .A1(n6177) );
  inv01 U3377 ( .Y(n6190), .A(n6201) );
  nand02 U3378 ( .Y(n6202), .A0(n6176), .A1(n6178) );
  inv01 U3379 ( .Y(n6192), .A(n6202) );
  nand02 U3380 ( .Y(n6203), .A0(n6177), .A1(n6179) );
  inv01 U3381 ( .Y(n6194), .A(n6203) );
  nand02 U3382 ( .Y(n6204), .A0(n6178), .A1(n6179) );
  inv01 U3383 ( .Y(n6196), .A(n6204) );
  nand02 U3384 ( .Y(n6205), .A0(n6181), .A1(n6183) );
  inv01 U3385 ( .Y(n6206), .A(n6205) );
  nand02 U3386 ( .Y(n6207), .A0(n6185), .A1(n6187) );
  inv01 U3387 ( .Y(n6208), .A(n6207) );
  nand02 U3388 ( .Y(n6209), .A0(n6206), .A1(n6208) );
  inv01 U3389 ( .Y(n6173), .A(n6209) );
  nand02 U3390 ( .Y(n6210), .A0(n6189), .A1(n6191) );
  inv01 U3391 ( .Y(n6211), .A(n6210) );
  nand02 U3392 ( .Y(n6212), .A0(n6193), .A1(n6195) );
  inv01 U3393 ( .Y(n6213), .A(n6212) );
  nand02 U3394 ( .Y(n6214), .A0(n6211), .A1(n6213) );
  inv01 U3395 ( .Y(n6174), .A(n6214) );
  inv02 U3396 ( .Y(n7858), .A(n7438) );
  nand02 U3397 ( .Y(n7971), .A0(n6215), .A1(n6216) );
  inv02 U3398 ( .Y(n6217), .A(n7649) );
  inv02 U3399 ( .Y(n6218), .A(n7578) );
  inv02 U3400 ( .Y(n6219), .A(n7594) );
  inv02 U3401 ( .Y(n6220), .A(n7825) );
  inv02 U3402 ( .Y(n6221), .A(n7819) );
  inv02 U3403 ( .Y(n6222), .A(n7827) );
  nand02 U3404 ( .Y(n6223), .A0(n6219), .A1(n6224) );
  nand02 U3405 ( .Y(n6225), .A0(n6220), .A1(n6226) );
  nand02 U3406 ( .Y(n6227), .A0(n6221), .A1(n6228) );
  nand02 U3407 ( .Y(n6229), .A0(n6221), .A1(n6230) );
  nand02 U3408 ( .Y(n6231), .A0(n6222), .A1(n6232) );
  nand02 U3409 ( .Y(n6233), .A0(n6222), .A1(n6234) );
  nand02 U3410 ( .Y(n6235), .A0(n6222), .A1(n6236) );
  nand02 U3411 ( .Y(n6237), .A0(n6222), .A1(n6238) );
  nand02 U3412 ( .Y(n6239), .A0(n6217), .A1(n6218) );
  inv01 U3413 ( .Y(n6224), .A(n6239) );
  nand02 U3414 ( .Y(n6240), .A0(n6217), .A1(n6218) );
  inv01 U3415 ( .Y(n6226), .A(n6240) );
  nand02 U3416 ( .Y(n6241), .A0(n6217), .A1(n6219) );
  inv01 U3417 ( .Y(n6228), .A(n6241) );
  nand02 U3418 ( .Y(n6242), .A0(n6217), .A1(n6220) );
  inv01 U3419 ( .Y(n6230), .A(n6242) );
  nand02 U3420 ( .Y(n6243), .A0(n6218), .A1(n6219) );
  inv01 U3421 ( .Y(n6232), .A(n6243) );
  nand02 U3422 ( .Y(n6244), .A0(n6218), .A1(n6220) );
  inv01 U3423 ( .Y(n6234), .A(n6244) );
  nand02 U3424 ( .Y(n6245), .A0(n6219), .A1(n6221) );
  inv01 U3425 ( .Y(n6236), .A(n6245) );
  nand02 U3426 ( .Y(n6246), .A0(n6220), .A1(n6221) );
  inv01 U3427 ( .Y(n6238), .A(n6246) );
  nand02 U3428 ( .Y(n6247), .A0(n6223), .A1(n6225) );
  inv01 U3429 ( .Y(n6248), .A(n6247) );
  nand02 U3430 ( .Y(n6249), .A0(n6227), .A1(n6229) );
  inv01 U3431 ( .Y(n6250), .A(n6249) );
  nand02 U3432 ( .Y(n6251), .A0(n6248), .A1(n6250) );
  inv01 U3433 ( .Y(n6215), .A(n6251) );
  nand02 U3434 ( .Y(n6252), .A0(n6231), .A1(n6233) );
  inv01 U3435 ( .Y(n6253), .A(n6252) );
  nand02 U3436 ( .Y(n6254), .A0(n6235), .A1(n6237) );
  inv01 U3437 ( .Y(n6255), .A(n6254) );
  nand02 U3438 ( .Y(n6256), .A0(n6253), .A1(n6255) );
  inv01 U3439 ( .Y(n6216), .A(n6256) );
  nand02 U3440 ( .Y(n7960), .A0(n6257), .A1(n6258) );
  inv02 U3441 ( .Y(n6259), .A(n7897) );
  inv02 U3442 ( .Y(n6260), .A(n7848) );
  inv02 U3443 ( .Y(n6261), .A(n7871) );
  inv02 U3444 ( .Y(n6262), .A(n7655) );
  inv02 U3445 ( .Y(n6263), .A(n7615) );
  inv02 U3446 ( .Y(n6264), .A(n7678) );
  nand02 U3447 ( .Y(n6265), .A0(n6261), .A1(n6266) );
  nand02 U3448 ( .Y(n6267), .A0(n6262), .A1(n6268) );
  nand02 U3449 ( .Y(n6269), .A0(n6263), .A1(n6270) );
  nand02 U3450 ( .Y(n6271), .A0(n6263), .A1(n6272) );
  nand02 U3451 ( .Y(n6273), .A0(n6264), .A1(n6274) );
  nand02 U3452 ( .Y(n6275), .A0(n6264), .A1(n6276) );
  nand02 U3453 ( .Y(n6277), .A0(n6264), .A1(n6278) );
  nand02 U3454 ( .Y(n6279), .A0(n6264), .A1(n6280) );
  nand02 U3455 ( .Y(n6281), .A0(n6259), .A1(n6260) );
  inv01 U3456 ( .Y(n6266), .A(n6281) );
  nand02 U3457 ( .Y(n6282), .A0(n6259), .A1(n6260) );
  inv01 U3458 ( .Y(n6268), .A(n6282) );
  nand02 U3459 ( .Y(n6283), .A0(n6259), .A1(n6261) );
  inv01 U3460 ( .Y(n6270), .A(n6283) );
  nand02 U3461 ( .Y(n6284), .A0(n6259), .A1(n6262) );
  inv01 U3462 ( .Y(n6272), .A(n6284) );
  nand02 U3463 ( .Y(n6285), .A0(n6260), .A1(n6261) );
  inv01 U3464 ( .Y(n6274), .A(n6285) );
  nand02 U3465 ( .Y(n6286), .A0(n6260), .A1(n6262) );
  inv01 U3466 ( .Y(n6276), .A(n6286) );
  nand02 U3467 ( .Y(n6287), .A0(n6261), .A1(n6263) );
  inv01 U3468 ( .Y(n6278), .A(n6287) );
  nand02 U3469 ( .Y(n6288), .A0(n6262), .A1(n6263) );
  inv01 U3470 ( .Y(n6280), .A(n6288) );
  nand02 U3471 ( .Y(n6289), .A0(n6265), .A1(n6267) );
  inv01 U3472 ( .Y(n6290), .A(n6289) );
  nand02 U3473 ( .Y(n6291), .A0(n6269), .A1(n6271) );
  inv01 U3474 ( .Y(n6292), .A(n6291) );
  nand02 U3475 ( .Y(n6293), .A0(n6290), .A1(n6292) );
  inv01 U3476 ( .Y(n6257), .A(n6293) );
  nand02 U3477 ( .Y(n6294), .A0(n6273), .A1(n6275) );
  inv01 U3478 ( .Y(n6295), .A(n6294) );
  nand02 U3479 ( .Y(n6296), .A0(n6277), .A1(n6279) );
  inv01 U3480 ( .Y(n6297), .A(n6296) );
  nand02 U3481 ( .Y(n6298), .A0(n6295), .A1(n6297) );
  inv01 U3482 ( .Y(n6258), .A(n6298) );
  nand02 U3483 ( .Y(n7870), .A0(n6299), .A1(n6300) );
  inv02 U3484 ( .Y(n6301), .A(n7846) );
  inv02 U3485 ( .Y(n6302), .A(n7872) );
  inv02 U3486 ( .Y(n6303), .A(n7871) );
  inv02 U3487 ( .Y(n6304), .A(n7624) );
  inv02 U3488 ( .Y(n6305), .A(n7283) );
  inv02 U3489 ( .Y(n6306), .A(n7677) );
  nand02 U3490 ( .Y(n6307), .A0(n6303), .A1(n6308) );
  nand02 U3491 ( .Y(n6309), .A0(n6304), .A1(n6310) );
  nand02 U3492 ( .Y(n6311), .A0(n6305), .A1(n6312) );
  nand02 U3493 ( .Y(n6313), .A0(n6305), .A1(n6314) );
  nand02 U3494 ( .Y(n6315), .A0(n6306), .A1(n6316) );
  nand02 U3495 ( .Y(n6317), .A0(n6306), .A1(n6318) );
  nand02 U3496 ( .Y(n6319), .A0(n6306), .A1(n6320) );
  nand02 U3497 ( .Y(n6321), .A0(n6306), .A1(n6322) );
  nand02 U3498 ( .Y(n6323), .A0(n6301), .A1(n6302) );
  inv01 U3499 ( .Y(n6308), .A(n6323) );
  nand02 U3500 ( .Y(n6324), .A0(n6301), .A1(n6302) );
  inv01 U3501 ( .Y(n6310), .A(n6324) );
  nand02 U3502 ( .Y(n6325), .A0(n6301), .A1(n6303) );
  inv01 U3503 ( .Y(n6312), .A(n6325) );
  nand02 U3504 ( .Y(n6326), .A0(n6301), .A1(n6304) );
  inv01 U3505 ( .Y(n6314), .A(n6326) );
  nand02 U3506 ( .Y(n6327), .A0(n6302), .A1(n6303) );
  inv01 U3507 ( .Y(n6316), .A(n6327) );
  nand02 U3508 ( .Y(n6328), .A0(n6302), .A1(n6304) );
  inv01 U3509 ( .Y(n6318), .A(n6328) );
  nand02 U3510 ( .Y(n6329), .A0(n6303), .A1(n6305) );
  inv01 U3511 ( .Y(n6320), .A(n6329) );
  nand02 U3512 ( .Y(n6330), .A0(n6304), .A1(n6305) );
  inv01 U3513 ( .Y(n6322), .A(n6330) );
  nand02 U3514 ( .Y(n6331), .A0(n6307), .A1(n6309) );
  inv01 U3515 ( .Y(n6332), .A(n6331) );
  nand02 U3516 ( .Y(n6333), .A0(n6311), .A1(n6313) );
  inv01 U3517 ( .Y(n6334), .A(n6333) );
  nand02 U3518 ( .Y(n6335), .A0(n6332), .A1(n6334) );
  inv01 U3519 ( .Y(n6299), .A(n6335) );
  nand02 U3520 ( .Y(n6336), .A0(n6315), .A1(n6317) );
  inv01 U3521 ( .Y(n6337), .A(n6336) );
  nand02 U3522 ( .Y(n6338), .A0(n6319), .A1(n6321) );
  inv01 U3523 ( .Y(n6339), .A(n6338) );
  nand02 U3524 ( .Y(n6340), .A0(n6337), .A1(n6339) );
  inv01 U3525 ( .Y(n6300), .A(n6340) );
  nand02 U3526 ( .Y(n7884), .A0(n6341), .A1(n6342) );
  inv02 U3527 ( .Y(n6343), .A(n7853) );
  inv02 U3528 ( .Y(n6344), .A(n7886) );
  inv02 U3529 ( .Y(n6345), .A(n7885) );
  inv02 U3530 ( .Y(n6346), .A(n7624) );
  inv02 U3531 ( .Y(n6347), .A(n7283) );
  inv02 U3532 ( .Y(n6348), .A(n7677) );
  nand02 U3533 ( .Y(n6349), .A0(n6345), .A1(n6350) );
  nand02 U3534 ( .Y(n6351), .A0(n6346), .A1(n6352) );
  nand02 U3535 ( .Y(n6353), .A0(n6347), .A1(n6354) );
  nand02 U3536 ( .Y(n6355), .A0(n6347), .A1(n6356) );
  nand02 U3537 ( .Y(n6357), .A0(n6348), .A1(n6358) );
  nand02 U3538 ( .Y(n6359), .A0(n6348), .A1(n6360) );
  nand02 U3539 ( .Y(n6361), .A0(n6348), .A1(n6362) );
  nand02 U3540 ( .Y(n6363), .A0(n6348), .A1(n6364) );
  nand02 U3541 ( .Y(n6365), .A0(n6343), .A1(n6344) );
  inv01 U3542 ( .Y(n6350), .A(n6365) );
  nand02 U3543 ( .Y(n6366), .A0(n6343), .A1(n6344) );
  inv01 U3544 ( .Y(n6352), .A(n6366) );
  nand02 U3545 ( .Y(n6367), .A0(n6343), .A1(n6345) );
  inv01 U3546 ( .Y(n6354), .A(n6367) );
  nand02 U3547 ( .Y(n6368), .A0(n6343), .A1(n6346) );
  inv01 U3548 ( .Y(n6356), .A(n6368) );
  nand02 U3549 ( .Y(n6369), .A0(n6344), .A1(n6345) );
  inv01 U3550 ( .Y(n6358), .A(n6369) );
  nand02 U3551 ( .Y(n6370), .A0(n6344), .A1(n6346) );
  inv01 U3552 ( .Y(n6360), .A(n6370) );
  nand02 U3553 ( .Y(n6371), .A0(n6345), .A1(n6347) );
  inv01 U3554 ( .Y(n6362), .A(n6371) );
  nand02 U3555 ( .Y(n6372), .A0(n6346), .A1(n6347) );
  inv01 U3556 ( .Y(n6364), .A(n6372) );
  nand02 U3557 ( .Y(n6373), .A0(n6349), .A1(n6351) );
  inv01 U3558 ( .Y(n6374), .A(n6373) );
  nand02 U3559 ( .Y(n6375), .A0(n6353), .A1(n6355) );
  inv01 U3560 ( .Y(n6376), .A(n6375) );
  nand02 U3561 ( .Y(n6377), .A0(n6374), .A1(n6376) );
  inv01 U3562 ( .Y(n6341), .A(n6377) );
  nand02 U3563 ( .Y(n6378), .A0(n6357), .A1(n6359) );
  inv01 U3564 ( .Y(n6379), .A(n6378) );
  nand02 U3565 ( .Y(n6380), .A0(n6361), .A1(n6363) );
  inv01 U3566 ( .Y(n6381), .A(n6380) );
  nand02 U3567 ( .Y(n6382), .A0(n6379), .A1(n6381) );
  inv01 U3568 ( .Y(n6342), .A(n6382) );
  inv02 U3569 ( .Y(n7825), .A(n7587) );
  inv02 U3570 ( .Y(n7827), .A(n7450) );
  inv02 U3571 ( .Y(n7871), .A(n7962) );
  inv02 U3572 ( .Y(n7885), .A(n7968) );
  nand02 U3573 ( .Y(n7970), .A0(n6383), .A1(n6384) );
  inv02 U3574 ( .Y(n6385), .A(n7923) );
  inv02 U3575 ( .Y(n6386), .A(n7861) );
  inv02 U3576 ( .Y(n6387), .A(n7958) );
  inv02 U3577 ( .Y(n6388), .A(n7653) );
  inv02 U3578 ( .Y(n6389), .A(n7615) );
  inv02 U3579 ( .Y(n6390), .A(n7678) );
  nand02 U3580 ( .Y(n6391), .A0(n6387), .A1(n6392) );
  nand02 U3581 ( .Y(n6393), .A0(n6388), .A1(n6394) );
  nand02 U3582 ( .Y(n6395), .A0(n6389), .A1(n6396) );
  nand02 U3583 ( .Y(n6397), .A0(n6389), .A1(n6398) );
  nand02 U3584 ( .Y(n6399), .A0(n6390), .A1(n6400) );
  nand02 U3585 ( .Y(n6401), .A0(n6390), .A1(n6402) );
  nand02 U3586 ( .Y(n6403), .A0(n6390), .A1(n6404) );
  nand02 U3587 ( .Y(n6405), .A0(n6390), .A1(n6406) );
  nand02 U3588 ( .Y(n6407), .A0(n6385), .A1(n6386) );
  inv01 U3589 ( .Y(n6392), .A(n6407) );
  nand02 U3590 ( .Y(n6408), .A0(n6385), .A1(n6386) );
  inv01 U3591 ( .Y(n6394), .A(n6408) );
  nand02 U3592 ( .Y(n6409), .A0(n6385), .A1(n6387) );
  inv01 U3593 ( .Y(n6396), .A(n6409) );
  nand02 U3594 ( .Y(n6410), .A0(n6385), .A1(n6388) );
  inv01 U3595 ( .Y(n6398), .A(n6410) );
  nand02 U3596 ( .Y(n6411), .A0(n6386), .A1(n6387) );
  inv01 U3597 ( .Y(n6400), .A(n6411) );
  nand02 U3598 ( .Y(n6412), .A0(n6386), .A1(n6388) );
  inv01 U3599 ( .Y(n6402), .A(n6412) );
  nand02 U3600 ( .Y(n6413), .A0(n6387), .A1(n6389) );
  inv01 U3601 ( .Y(n6404), .A(n6413) );
  nand02 U3602 ( .Y(n6414), .A0(n6388), .A1(n6389) );
  inv01 U3603 ( .Y(n6406), .A(n6414) );
  nand02 U3604 ( .Y(n6415), .A0(n6391), .A1(n6393) );
  inv01 U3605 ( .Y(n6416), .A(n6415) );
  nand02 U3606 ( .Y(n6417), .A0(n6395), .A1(n6397) );
  inv01 U3607 ( .Y(n6418), .A(n6417) );
  nand02 U3608 ( .Y(n6419), .A0(n6416), .A1(n6418) );
  inv01 U3609 ( .Y(n6383), .A(n6419) );
  nand02 U3610 ( .Y(n6420), .A0(n6399), .A1(n6401) );
  inv01 U3611 ( .Y(n6421), .A(n6420) );
  nand02 U3612 ( .Y(n6422), .A0(n6403), .A1(n6405) );
  inv01 U3613 ( .Y(n6423), .A(n6422) );
  nand02 U3614 ( .Y(n6424), .A0(n6421), .A1(n6423) );
  inv01 U3615 ( .Y(n6384), .A(n6424) );
  inv02 U3616 ( .Y(n7958), .A(n7971) );
  nand02 U3617 ( .Y(n7918), .A0(n6425), .A1(n6426) );
  inv02 U3618 ( .Y(n6427), .A(n7639) );
  inv02 U3619 ( .Y(n6428), .A(n7586) );
  inv02 U3620 ( .Y(n6429), .A(n7596) );
  inv02 U3621 ( .Y(n6430), .A(n7862) );
  inv02 U3622 ( .Y(n6431), .A(n7861) );
  inv02 U3623 ( .Y(n6432), .A(n7920) );
  nand02 U3624 ( .Y(n6433), .A0(n6429), .A1(n6434) );
  nand02 U3625 ( .Y(n6435), .A0(n6430), .A1(n6436) );
  nand02 U3626 ( .Y(n6437), .A0(n6431), .A1(n6438) );
  nand02 U3627 ( .Y(n6439), .A0(n6431), .A1(n6440) );
  nand02 U3628 ( .Y(n6441), .A0(n6432), .A1(n6442) );
  nand02 U3629 ( .Y(n6443), .A0(n6432), .A1(n6444) );
  nand02 U3630 ( .Y(n6445), .A0(n6432), .A1(n6446) );
  nand02 U3631 ( .Y(n6447), .A0(n6432), .A1(n6448) );
  nand02 U3632 ( .Y(n6449), .A0(n6427), .A1(n6428) );
  inv01 U3633 ( .Y(n6434), .A(n6449) );
  nand02 U3634 ( .Y(n6450), .A0(n6427), .A1(n6428) );
  inv01 U3635 ( .Y(n6436), .A(n6450) );
  nand02 U3636 ( .Y(n6451), .A0(n6427), .A1(n6429) );
  inv01 U3637 ( .Y(n6438), .A(n6451) );
  nand02 U3638 ( .Y(n6452), .A0(n6427), .A1(n6430) );
  inv01 U3639 ( .Y(n6440), .A(n6452) );
  nand02 U3640 ( .Y(n6453), .A0(n6428), .A1(n6429) );
  inv01 U3641 ( .Y(n6442), .A(n6453) );
  nand02 U3642 ( .Y(n6454), .A0(n6428), .A1(n6430) );
  inv01 U3643 ( .Y(n6444), .A(n6454) );
  nand02 U3644 ( .Y(n6455), .A0(n6429), .A1(n6431) );
  inv01 U3645 ( .Y(n6446), .A(n6455) );
  nand02 U3646 ( .Y(n6456), .A0(n6430), .A1(n6431) );
  inv01 U3647 ( .Y(n6448), .A(n6456) );
  nand02 U3648 ( .Y(n6457), .A0(n6433), .A1(n6435) );
  inv01 U3649 ( .Y(n6458), .A(n6457) );
  nand02 U3650 ( .Y(n6459), .A0(n6437), .A1(n6439) );
  inv01 U3651 ( .Y(n6460), .A(n6459) );
  nand02 U3652 ( .Y(n6461), .A0(n6458), .A1(n6460) );
  inv01 U3653 ( .Y(n6425), .A(n6461) );
  nand02 U3654 ( .Y(n6462), .A0(n6441), .A1(n6443) );
  inv01 U3655 ( .Y(n6463), .A(n6462) );
  nand02 U3656 ( .Y(n6464), .A0(n6445), .A1(n6447) );
  inv01 U3657 ( .Y(n6465), .A(n6464) );
  nand02 U3658 ( .Y(n6466), .A0(n6463), .A1(n6465) );
  inv01 U3659 ( .Y(n6426), .A(n6466) );
  inv02 U3660 ( .Y(n7862), .A(n7563) );
  inv02 U3661 ( .Y(n7920), .A(n7459) );
  nand02 U3662 ( .Y(n7929), .A0(n6467), .A1(n6468) );
  inv02 U3663 ( .Y(n6469), .A(n7640) );
  inv02 U3664 ( .Y(n6470), .A(n7431) );
  inv02 U3665 ( .Y(n6471), .A(n7919) );
  inv02 U3666 ( .Y(n6472), .A(n7930) );
  inv02 U3667 ( .Y(n6473), .A(n7586) );
  inv02 U3668 ( .Y(n6474), .A(n7931) );
  nand02 U3669 ( .Y(n6475), .A0(n6471), .A1(n6476) );
  nand02 U3670 ( .Y(n6477), .A0(n6472), .A1(n6478) );
  nand02 U3671 ( .Y(n6479), .A0(n6473), .A1(n6480) );
  nand02 U3672 ( .Y(n6481), .A0(n6473), .A1(n6482) );
  nand02 U3673 ( .Y(n6483), .A0(n6474), .A1(n6484) );
  nand02 U3674 ( .Y(n6485), .A0(n6474), .A1(n6486) );
  nand02 U3675 ( .Y(n6487), .A0(n6474), .A1(n6488) );
  nand02 U3676 ( .Y(n6489), .A0(n6474), .A1(n6490) );
  nand02 U3677 ( .Y(n6491), .A0(n6469), .A1(n6470) );
  inv01 U3678 ( .Y(n6476), .A(n6491) );
  nand02 U3679 ( .Y(n6492), .A0(n6469), .A1(n6470) );
  inv01 U3680 ( .Y(n6478), .A(n6492) );
  nand02 U3681 ( .Y(n6493), .A0(n6469), .A1(n6471) );
  inv01 U3682 ( .Y(n6480), .A(n6493) );
  nand02 U3683 ( .Y(n6494), .A0(n6469), .A1(n6472) );
  inv01 U3684 ( .Y(n6482), .A(n6494) );
  nand02 U3685 ( .Y(n6495), .A0(n6470), .A1(n6471) );
  inv01 U3686 ( .Y(n6484), .A(n6495) );
  nand02 U3687 ( .Y(n6496), .A0(n6470), .A1(n6472) );
  inv01 U3688 ( .Y(n6486), .A(n6496) );
  nand02 U3689 ( .Y(n6497), .A0(n6471), .A1(n6473) );
  inv01 U3690 ( .Y(n6488), .A(n6497) );
  nand02 U3691 ( .Y(n6498), .A0(n6472), .A1(n6473) );
  inv01 U3692 ( .Y(n6490), .A(n6498) );
  nand02 U3693 ( .Y(n6499), .A0(n6475), .A1(n6477) );
  inv01 U3694 ( .Y(n6500), .A(n6499) );
  nand02 U3695 ( .Y(n6501), .A0(n6479), .A1(n6481) );
  inv01 U3696 ( .Y(n6502), .A(n6501) );
  nand02 U3697 ( .Y(n6503), .A0(n6500), .A1(n6502) );
  inv01 U3698 ( .Y(n6467), .A(n6503) );
  nand02 U3699 ( .Y(n6504), .A0(n6483), .A1(n6485) );
  inv01 U3700 ( .Y(n6505), .A(n6504) );
  nand02 U3701 ( .Y(n6506), .A0(n6487), .A1(n6489) );
  inv01 U3702 ( .Y(n6507), .A(n6506) );
  nand02 U3703 ( .Y(n6508), .A0(n6505), .A1(n6507) );
  inv01 U3704 ( .Y(n6468), .A(n6508) );
  nand02 U3705 ( .Y(n7915), .A0(n6509), .A1(n6510) );
  inv02 U3706 ( .Y(n6511), .A(n7821) );
  inv02 U3707 ( .Y(n6512), .A(n7917) );
  inv02 U3708 ( .Y(n6513), .A(n7916) );
  inv02 U3709 ( .Y(n6514), .A(n7676) );
  inv02 U3710 ( .Y(n6515), .A(n7678) );
  inv02 U3711 ( .Y(n6516), .A(n7648) );
  nand02 U3712 ( .Y(n6517), .A0(n6513), .A1(n6518) );
  nand02 U3713 ( .Y(n6519), .A0(n6514), .A1(n6520) );
  nand02 U3714 ( .Y(n6521), .A0(n6515), .A1(n6522) );
  nand02 U3715 ( .Y(n6523), .A0(n6515), .A1(n6524) );
  nand02 U3716 ( .Y(n6525), .A0(n6516), .A1(n6526) );
  nand02 U3717 ( .Y(n6527), .A0(n6516), .A1(n6528) );
  nand02 U3718 ( .Y(n6529), .A0(n6516), .A1(n6530) );
  nand02 U3719 ( .Y(n6531), .A0(n6516), .A1(n6532) );
  nand02 U3720 ( .Y(n6533), .A0(n6511), .A1(n6512) );
  inv01 U3721 ( .Y(n6518), .A(n6533) );
  nand02 U3722 ( .Y(n6534), .A0(n6511), .A1(n6512) );
  inv01 U3723 ( .Y(n6520), .A(n6534) );
  nand02 U3724 ( .Y(n6535), .A0(n6511), .A1(n6513) );
  inv01 U3725 ( .Y(n6522), .A(n6535) );
  nand02 U3726 ( .Y(n6536), .A0(n6511), .A1(n6514) );
  inv01 U3727 ( .Y(n6524), .A(n6536) );
  nand02 U3728 ( .Y(n6537), .A0(n6512), .A1(n6513) );
  inv01 U3729 ( .Y(n6526), .A(n6537) );
  nand02 U3730 ( .Y(n6538), .A0(n6512), .A1(n6514) );
  inv01 U3731 ( .Y(n6528), .A(n6538) );
  nand02 U3732 ( .Y(n6539), .A0(n6513), .A1(n6515) );
  inv01 U3733 ( .Y(n6530), .A(n6539) );
  nand02 U3734 ( .Y(n6540), .A0(n6514), .A1(n6515) );
  inv01 U3735 ( .Y(n6532), .A(n6540) );
  nand02 U3736 ( .Y(n6541), .A0(n6517), .A1(n6519) );
  inv01 U3737 ( .Y(n6542), .A(n6541) );
  nand02 U3738 ( .Y(n6543), .A0(n6521), .A1(n6523) );
  inv01 U3739 ( .Y(n6544), .A(n6543) );
  nand02 U3740 ( .Y(n6545), .A0(n6542), .A1(n6544) );
  inv01 U3741 ( .Y(n6509), .A(n6545) );
  nand02 U3742 ( .Y(n6546), .A0(n6525), .A1(n6527) );
  inv01 U3743 ( .Y(n6547), .A(n6546) );
  nand02 U3744 ( .Y(n6548), .A0(n6529), .A1(n6531) );
  inv01 U3745 ( .Y(n6549), .A(n6548) );
  nand02 U3746 ( .Y(n6550), .A0(n6547), .A1(n6549) );
  inv01 U3747 ( .Y(n6510), .A(n6550) );
  inv02 U3748 ( .Y(n7931), .A(n7444) );
  inv02 U3749 ( .Y(n7821), .A(n7918) );
  inv01 U3750 ( .Y(n8025), .A(n6551) );
  inv01 U3751 ( .Y(n6552), .A(n8020) );
  inv01 U3752 ( .Y(n6553), .A(n8032) );
  inv01 U3753 ( .Y(n6554), .A(n8021) );
  inv01 U3754 ( .Y(n6555), .A(n4771) );
  nand02 U3755 ( .Y(n6551), .A0(n6556), .A1(n6557) );
  nand02 U3756 ( .Y(n6558), .A0(n6552), .A1(n6553) );
  inv01 U3757 ( .Y(n6556), .A(n6558) );
  nand02 U3758 ( .Y(n6559), .A0(n6554), .A1(n6555) );
  inv01 U3759 ( .Y(n6557), .A(n6559) );
  nand02 U3760 ( .Y(n7926), .A0(n6560), .A1(n6561) );
  inv02 U3761 ( .Y(n6562), .A(n7832) );
  inv02 U3762 ( .Y(n6563), .A(n7928) );
  inv02 U3763 ( .Y(n6564), .A(n7927) );
  inv02 U3764 ( .Y(n6565), .A(n7676) );
  inv02 U3765 ( .Y(n6566), .A(n7678) );
  inv02 U3766 ( .Y(n6567), .A(n7648) );
  nand02 U3767 ( .Y(n6568), .A0(n6564), .A1(n6569) );
  nand02 U3768 ( .Y(n6570), .A0(n6565), .A1(n6571) );
  nand02 U3769 ( .Y(n6572), .A0(n6566), .A1(n6573) );
  nand02 U3770 ( .Y(n6574), .A0(n6566), .A1(n6575) );
  nand02 U3771 ( .Y(n6576), .A0(n6567), .A1(n6577) );
  nand02 U3772 ( .Y(n6578), .A0(n6567), .A1(n6579) );
  nand02 U3773 ( .Y(n6580), .A0(n6567), .A1(n6581) );
  nand02 U3774 ( .Y(n6582), .A0(n6567), .A1(n6583) );
  nand02 U3775 ( .Y(n6584), .A0(n6562), .A1(n6563) );
  inv01 U3776 ( .Y(n6569), .A(n6584) );
  nand02 U3777 ( .Y(n6585), .A0(n6562), .A1(n6563) );
  inv01 U3778 ( .Y(n6571), .A(n6585) );
  nand02 U3779 ( .Y(n6586), .A0(n6562), .A1(n6564) );
  inv01 U3780 ( .Y(n6573), .A(n6586) );
  nand02 U3781 ( .Y(n6587), .A0(n6562), .A1(n6565) );
  inv01 U3782 ( .Y(n6575), .A(n6587) );
  nand02 U3783 ( .Y(n6588), .A0(n6563), .A1(n6564) );
  inv01 U3784 ( .Y(n6577), .A(n6588) );
  nand02 U3785 ( .Y(n6589), .A0(n6563), .A1(n6565) );
  inv01 U3786 ( .Y(n6579), .A(n6589) );
  nand02 U3787 ( .Y(n6590), .A0(n6564), .A1(n6566) );
  inv01 U3788 ( .Y(n6581), .A(n6590) );
  nand02 U3789 ( .Y(n6591), .A0(n6565), .A1(n6566) );
  inv01 U3790 ( .Y(n6583), .A(n6591) );
  nand02 U3791 ( .Y(n6592), .A0(n6568), .A1(n6570) );
  inv01 U3792 ( .Y(n6593), .A(n6592) );
  nand02 U3793 ( .Y(n6594), .A0(n6572), .A1(n6574) );
  inv01 U3794 ( .Y(n6595), .A(n6594) );
  nand02 U3795 ( .Y(n6596), .A0(n6593), .A1(n6595) );
  inv01 U3796 ( .Y(n6560), .A(n6596) );
  nand02 U3797 ( .Y(n6597), .A0(n6576), .A1(n6578) );
  inv01 U3798 ( .Y(n6598), .A(n6597) );
  nand02 U3799 ( .Y(n6599), .A0(n6580), .A1(n6582) );
  inv01 U3800 ( .Y(n6600), .A(n6599) );
  nand02 U3801 ( .Y(n6601), .A0(n6598), .A1(n6600) );
  inv01 U3802 ( .Y(n6561), .A(n6601) );
  inv02 U3803 ( .Y(n7832), .A(n7929) );
  inv01 U3804 ( .Y(n8026), .A(n6602) );
  inv01 U3805 ( .Y(n6603), .A(n8019) );
  inv01 U3806 ( .Y(n6604), .A(n8018) );
  inv01 U3807 ( .Y(n6605), .A(n4748) );
  inv01 U3808 ( .Y(n6606), .A(n6969) );
  nand02 U3809 ( .Y(n6602), .A0(n6607), .A1(n6608) );
  nand02 U3810 ( .Y(n6609), .A0(n6603), .A1(n6604) );
  inv01 U3811 ( .Y(n6607), .A(n6609) );
  nand02 U3812 ( .Y(n6610), .A0(n6605), .A1(n6606) );
  inv01 U3813 ( .Y(n6608), .A(n6610) );
  nand02 U3814 ( .Y(n7907), .A0(n6611), .A1(n6612) );
  inv02 U3815 ( .Y(n6613), .A(n7910) );
  inv02 U3816 ( .Y(n6614), .A(n7909) );
  inv02 U3817 ( .Y(n6615), .A(n7908) );
  inv02 U3818 ( .Y(n6616), .A(n7669) );
  inv02 U3819 ( .Y(n6617), .A(n7678) );
  inv02 U3820 ( .Y(n6618), .A(n7676) );
  nand02 U3821 ( .Y(n6619), .A0(n6615), .A1(n6620) );
  nand02 U3822 ( .Y(n6621), .A0(n6616), .A1(n6622) );
  nand02 U3823 ( .Y(n6623), .A0(n6617), .A1(n6624) );
  nand02 U3824 ( .Y(n6625), .A0(n6617), .A1(n6626) );
  nand02 U3825 ( .Y(n6627), .A0(n6618), .A1(n6628) );
  nand02 U3826 ( .Y(n6629), .A0(n6618), .A1(n6630) );
  nand02 U3827 ( .Y(n6631), .A0(n6618), .A1(n6632) );
  nand02 U3828 ( .Y(n6633), .A0(n6618), .A1(n6634) );
  nand02 U3829 ( .Y(n6635), .A0(n6613), .A1(n6614) );
  inv01 U3830 ( .Y(n6620), .A(n6635) );
  nand02 U3831 ( .Y(n6636), .A0(n6613), .A1(n6614) );
  inv01 U3832 ( .Y(n6622), .A(n6636) );
  nand02 U3833 ( .Y(n6637), .A0(n6613), .A1(n6615) );
  inv01 U3834 ( .Y(n6624), .A(n6637) );
  nand02 U3835 ( .Y(n6638), .A0(n6613), .A1(n6616) );
  inv01 U3836 ( .Y(n6626), .A(n6638) );
  nand02 U3837 ( .Y(n6639), .A0(n6614), .A1(n6615) );
  inv01 U3838 ( .Y(n6628), .A(n6639) );
  nand02 U3839 ( .Y(n6640), .A0(n6614), .A1(n6616) );
  inv01 U3840 ( .Y(n6630), .A(n6640) );
  nand02 U3841 ( .Y(n6641), .A0(n6615), .A1(n6617) );
  inv01 U3842 ( .Y(n6632), .A(n6641) );
  nand02 U3843 ( .Y(n6642), .A0(n6616), .A1(n6617) );
  inv01 U3844 ( .Y(n6634), .A(n6642) );
  nand02 U3845 ( .Y(n6643), .A0(n6619), .A1(n6621) );
  inv01 U3846 ( .Y(n6644), .A(n6643) );
  nand02 U3847 ( .Y(n6645), .A0(n6623), .A1(n6625) );
  inv01 U3848 ( .Y(n6646), .A(n6645) );
  nand02 U3849 ( .Y(n6647), .A0(n6644), .A1(n6646) );
  inv01 U3850 ( .Y(n6611), .A(n6647) );
  nand02 U3851 ( .Y(n6648), .A0(n6627), .A1(n6629) );
  inv01 U3852 ( .Y(n6649), .A(n6648) );
  nand02 U3853 ( .Y(n6650), .A0(n6631), .A1(n6633) );
  inv01 U3854 ( .Y(n6651), .A(n6650) );
  nand02 U3855 ( .Y(n6652), .A0(n6649), .A1(n6651) );
  inv01 U3856 ( .Y(n6612), .A(n6652) );
  inv04 U3857 ( .Y(n7764), .A(n6653) );
  inv01 U3858 ( .Y(n6654), .A(opa_i[8]) );
  inv01 U3859 ( .Y(n6655), .A(opa_i[9]) );
  inv01 U3860 ( .Y(n6656), .A(opa_i[7]) );
  nand02 U3861 ( .Y(n6653), .A0(n6656), .A1(n6657) );
  nand02 U3862 ( .Y(n6658), .A0(n6654), .A1(n6655) );
  inv01 U3863 ( .Y(n6657), .A(n6658) );
  buf08 U3864 ( .Y(n7669), .A(n7896) );
  or02 U3865 ( .Y(n6659), .A0(fract_28_i[24]), .A1(fract_28_i[23]) );
  inv01 U3866 ( .Y(n6660), .A(n6659) );
  inv04 U3867 ( .Y(n7759), .A(n6661) );
  inv01 U3868 ( .Y(n6662), .A(opa_i[15]) );
  inv01 U3869 ( .Y(n6663), .A(opa_i[16]) );
  inv01 U3870 ( .Y(n6664), .A(opa_i[14]) );
  nand02 U3871 ( .Y(n6661), .A0(n6664), .A1(n6665) );
  nand02 U3872 ( .Y(n6666), .A0(n6662), .A1(n6663) );
  inv01 U3873 ( .Y(n6665), .A(n6666) );
  nand02 U3874 ( .Y(n7754), .A0(n6667), .A1(n6668) );
  inv02 U3875 ( .Y(n6669), .A(n7684) );
  inv02 U3876 ( .Y(n6670), .A(n7716) );
  inv02 U3877 ( .Y(n6671), .A(n7713) );
  inv02 U3878 ( .Y(n6672), .A(n____return2766_26_) );
  inv02 U3879 ( .Y(n6673), .A(n____return2766_25_) );
  inv02 U3880 ( .Y(n6674), .A(s_fracto28_1[25]) );
  nand02 U3881 ( .Y(n6675), .A0(n6671), .A1(n6676) );
  nand02 U3882 ( .Y(n6677), .A0(n6672), .A1(n6678) );
  nand02 U3883 ( .Y(n6679), .A0(n6673), .A1(n6680) );
  nand02 U3884 ( .Y(n6681), .A0(n6673), .A1(n6682) );
  nand02 U3885 ( .Y(n6683), .A0(n6674), .A1(n6684) );
  nand02 U3886 ( .Y(n6685), .A0(n6674), .A1(n6686) );
  nand02 U3887 ( .Y(n6687), .A0(n6674), .A1(n6688) );
  nand02 U3888 ( .Y(n6689), .A0(n6674), .A1(n6690) );
  nand02 U3889 ( .Y(n6691), .A0(n6669), .A1(n6670) );
  inv01 U3890 ( .Y(n6676), .A(n6691) );
  nand02 U3891 ( .Y(n6692), .A0(n6669), .A1(n6670) );
  inv01 U3892 ( .Y(n6678), .A(n6692) );
  nand02 U3893 ( .Y(n6693), .A0(n6669), .A1(n6671) );
  inv01 U3894 ( .Y(n6680), .A(n6693) );
  nand02 U3895 ( .Y(n6694), .A0(n6669), .A1(n6672) );
  inv01 U3896 ( .Y(n6682), .A(n6694) );
  nand02 U3897 ( .Y(n6695), .A0(n6670), .A1(n6671) );
  inv01 U3898 ( .Y(n6684), .A(n6695) );
  nand02 U3899 ( .Y(n6696), .A0(n6670), .A1(n6672) );
  inv01 U3900 ( .Y(n6686), .A(n6696) );
  nand02 U3901 ( .Y(n6697), .A0(n6671), .A1(n6673) );
  inv01 U3902 ( .Y(n6688), .A(n6697) );
  nand02 U3903 ( .Y(n6698), .A0(n6672), .A1(n6673) );
  inv01 U3904 ( .Y(n6690), .A(n6698) );
  nand02 U3905 ( .Y(n6699), .A0(n6675), .A1(n6677) );
  inv01 U3906 ( .Y(n6700), .A(n6699) );
  nand02 U3907 ( .Y(n6701), .A0(n6679), .A1(n6681) );
  inv01 U3908 ( .Y(n6702), .A(n6701) );
  nand02 U3909 ( .Y(n6703), .A0(n6700), .A1(n6702) );
  inv01 U3910 ( .Y(n6667), .A(n6703) );
  nand02 U3911 ( .Y(n6704), .A0(n6683), .A1(n6685) );
  inv01 U3912 ( .Y(n6705), .A(n6704) );
  nand02 U3913 ( .Y(n6706), .A0(n6687), .A1(n6689) );
  inv01 U3914 ( .Y(n6707), .A(n6706) );
  nand02 U3915 ( .Y(n6708), .A0(n6705), .A1(n6707) );
  inv01 U3916 ( .Y(n6668), .A(n6708) );
  nand02 U3917 ( .Y(n7864), .A0(n6709), .A1(n6710) );
  inv02 U3918 ( .Y(n6711), .A(n7833) );
  inv02 U3919 ( .Y(n6712), .A(n7830) );
  inv02 U3920 ( .Y(n6713), .A(n7834) );
  inv02 U3921 ( .Y(n6714), .A(n7670) );
  inv02 U3922 ( .Y(n6715), .A(n7677) );
  inv02 U3923 ( .Y(n6716), .A(n7672) );
  nand02 U3924 ( .Y(n6717), .A0(n6713), .A1(n6718) );
  nand02 U3925 ( .Y(n6719), .A0(n6714), .A1(n6720) );
  nand02 U3926 ( .Y(n6721), .A0(n6715), .A1(n6722) );
  nand02 U3927 ( .Y(n6723), .A0(n6715), .A1(n6724) );
  nand02 U3928 ( .Y(n6725), .A0(n6716), .A1(n6726) );
  nand02 U3929 ( .Y(n6727), .A0(n6716), .A1(n6728) );
  nand02 U3930 ( .Y(n6729), .A0(n6716), .A1(n6730) );
  nand02 U3931 ( .Y(n6731), .A0(n6716), .A1(n6732) );
  nand02 U3932 ( .Y(n6733), .A0(n6711), .A1(n6712) );
  inv01 U3933 ( .Y(n6718), .A(n6733) );
  nand02 U3934 ( .Y(n6734), .A0(n6711), .A1(n6712) );
  inv01 U3935 ( .Y(n6720), .A(n6734) );
  nand02 U3936 ( .Y(n6735), .A0(n6711), .A1(n6713) );
  inv01 U3937 ( .Y(n6722), .A(n6735) );
  nand02 U3938 ( .Y(n6736), .A0(n6711), .A1(n6714) );
  inv01 U3939 ( .Y(n6724), .A(n6736) );
  nand02 U3940 ( .Y(n6737), .A0(n6712), .A1(n6713) );
  inv01 U3941 ( .Y(n6726), .A(n6737) );
  nand02 U3942 ( .Y(n6738), .A0(n6712), .A1(n6714) );
  inv01 U3943 ( .Y(n6728), .A(n6738) );
  nand02 U3944 ( .Y(n6739), .A0(n6713), .A1(n6715) );
  inv01 U3945 ( .Y(n6730), .A(n6739) );
  nand02 U3946 ( .Y(n6740), .A0(n6714), .A1(n6715) );
  inv01 U3947 ( .Y(n6732), .A(n6740) );
  nand02 U3948 ( .Y(n6741), .A0(n6717), .A1(n6719) );
  inv01 U3949 ( .Y(n6742), .A(n6741) );
  nand02 U3950 ( .Y(n6743), .A0(n6721), .A1(n6723) );
  inv01 U3951 ( .Y(n6744), .A(n6743) );
  nand02 U3952 ( .Y(n6745), .A0(n6742), .A1(n6744) );
  inv01 U3953 ( .Y(n6709), .A(n6745) );
  nand02 U3954 ( .Y(n6746), .A0(n6725), .A1(n6727) );
  inv01 U3955 ( .Y(n6747), .A(n6746) );
  nand02 U3956 ( .Y(n6748), .A0(n6729), .A1(n6731) );
  inv01 U3957 ( .Y(n6749), .A(n6748) );
  nand02 U3958 ( .Y(n6750), .A0(n6747), .A1(n6749) );
  inv01 U3959 ( .Y(n6710), .A(n6750) );
  nand02 U3960 ( .Y(n7990), .A0(n6751), .A1(n6752) );
  inv02 U3961 ( .Y(n6753), .A(n7831) );
  inv02 U3962 ( .Y(n6754), .A(n7833) );
  inv02 U3963 ( .Y(n6755), .A(n7835) );
  inv02 U3964 ( .Y(n6756), .A(n7670) );
  inv02 U3965 ( .Y(n6757), .A(n7677) );
  inv02 U3966 ( .Y(n6758), .A(n7673) );
  nand02 U3967 ( .Y(n6759), .A0(n6755), .A1(n6760) );
  nand02 U3968 ( .Y(n6761), .A0(n6756), .A1(n6762) );
  nand02 U3969 ( .Y(n6763), .A0(n6757), .A1(n6764) );
  nand02 U3970 ( .Y(n6765), .A0(n6757), .A1(n6766) );
  nand02 U3971 ( .Y(n6767), .A0(n6758), .A1(n6768) );
  nand02 U3972 ( .Y(n6769), .A0(n6758), .A1(n6770) );
  nand02 U3973 ( .Y(n6771), .A0(n6758), .A1(n6772) );
  nand02 U3974 ( .Y(n6773), .A0(n6758), .A1(n6774) );
  nand02 U3975 ( .Y(n6775), .A0(n6753), .A1(n6754) );
  inv01 U3976 ( .Y(n6760), .A(n6775) );
  nand02 U3977 ( .Y(n6776), .A0(n6753), .A1(n6754) );
  inv01 U3978 ( .Y(n6762), .A(n6776) );
  nand02 U3979 ( .Y(n6777), .A0(n6753), .A1(n6755) );
  inv01 U3980 ( .Y(n6764), .A(n6777) );
  nand02 U3981 ( .Y(n6778), .A0(n6753), .A1(n6756) );
  inv01 U3982 ( .Y(n6766), .A(n6778) );
  nand02 U3983 ( .Y(n6779), .A0(n6754), .A1(n6755) );
  inv01 U3984 ( .Y(n6768), .A(n6779) );
  nand02 U3985 ( .Y(n6780), .A0(n6754), .A1(n6756) );
  inv01 U3986 ( .Y(n6770), .A(n6780) );
  nand02 U3987 ( .Y(n6781), .A0(n6755), .A1(n6757) );
  inv01 U3988 ( .Y(n6772), .A(n6781) );
  nand02 U3989 ( .Y(n6782), .A0(n6756), .A1(n6757) );
  inv01 U3990 ( .Y(n6774), .A(n6782) );
  nand02 U3991 ( .Y(n6783), .A0(n6759), .A1(n6761) );
  inv01 U3992 ( .Y(n6784), .A(n6783) );
  nand02 U3993 ( .Y(n6785), .A0(n6763), .A1(n6765) );
  inv01 U3994 ( .Y(n6786), .A(n6785) );
  nand02 U3995 ( .Y(n6787), .A0(n6784), .A1(n6786) );
  inv01 U3996 ( .Y(n6751), .A(n6787) );
  nand02 U3997 ( .Y(n6788), .A0(n6767), .A1(n6769) );
  inv01 U3998 ( .Y(n6789), .A(n6788) );
  nand02 U3999 ( .Y(n6790), .A0(n6771), .A1(n6773) );
  inv01 U4000 ( .Y(n6791), .A(n6790) );
  nand02 U4001 ( .Y(n6792), .A0(n6789), .A1(n6791) );
  inv01 U4002 ( .Y(n6752), .A(n6792) );
  buf08 U4003 ( .Y(n7670), .A(n7826) );
  nand02 U4004 ( .Y(n7838), .A0(n6793), .A1(n6794) );
  inv02 U4005 ( .Y(n6795), .A(n7842) );
  inv02 U4006 ( .Y(n6796), .A(n7840) );
  inv02 U4007 ( .Y(n6797), .A(n7839) );
  inv02 U4008 ( .Y(n6798), .A(n7671) );
  inv02 U4009 ( .Y(n6799), .A(n7670) );
  inv02 U4010 ( .Y(n6800), .A(n7678) );
  nand02 U4011 ( .Y(n6801), .A0(n6797), .A1(n6802) );
  nand02 U4012 ( .Y(n6803), .A0(n6798), .A1(n6804) );
  nand02 U4013 ( .Y(n6805), .A0(n6799), .A1(n6806) );
  nand02 U4014 ( .Y(n6807), .A0(n6799), .A1(n6808) );
  nand02 U4015 ( .Y(n6809), .A0(n6800), .A1(n6810) );
  nand02 U4016 ( .Y(n6811), .A0(n6800), .A1(n6812) );
  nand02 U4017 ( .Y(n6813), .A0(n6800), .A1(n6814) );
  nand02 U4018 ( .Y(n6815), .A0(n6800), .A1(n6816) );
  nand02 U4019 ( .Y(n6817), .A0(n6795), .A1(n6796) );
  inv01 U4020 ( .Y(n6802), .A(n6817) );
  nand02 U4021 ( .Y(n6818), .A0(n6795), .A1(n6796) );
  inv01 U4022 ( .Y(n6804), .A(n6818) );
  nand02 U4023 ( .Y(n6819), .A0(n6795), .A1(n6797) );
  inv01 U4024 ( .Y(n6806), .A(n6819) );
  nand02 U4025 ( .Y(n6820), .A0(n6795), .A1(n6798) );
  inv01 U4026 ( .Y(n6808), .A(n6820) );
  nand02 U4027 ( .Y(n6821), .A0(n6796), .A1(n6797) );
  inv01 U4028 ( .Y(n6810), .A(n6821) );
  nand02 U4029 ( .Y(n6822), .A0(n6796), .A1(n6798) );
  inv01 U4030 ( .Y(n6812), .A(n6822) );
  nand02 U4031 ( .Y(n6823), .A0(n6797), .A1(n6799) );
  inv01 U4032 ( .Y(n6814), .A(n6823) );
  nand02 U4033 ( .Y(n6824), .A0(n6798), .A1(n6799) );
  inv01 U4034 ( .Y(n6816), .A(n6824) );
  nand02 U4035 ( .Y(n6825), .A0(n6801), .A1(n6803) );
  inv01 U4036 ( .Y(n6826), .A(n6825) );
  nand02 U4037 ( .Y(n6827), .A0(n6805), .A1(n6807) );
  inv01 U4038 ( .Y(n6828), .A(n6827) );
  nand02 U4039 ( .Y(n6829), .A0(n6826), .A1(n6828) );
  inv01 U4040 ( .Y(n6793), .A(n6829) );
  nand02 U4041 ( .Y(n6830), .A0(n6809), .A1(n6811) );
  inv01 U4042 ( .Y(n6831), .A(n6830) );
  nand02 U4043 ( .Y(n6832), .A0(n6813), .A1(n6815) );
  inv01 U4044 ( .Y(n6833), .A(n6832) );
  nand02 U4045 ( .Y(n6834), .A0(n6831), .A1(n6833) );
  inv01 U4046 ( .Y(n6794), .A(n6834) );
  nand02 U4047 ( .Y(n7979), .A0(n6835), .A1(n6836) );
  inv02 U4048 ( .Y(n6837), .A(n7840) );
  inv02 U4049 ( .Y(n6838), .A(n7839) );
  inv02 U4050 ( .Y(n6839), .A(n7677) );
  inv02 U4051 ( .Y(n6840), .A(n7676) );
  inv02 U4052 ( .Y(n6841), .A(n7675) );
  nand02 U4053 ( .Y(n6842), .A0(n6838), .A1(n6843) );
  nand02 U4054 ( .Y(n6844), .A0(n6839), .A1(n6845) );
  nand02 U4055 ( .Y(n6846), .A0(n6840), .A1(n6847) );
  nand02 U4056 ( .Y(n6848), .A0(n6840), .A1(n6849) );
  nand02 U4057 ( .Y(n6850), .A0(n6841), .A1(n6851) );
  nand02 U4058 ( .Y(n6852), .A0(n6841), .A1(n6853) );
  nand02 U4059 ( .Y(n6854), .A0(n6841), .A1(n6855) );
  nand02 U4060 ( .Y(n6856), .A0(n6841), .A1(n6857) );
  nand02 U4061 ( .Y(n6858), .A0(n6837), .A1(n5608) );
  inv01 U4062 ( .Y(n6843), .A(n6858) );
  nand02 U4063 ( .Y(n6859), .A0(n6837), .A1(n5608) );
  inv01 U4064 ( .Y(n6845), .A(n6859) );
  nand02 U4065 ( .Y(n6860), .A0(n6837), .A1(n6838) );
  inv01 U4066 ( .Y(n6847), .A(n6860) );
  nand02 U4067 ( .Y(n6861), .A0(n6837), .A1(n6839) );
  inv01 U4068 ( .Y(n6849), .A(n6861) );
  nand02 U4069 ( .Y(n6862), .A0(n5608), .A1(n6838) );
  inv01 U4070 ( .Y(n6851), .A(n6862) );
  nand02 U4071 ( .Y(n6863), .A0(n5608), .A1(n6839) );
  inv01 U4072 ( .Y(n6853), .A(n6863) );
  nand02 U4073 ( .Y(n6864), .A0(n6838), .A1(n6840) );
  inv01 U4074 ( .Y(n6855), .A(n6864) );
  nand02 U4075 ( .Y(n6865), .A0(n6839), .A1(n6840) );
  inv01 U4076 ( .Y(n6857), .A(n6865) );
  nand02 U4077 ( .Y(n6866), .A0(n6842), .A1(n6844) );
  inv01 U4078 ( .Y(n6867), .A(n6866) );
  nand02 U4079 ( .Y(n6868), .A0(n6846), .A1(n6848) );
  inv01 U4080 ( .Y(n6869), .A(n6868) );
  nand02 U4081 ( .Y(n6870), .A0(n6867), .A1(n6869) );
  inv01 U4082 ( .Y(n6835), .A(n6870) );
  nand02 U4083 ( .Y(n6871), .A0(n6850), .A1(n6852) );
  inv01 U4084 ( .Y(n6872), .A(n6871) );
  nand02 U4085 ( .Y(n6873), .A0(n6854), .A1(n6856) );
  inv01 U4086 ( .Y(n6874), .A(n6873) );
  nand02 U4087 ( .Y(n6875), .A0(n6872), .A1(n6874) );
  inv01 U4088 ( .Y(n6836), .A(n6875) );
  inv02 U4089 ( .Y(n7839), .A(n7507) );
  inv02 U4090 ( .Y(n7842), .A(n7571) );
  nand02 U4091 ( .Y(n7948), .A0(n6876), .A1(n6877) );
  inv02 U4092 ( .Y(n6878), .A(n7835) );
  inv02 U4093 ( .Y(n6879), .A(n7935) );
  inv02 U4094 ( .Y(n6880), .A(n7677) );
  inv02 U4095 ( .Y(n6881), .A(n7668) );
  inv02 U4096 ( .Y(n6882), .A(n7675) );
  nand02 U4097 ( .Y(n6883), .A0(n5913), .A1(n6884) );
  nand02 U4098 ( .Y(n6885), .A0(n6880), .A1(n6886) );
  nand02 U4099 ( .Y(n6887), .A0(n6881), .A1(n6888) );
  nand02 U4100 ( .Y(n6889), .A0(n6881), .A1(n6890) );
  nand02 U4101 ( .Y(n6891), .A0(n6882), .A1(n6892) );
  nand02 U4102 ( .Y(n6893), .A0(n6882), .A1(n6894) );
  nand02 U4103 ( .Y(n6895), .A0(n6882), .A1(n6896) );
  nand02 U4104 ( .Y(n6897), .A0(n6882), .A1(n6898) );
  nand02 U4105 ( .Y(n6899), .A0(n6878), .A1(n6879) );
  inv01 U4106 ( .Y(n6884), .A(n6899) );
  nand02 U4107 ( .Y(n6900), .A0(n6878), .A1(n6879) );
  inv01 U4108 ( .Y(n6886), .A(n6900) );
  nand02 U4109 ( .Y(n6901), .A0(n6878), .A1(n6753) );
  inv01 U4110 ( .Y(n6888), .A(n6901) );
  nand02 U4111 ( .Y(n6902), .A0(n6878), .A1(n6880) );
  inv01 U4112 ( .Y(n6890), .A(n6902) );
  nand02 U4113 ( .Y(n6903), .A0(n6879), .A1(n5567) );
  inv01 U4114 ( .Y(n6892), .A(n6903) );
  nand02 U4115 ( .Y(n6904), .A0(n6879), .A1(n6880) );
  inv01 U4116 ( .Y(n6894), .A(n6904) );
  nand02 U4117 ( .Y(n6905), .A0(n5272), .A1(n6881) );
  inv01 U4118 ( .Y(n6896), .A(n6905) );
  nand02 U4119 ( .Y(n6906), .A0(n6880), .A1(n6881) );
  inv01 U4120 ( .Y(n6898), .A(n6906) );
  nand02 U4121 ( .Y(n6907), .A0(n6883), .A1(n6885) );
  inv01 U4122 ( .Y(n6908), .A(n6907) );
  nand02 U4123 ( .Y(n6909), .A0(n6887), .A1(n6889) );
  inv01 U4124 ( .Y(n6910), .A(n6909) );
  nand02 U4125 ( .Y(n6911), .A0(n6908), .A1(n6910) );
  inv01 U4126 ( .Y(n6876), .A(n6911) );
  nand02 U4127 ( .Y(n6912), .A0(n6891), .A1(n6893) );
  inv01 U4128 ( .Y(n6913), .A(n6912) );
  nand02 U4129 ( .Y(n6914), .A0(n6895), .A1(n6897) );
  inv01 U4130 ( .Y(n6915), .A(n6914) );
  nand02 U4131 ( .Y(n6916), .A0(n6913), .A1(n6915) );
  inv01 U4132 ( .Y(n6877), .A(n6916) );
  inv02 U4133 ( .Y(n7835), .A(n7579) );
  inv04 U4134 ( .Y(n7760), .A(n6917) );
  inv01 U4135 ( .Y(n6918), .A(opa_i[18]) );
  inv01 U4136 ( .Y(n6919), .A(opa_i[19]) );
  inv01 U4137 ( .Y(n6920), .A(opa_i[17]) );
  nand02 U4138 ( .Y(n6917), .A0(n6920), .A1(n6921) );
  nand02 U4139 ( .Y(n6922), .A0(n6918), .A1(n6919) );
  inv01 U4140 ( .Y(n6921), .A(n6922) );
  inv01 U4141 ( .Y(n7937), .A(n6923) );
  nor02 U4142 ( .Y(n6924), .A0(n7892), .A1(n6925) );
  nor02 U4143 ( .Y(n6926), .A0(n7892), .A1(n6927) );
  nor02 U4144 ( .Y(n6928), .A0(n7892), .A1(n6929) );
  nor02 U4145 ( .Y(n6930), .A0(n7892), .A1(n6931) );
  nor02 U4146 ( .Y(n6932), .A0(n7668), .A1(n6933) );
  nor02 U4147 ( .Y(n6934), .A0(n7668), .A1(n6935) );
  nor02 U4148 ( .Y(n6936), .A0(n7668), .A1(n6937) );
  nor02 U4149 ( .Y(n6938), .A0(n7668), .A1(n6939) );
  nor02 U4150 ( .Y(n6923), .A0(n6940), .A1(n6941) );
  nor02 U4151 ( .Y(n6942), .A0(n7938), .A1(n7897) );
  inv01 U4152 ( .Y(n6925), .A(n6942) );
  nor02 U4153 ( .Y(n6943), .A0(n7674), .A1(n7897) );
  inv01 U4154 ( .Y(n6927), .A(n6943) );
  nor02 U4155 ( .Y(n6944), .A0(n7938), .A1(n7676) );
  inv01 U4156 ( .Y(n6929), .A(n6944) );
  nor02 U4157 ( .Y(n6945), .A0(n7674), .A1(n7676) );
  inv01 U4158 ( .Y(n6931), .A(n6945) );
  nor02 U4159 ( .Y(n6946), .A0(n7938), .A1(n7897) );
  inv01 U4160 ( .Y(n6933), .A(n6946) );
  nor02 U4161 ( .Y(n6947), .A0(n7674), .A1(n7897) );
  inv01 U4162 ( .Y(n6935), .A(n6947) );
  nor02 U4163 ( .Y(n6948), .A0(n7938), .A1(n7676) );
  inv01 U4164 ( .Y(n6937), .A(n6948) );
  nor02 U4165 ( .Y(n6949), .A0(n7674), .A1(n7676) );
  inv01 U4166 ( .Y(n6939), .A(n6949) );
  nor02 U4167 ( .Y(n6950), .A0(n6924), .A1(n6926) );
  inv01 U4168 ( .Y(n6951), .A(n6950) );
  nor02 U4169 ( .Y(n6952), .A0(n6928), .A1(n6930) );
  inv01 U4170 ( .Y(n6953), .A(n6952) );
  nor02 U4171 ( .Y(n6954), .A0(n6951), .A1(n6953) );
  inv01 U4172 ( .Y(n6940), .A(n6954) );
  nor02 U4173 ( .Y(n6955), .A0(n6932), .A1(n6934) );
  inv01 U4174 ( .Y(n6956), .A(n6955) );
  nor02 U4175 ( .Y(n6957), .A0(n6936), .A1(n6938) );
  inv01 U4176 ( .Y(n6958), .A(n6957) );
  nor02 U4177 ( .Y(n6959), .A0(n6956), .A1(n6958) );
  inv01 U4178 ( .Y(n6941), .A(n6959) );
  buf08 U4179 ( .Y(n7676), .A(n7847) );
  buf04 U4180 ( .Y(n7668), .A(n7896) );
  inv02 U4181 ( .Y(n8048), .A(n6960) );
  inv01 U4182 ( .Y(n6961), .A(exp_i[1]) );
  inv01 U4183 ( .Y(n6962), .A(fract_28_i[27]) );
  inv08 U4184 ( .Y(n6963), .A(exp_i[0]) );
  nor02 U4185 ( .Y(n6960), .A0(n6963), .A1(n6964) );
  nor02 U4186 ( .Y(n6965), .A0(n6961), .A1(n6962) );
  inv01 U4187 ( .Y(n6964), .A(n6965) );
  buf02 U4188 ( .Y(n6966), .A(n8103) );
  buf02 U4189 ( .Y(n6967), .A(n8103) );
  or02 U4190 ( .Y(n6968), .A0(n4780), .A1(n8024) );
  inv02 U4191 ( .Y(n6969), .A(n6968) );
  inv02 U4192 ( .Y(n8104), .A(n6970) );
  nand02 U4193 ( .Y(n6970), .A0(n4513), .A1(n6971) );
  nand02 U4194 ( .Y(n6972), .A0(n7882), .A1(n7954) );
  inv01 U4195 ( .Y(n6971), .A(n6972) );
  inv02 U4196 ( .Y(n8105), .A(n6973) );
  nand02 U4197 ( .Y(n6973), .A0(n4746), .A1(n6974) );
  nand02 U4198 ( .Y(n6975), .A0(n7961), .A1(n7949) );
  inv01 U4199 ( .Y(n6974), .A(n6975) );
  or04 U4200 ( .Y(n6976), .A0(n7745), .A1(n7747), .A2(n7749), .A3(n7324) );
  inv01 U4201 ( .Y(n6977), .A(n6976) );
  or04 U4202 ( .Y(n6978), .A0(n7803), .A1(n7740), .A2(n7744), .A3(n7742) );
  inv01 U4203 ( .Y(n6979), .A(n6978) );
  inv02 U4204 ( .Y(n8030), .A(n6980) );
  nor02 U4205 ( .Y(n6981), .A0(n7707), .A1(n7387) );
  inv01 U4206 ( .Y(n6982), .A(n8045) );
  nor02 U4207 ( .Y(n6980), .A0(n6981), .A1(n6982) );
  inv01 U4208 ( .Y(n7765), .A(n6983) );
  inv01 U4209 ( .Y(n6984), .A(opb_i[0]) );
  inv01 U4210 ( .Y(n6985), .A(opb_i[10]) );
  inv01 U4211 ( .Y(n6986), .A(n7772) );
  inv01 U4212 ( .Y(n6987), .A(opb_i[11]) );
  nand02 U4213 ( .Y(n6983), .A0(n6988), .A1(n6989) );
  nand02 U4214 ( .Y(n6990), .A0(n6984), .A1(n6985) );
  inv01 U4215 ( .Y(n6988), .A(n6990) );
  nand02 U4216 ( .Y(n6991), .A0(n6986), .A1(n6987) );
  inv01 U4217 ( .Y(n6989), .A(n6991) );
  nand02 U4218 ( .Y(n7743), .A0(n6992), .A1(n6993) );
  inv01 U4219 ( .Y(n6994), .A(n____return2548_4_) );
  inv01 U4220 ( .Y(n6995), .A(s_expo9_1[4]) );
  inv01 U4221 ( .Y(n6996), .A(n7667) );
  nand02 U4222 ( .Y(n6992), .A0(n7667), .A1(n6994) );
  nand02 U4223 ( .Y(n6993), .A0(n6995), .A1(n6996) );
  nand02 U4224 ( .Y(n7741), .A0(n6997), .A1(n6998) );
  inv01 U4225 ( .Y(n6999), .A(n____return2548_5_) );
  inv01 U4226 ( .Y(n7000), .A(s_expo9_1[5]) );
  inv01 U4227 ( .Y(n7001), .A(n7667) );
  nand02 U4228 ( .Y(n6997), .A0(n7667), .A1(n6999) );
  nand02 U4229 ( .Y(n6998), .A0(n7000), .A1(n7001) );
  inv01 U4230 ( .Y(n8110), .A(n7002) );
  inv01 U4231 ( .Y(n7003), .A(n7316) );
  inv01 U4232 ( .Y(n7004), .A(n8078) );
  inv01 U4233 ( .Y(n7005), .A(n8077) );
  inv01 U4234 ( .Y(n7006), .A(n8082) );
  nand02 U4235 ( .Y(n7002), .A0(n7007), .A1(n7008) );
  nand02 U4236 ( .Y(n7009), .A0(n7003), .A1(n7004) );
  inv01 U4237 ( .Y(n7007), .A(n7009) );
  nand02 U4238 ( .Y(n7010), .A0(n7005), .A1(n7006) );
  inv01 U4239 ( .Y(n7008), .A(n7010) );
  buf02 U4240 ( .Y(n7011), .A(n7681) );
  buf02 U4241 ( .Y(n7012), .A(n7685) );
  inv08 U4242 ( .Y(n7716), .A(n7011) );
  inv08 U4243 ( .Y(n7713), .A(n7012) );
  nand02 U4244 ( .Y(s_output_o[31]), .A0(n7013), .A1(n7014) );
  inv01 U4245 ( .Y(n7015), .A(n7726) );
  inv01 U4246 ( .Y(n7016), .A(n7725) );
  inv01 U4247 ( .Y(n7017), .A(n7724) );
  inv01 U4248 ( .Y(n7018), .A(n7728) );
  inv01 U4249 ( .Y(n7019), .A(n7727) );
  nand02 U4250 ( .Y(n7013), .A0(n7017), .A1(n7020) );
  nand02 U4251 ( .Y(n7014), .A0(n7018), .A1(n7019) );
  nand02 U4252 ( .Y(n7021), .A0(n7015), .A1(n7016) );
  inv01 U4253 ( .Y(n7020), .A(n7021) );
  inv02 U4254 ( .Y(n7728), .A(sign_i) );
  inv01 U4255 ( .Y(n8112), .A(n7022) );
  inv01 U4256 ( .Y(n7023), .A(n8063) );
  inv01 U4257 ( .Y(n7024), .A(n8065) );
  inv01 U4258 ( .Y(n7025), .A(n8064) );
  inv01 U4259 ( .Y(n7026), .A(n8067) );
  nand02 U4260 ( .Y(n7022), .A0(n7027), .A1(n7028) );
  nand02 U4261 ( .Y(n7029), .A0(n7023), .A1(n7024) );
  inv01 U4262 ( .Y(n7027), .A(n7029) );
  nand02 U4263 ( .Y(n7030), .A0(n7025), .A1(n7026) );
  inv01 U4264 ( .Y(n7028), .A(n7030) );
  inv01 U4265 ( .Y(n7766), .A(n7031) );
  inv01 U4266 ( .Y(n7032), .A(opb_i[18]) );
  inv01 U4267 ( .Y(n7033), .A(opb_i[16]) );
  inv01 U4268 ( .Y(n7034), .A(opb_i[19]) );
  inv01 U4269 ( .Y(n7035), .A(n7771) );
  nand02 U4270 ( .Y(n7031), .A0(n7036), .A1(n7037) );
  nand02 U4271 ( .Y(n7038), .A0(n7032), .A1(n7033) );
  inv01 U4272 ( .Y(n7036), .A(n7038) );
  nand02 U4273 ( .Y(n7039), .A0(n7034), .A1(n7035) );
  inv01 U4274 ( .Y(n7037), .A(n7039) );
  inv01 U4275 ( .Y(n7767), .A(n7040) );
  inv01 U4276 ( .Y(n7041), .A(opb_i[20]) );
  inv01 U4277 ( .Y(n7042), .A(opb_i[2]) );
  inv01 U4278 ( .Y(n7043), .A(opb_i[1]) );
  inv01 U4279 ( .Y(n7044), .A(n7770) );
  nand02 U4280 ( .Y(n7040), .A0(n7045), .A1(n7046) );
  nand02 U4281 ( .Y(n7047), .A0(n7041), .A1(n7042) );
  inv01 U4282 ( .Y(n7045), .A(n7047) );
  nand02 U4283 ( .Y(n7048), .A0(n7043), .A1(n7044) );
  inv01 U4284 ( .Y(n7046), .A(n7048) );
  nand02 U4285 ( .Y(n8088), .A0(n7049), .A1(n7050) );
  inv02 U4286 ( .Y(n7051), .A(n7316) );
  inv02 U4287 ( .Y(n7052), .A(n8089) );
  inv01 U4288 ( .Y(n7053), .A(n7428) );
  inv01 U4289 ( .Y(n7054), .A(fract_28_i[22]) );
  inv01 U4290 ( .Y(n7055), .A(n6660) );
  inv01 U4291 ( .Y(n7056), .A(n8072) );
  nand02 U4292 ( .Y(n7057), .A0(n7053), .A1(n7058) );
  nand02 U4293 ( .Y(n7059), .A0(n7054), .A1(n7060) );
  nand02 U4294 ( .Y(n7061), .A0(n7055), .A1(n7062) );
  nand02 U4295 ( .Y(n7063), .A0(n7056), .A1(n7064) );
  nand02 U4296 ( .Y(n7065), .A0(n7056), .A1(n7066) );
  nand02 U4297 ( .Y(n7067), .A0(n7056), .A1(n7068) );
  nand02 U4298 ( .Y(n7069), .A0(n7051), .A1(n7052) );
  inv01 U4299 ( .Y(n7058), .A(n7069) );
  nand02 U4300 ( .Y(n7070), .A0(n7051), .A1(n7052) );
  inv01 U4301 ( .Y(n7060), .A(n7070) );
  nand02 U4302 ( .Y(n7071), .A0(n7051), .A1(n7052) );
  inv01 U4303 ( .Y(n7062), .A(n7071) );
  nand02 U4304 ( .Y(n7072), .A0(n7051), .A1(n7053) );
  inv01 U4305 ( .Y(n7064), .A(n7072) );
  nand02 U4306 ( .Y(n7073), .A0(n7051), .A1(n7054) );
  inv01 U4307 ( .Y(n7066), .A(n7073) );
  nand02 U4308 ( .Y(n7074), .A0(n7051), .A1(n7055) );
  inv01 U4309 ( .Y(n7068), .A(n7074) );
  nand02 U4310 ( .Y(n7075), .A0(n7057), .A1(n7059) );
  inv01 U4311 ( .Y(n7076), .A(n7075) );
  nand02 U4312 ( .Y(n7077), .A0(n7061), .A1(n7076) );
  inv01 U4313 ( .Y(n7049), .A(n7077) );
  nand02 U4314 ( .Y(n7078), .A0(n7063), .A1(n7065) );
  inv01 U4315 ( .Y(n7079), .A(n7078) );
  nand02 U4316 ( .Y(n7080), .A0(n7067), .A1(n7079) );
  inv01 U4317 ( .Y(n7050), .A(n7080) );
  xor2 U4318 ( .Y(n7081), .A0(exp_i[3]), .A1(n4649) );
  inv02 U4319 ( .Y(n7082), .A(n7081) );
  nand02 U4320 ( .Y(n8109), .A0(n7083), .A1(n7084) );
  inv02 U4321 ( .Y(n7085), .A(n8072) );
  inv02 U4322 ( .Y(n7086), .A(n7900) );
  inv02 U4323 ( .Y(n7087), .A(fract_28_i[23]) );
  inv02 U4324 ( .Y(n7088), .A(n7911) );
  inv02 U4325 ( .Y(n7089), .A(n7429) );
  inv02 U4326 ( .Y(n7090), .A(fract_28_i[25]) );
  inv02 U4327 ( .Y(n7091), .A(fract_28_i[21]) );
  nand02 U4328 ( .Y(n7092), .A0(n7087), .A1(n7093) );
  nand02 U4329 ( .Y(n7094), .A0(n7088), .A1(n7095) );
  nand02 U4330 ( .Y(n7096), .A0(n7089), .A1(n7097) );
  nand02 U4331 ( .Y(n7098), .A0(n7090), .A1(n7099) );
  nand02 U4332 ( .Y(n7100), .A0(n7090), .A1(n7101) );
  nand02 U4333 ( .Y(n7102), .A0(n7090), .A1(n7103) );
  nand02 U4334 ( .Y(n7104), .A0(n7091), .A1(n7105) );
  nand02 U4335 ( .Y(n7106), .A0(n7091), .A1(n7107) );
  nand02 U4336 ( .Y(n7108), .A0(n7091), .A1(n7109) );
  nand02 U4337 ( .Y(n7110), .A0(n7091), .A1(n7111) );
  nand02 U4338 ( .Y(n7112), .A0(n7091), .A1(n7113) );
  nand02 U4339 ( .Y(n7114), .A0(n7091), .A1(n7115) );
  nand02 U4340 ( .Y(n7116), .A0(n7085), .A1(n7086) );
  inv01 U4341 ( .Y(n7093), .A(n7116) );
  nand02 U4342 ( .Y(n7117), .A0(n7085), .A1(n7086) );
  inv01 U4343 ( .Y(n7095), .A(n7117) );
  nand02 U4344 ( .Y(n7118), .A0(n7085), .A1(n7086) );
  inv01 U4345 ( .Y(n7097), .A(n7118) );
  nand02 U4346 ( .Y(n7119), .A0(n7085), .A1(n7087) );
  inv01 U4347 ( .Y(n7099), .A(n7119) );
  nand02 U4348 ( .Y(n7120), .A0(n7085), .A1(n7088) );
  inv01 U4349 ( .Y(n7101), .A(n7120) );
  nand02 U4350 ( .Y(n7121), .A0(n7085), .A1(n7089) );
  inv01 U4351 ( .Y(n7103), .A(n7121) );
  nand02 U4352 ( .Y(n7122), .A0(n7086), .A1(n7087) );
  inv01 U4353 ( .Y(n7105), .A(n7122) );
  nand02 U4354 ( .Y(n7123), .A0(n7086), .A1(n7088) );
  inv01 U4355 ( .Y(n7107), .A(n7123) );
  nand02 U4356 ( .Y(n7124), .A0(n7086), .A1(n7089) );
  inv01 U4357 ( .Y(n7109), .A(n7124) );
  nand02 U4358 ( .Y(n7125), .A0(n7087), .A1(n7090) );
  inv01 U4359 ( .Y(n7111), .A(n7125) );
  nand02 U4360 ( .Y(n7126), .A0(n7088), .A1(n7090) );
  inv01 U4361 ( .Y(n7113), .A(n7126) );
  nand02 U4362 ( .Y(n7127), .A0(n7089), .A1(n7090) );
  inv01 U4363 ( .Y(n7115), .A(n7127) );
  nand02 U4364 ( .Y(n7128), .A0(n7092), .A1(n7094) );
  inv01 U4365 ( .Y(n7129), .A(n7128) );
  nand02 U4366 ( .Y(n7130), .A0(n7096), .A1(n7129) );
  inv01 U4367 ( .Y(n7131), .A(n7130) );
  nand02 U4368 ( .Y(n7132), .A0(n7098), .A1(n7100) );
  inv01 U4369 ( .Y(n7133), .A(n7132) );
  nand02 U4370 ( .Y(n7134), .A0(n7102), .A1(n7133) );
  inv01 U4371 ( .Y(n7135), .A(n7134) );
  nand02 U4372 ( .Y(n7136), .A0(n7131), .A1(n7135) );
  inv01 U4373 ( .Y(n7083), .A(n7136) );
  nand02 U4374 ( .Y(n7137), .A0(n7104), .A1(n7106) );
  inv01 U4375 ( .Y(n7138), .A(n7137) );
  nand02 U4376 ( .Y(n7139), .A0(n7108), .A1(n7138) );
  inv01 U4377 ( .Y(n7140), .A(n7139) );
  nand02 U4378 ( .Y(n7141), .A0(n7110), .A1(n7112) );
  inv01 U4379 ( .Y(n7142), .A(n7141) );
  nand02 U4380 ( .Y(n7143), .A0(n7114), .A1(n7142) );
  inv01 U4381 ( .Y(n7144), .A(n7143) );
  nand02 U4382 ( .Y(n7145), .A0(n7140), .A1(n7144) );
  inv01 U4383 ( .Y(n7084), .A(n7145) );
  nand02 U4384 ( .Y(n8071), .A0(n7146), .A1(n7147) );
  inv02 U4385 ( .Y(n7148), .A(n7316) );
  inv02 U4386 ( .Y(n7149), .A(n8074) );
  inv01 U4387 ( .Y(n7150), .A(n8072) );
  inv01 U4388 ( .Y(n7151), .A(fract_28_i[20]) );
  inv01 U4389 ( .Y(n7152), .A(n7604) );
  inv01 U4390 ( .Y(n7153), .A(n7428) );
  nand02 U4391 ( .Y(n7154), .A0(n7150), .A1(n7155) );
  nand02 U4392 ( .Y(n7156), .A0(n7151), .A1(n7157) );
  nand02 U4393 ( .Y(n7158), .A0(n7152), .A1(n7159) );
  nand02 U4394 ( .Y(n7160), .A0(n7153), .A1(n7161) );
  nand02 U4395 ( .Y(n7162), .A0(n7153), .A1(n7163) );
  nand02 U4396 ( .Y(n7164), .A0(n7153), .A1(n7165) );
  nand02 U4397 ( .Y(n7166), .A0(n7148), .A1(n7149) );
  inv01 U4398 ( .Y(n7155), .A(n7166) );
  nand02 U4399 ( .Y(n7167), .A0(n7148), .A1(n7149) );
  inv01 U4400 ( .Y(n7157), .A(n7167) );
  nand02 U4401 ( .Y(n7168), .A0(n7148), .A1(n7149) );
  inv01 U4402 ( .Y(n7159), .A(n7168) );
  nand02 U4403 ( .Y(n7169), .A0(n7148), .A1(n7150) );
  inv01 U4404 ( .Y(n7161), .A(n7169) );
  nand02 U4405 ( .Y(n7170), .A0(n7148), .A1(n7151) );
  inv01 U4406 ( .Y(n7163), .A(n7170) );
  nand02 U4407 ( .Y(n7171), .A0(n7148), .A1(n7152) );
  inv01 U4408 ( .Y(n7165), .A(n7171) );
  nand02 U4409 ( .Y(n7172), .A0(n7154), .A1(n7156) );
  inv01 U4410 ( .Y(n7173), .A(n7172) );
  nand02 U4411 ( .Y(n7174), .A0(n7158), .A1(n7173) );
  inv01 U4412 ( .Y(n7146), .A(n7174) );
  nand02 U4413 ( .Y(n7175), .A0(n7160), .A1(n7162) );
  inv01 U4414 ( .Y(n7176), .A(n7175) );
  nand02 U4415 ( .Y(n7177), .A0(n7164), .A1(n7176) );
  inv01 U4416 ( .Y(n7147), .A(n7177) );
  inv01 U4417 ( .Y(n7768), .A(n7178) );
  inv01 U4418 ( .Y(n7179), .A(opb_i[5]) );
  inv01 U4419 ( .Y(n7180), .A(opb_i[6]) );
  inv01 U4420 ( .Y(n7181), .A(opb_i[4]) );
  inv01 U4421 ( .Y(n7182), .A(n7769) );
  nand02 U4422 ( .Y(n7178), .A0(n7183), .A1(n7184) );
  nand02 U4423 ( .Y(n7185), .A0(n7179), .A1(n7180) );
  inv01 U4424 ( .Y(n7183), .A(n7185) );
  nand02 U4425 ( .Y(n7186), .A0(n7181), .A1(n7182) );
  inv01 U4426 ( .Y(n7184), .A(n7186) );
  or02 U4427 ( .Y(n7187), .A0(n8030), .A1(n8041) );
  inv02 U4428 ( .Y(n7188), .A(n7187) );
  xor2 U4429 ( .Y(n7189), .A0(n8040), .A1(exp_i[6]) );
  inv02 U4430 ( .Y(n7190), .A(n7189) );
  buf02 U4431 ( .Y(n7191), .A(n4247) );
  nand02 U4432 ( .Y(n7802), .A0(n7192), .A1(n7193) );
  inv02 U4433 ( .Y(n7194), .A(n6977) );
  inv02 U4434 ( .Y(n7195), .A(n6979) );
  inv02 U4435 ( .Y(n7196), .A(n4714) );
  inv02 U4436 ( .Y(n7197), .A(n____return2864_1_) );
  inv02 U4437 ( .Y(n7198), .A(n____return2864_2_) );
  inv02 U4438 ( .Y(n7199), .A(n4710) );
  inv02 U4439 ( .Y(n7200), .A(s_expo9_2[5]) );
  inv02 U4440 ( .Y(n7201), .A(s_expo9_2[4]) );
  nand02 U4441 ( .Y(n7202), .A0(n7194), .A1(n7195) );
  nand02 U4442 ( .Y(n7203), .A0(n7194), .A1(n7196) );
  nand02 U4443 ( .Y(n7204), .A0(n7194), .A1(n7197) );
  nand02 U4444 ( .Y(n7205), .A0(n7194), .A1(n7198) );
  nand02 U4445 ( .Y(n7206), .A0(n7195), .A1(n7199) );
  nand02 U4446 ( .Y(n7207), .A0(n7196), .A1(n7199) );
  nand02 U4447 ( .Y(n7208), .A0(n7197), .A1(n7199) );
  nand02 U4448 ( .Y(n7209), .A0(n7198), .A1(n7199) );
  nand02 U4449 ( .Y(n7210), .A0(n7195), .A1(n7200) );
  nand02 U4450 ( .Y(n7211), .A0(n7196), .A1(n7200) );
  nand02 U4451 ( .Y(n7212), .A0(n7197), .A1(n7200) );
  nand02 U4452 ( .Y(n7213), .A0(n7198), .A1(n7200) );
  nand02 U4453 ( .Y(n7214), .A0(n7195), .A1(n7201) );
  nand02 U4454 ( .Y(n7215), .A0(n7196), .A1(n7201) );
  nand02 U4455 ( .Y(n7216), .A0(n7197), .A1(n7201) );
  nand02 U4456 ( .Y(n7217), .A0(n7198), .A1(n7201) );
  nand02 U4457 ( .Y(n7218), .A0(n7202), .A1(n7203) );
  inv01 U4458 ( .Y(n7219), .A(n7218) );
  nand02 U4459 ( .Y(n7220), .A0(n7204), .A1(n7205) );
  inv01 U4460 ( .Y(n7221), .A(n7220) );
  nand02 U4461 ( .Y(n7222), .A0(n7219), .A1(n7221) );
  inv01 U4462 ( .Y(n7223), .A(n7222) );
  nand02 U4463 ( .Y(n7224), .A0(n7206), .A1(n7207) );
  inv01 U4464 ( .Y(n7225), .A(n7224) );
  nand02 U4465 ( .Y(n7226), .A0(n7208), .A1(n7209) );
  inv01 U4466 ( .Y(n7227), .A(n7226) );
  nand02 U4467 ( .Y(n7228), .A0(n7225), .A1(n7227) );
  inv01 U4468 ( .Y(n7229), .A(n7228) );
  nand02 U4469 ( .Y(n7230), .A0(n7223), .A1(n7229) );
  inv01 U4470 ( .Y(n7192), .A(n7230) );
  nand02 U4471 ( .Y(n7231), .A0(n7210), .A1(n7211) );
  inv01 U4472 ( .Y(n7232), .A(n7231) );
  nand02 U4473 ( .Y(n7233), .A0(n7212), .A1(n7213) );
  inv01 U4474 ( .Y(n7234), .A(n7233) );
  nand02 U4475 ( .Y(n7235), .A0(n7232), .A1(n7234) );
  inv01 U4476 ( .Y(n7236), .A(n7235) );
  nand02 U4477 ( .Y(n7237), .A0(n7214), .A1(n7215) );
  inv01 U4478 ( .Y(n7238), .A(n7237) );
  nand02 U4479 ( .Y(n7239), .A0(n7216), .A1(n7217) );
  inv01 U4480 ( .Y(n7240), .A(n7239) );
  nand02 U4481 ( .Y(n7241), .A0(n7238), .A1(n7240) );
  inv01 U4482 ( .Y(n7242), .A(n7241) );
  nand02 U4483 ( .Y(n7243), .A0(n7236), .A1(n7242) );
  inv01 U4484 ( .Y(n7193), .A(n7243) );
  inv02 U4485 ( .Y(s_expo9_2[4]), .A(n7743) );
  inv02 U4486 ( .Y(s_expo9_2[5]), .A(n7741) );
  or02 U4487 ( .Y(n7244), .A0(fract_28_i[21]), .A1(fract_28_i[20]) );
  inv02 U4488 ( .Y(n7245), .A(n7244) );
  inv01 U4489 ( .Y(n7916), .A(n7246) );
  nor02 U4490 ( .Y(n7247), .A0(n7947), .A1(n7703) );
  nor02 U4491 ( .Y(n7248), .A0(n7943), .A1(n7702) );
  inv01 U4492 ( .Y(n7249), .A(n4349) );
  nor02 U4493 ( .Y(n7246), .A0(n7249), .A1(n7250) );
  nor02 U4494 ( .Y(n7251), .A0(n7247), .A1(n7248) );
  inv01 U4495 ( .Y(n7250), .A(n7251) );
  inv01 U4496 ( .Y(n7853), .A(n7252) );
  nor02 U4497 ( .Y(n7253), .A0(n7873), .A1(n7698) );
  nor02 U4498 ( .Y(n7254), .A0(n7887), .A1(n7701) );
  inv01 U4499 ( .Y(n7255), .A(n7888) );
  nor02 U4500 ( .Y(n7252), .A0(n7255), .A1(n7256) );
  nor02 U4501 ( .Y(n7257), .A0(n7253), .A1(n7254) );
  inv01 U4502 ( .Y(n7256), .A(n7257) );
  inv01 U4503 ( .Y(n7899), .A(n7258) );
  nor02 U4504 ( .Y(n7259), .A0(n7941), .A1(n7703) );
  nor02 U4505 ( .Y(n7260), .A0(n7932), .A1(n7702) );
  inv01 U4506 ( .Y(n7261), .A(n4434) );
  nor02 U4507 ( .Y(n7258), .A0(n7261), .A1(n7262) );
  nor02 U4508 ( .Y(n7263), .A0(n7259), .A1(n7260) );
  inv01 U4509 ( .Y(n7262), .A(n7263) );
  inv01 U4510 ( .Y(n7868), .A(n7264) );
  nor02 U4511 ( .Y(n7265), .A0(n7954), .A1(n7700) );
  nor02 U4512 ( .Y(n7266), .A0(n7882), .A1(n7701) );
  inv01 U4513 ( .Y(n7267), .A(n8010) );
  nor02 U4514 ( .Y(n7264), .A0(n7267), .A1(n7268) );
  nor02 U4515 ( .Y(n7269), .A0(n7265), .A1(n7266) );
  inv01 U4516 ( .Y(n7268), .A(n7269) );
  inv01 U4517 ( .Y(n7860), .A(n7270) );
  nor02 U4518 ( .Y(n7271), .A0(n7887), .A1(n7700) );
  nor02 U4519 ( .Y(n7272), .A0(n7954), .A1(n7701) );
  inv01 U4520 ( .Y(n7273), .A(n4381) );
  nor02 U4521 ( .Y(n7270), .A0(n7273), .A1(n7274) );
  nor02 U4522 ( .Y(n7275), .A0(n7271), .A1(n7272) );
  inv01 U4523 ( .Y(n7274), .A(n7275) );
  inv02 U4524 ( .Y(n7954), .A(fract_28_i[7]) );
  inv01 U4525 ( .Y(n7910), .A(n7276) );
  nor02 U4526 ( .Y(n7277), .A0(n7943), .A1(n7703) );
  nor02 U4527 ( .Y(n7278), .A0(n7941), .A1(n7702) );
  inv01 U4528 ( .Y(n7279), .A(n4416) );
  nor02 U4529 ( .Y(n7276), .A0(n7279), .A1(n7280) );
  nor02 U4530 ( .Y(n7281), .A0(n7277), .A1(n7278) );
  inv01 U4531 ( .Y(n7280), .A(n7281) );
  nand02 U4532 ( .Y(n7282), .A0(n8007), .A1(n7311) );
  inv02 U4533 ( .Y(n7283), .A(n7282) );
  inv01 U4534 ( .Y(n7846), .A(n7284) );
  nor02 U4535 ( .Y(n7285), .A0(n7875), .A1(n7699) );
  nor02 U4536 ( .Y(n7286), .A0(n7873), .A1(n7701) );
  inv01 U4537 ( .Y(n7287), .A(n7877) );
  nor02 U4538 ( .Y(n7284), .A0(n7287), .A1(n7288) );
  nor02 U4539 ( .Y(n7289), .A0(n7285), .A1(n7286) );
  inv01 U4540 ( .Y(n7288), .A(n7289) );
  inv01 U4541 ( .Y(n7927), .A(n7290) );
  nor02 U4542 ( .Y(n7291), .A0(n7949), .A1(n7703) );
  nor02 U4543 ( .Y(n7292), .A0(n7947), .A1(n7702) );
  inv01 U4544 ( .Y(n7293), .A(n7950) );
  nor02 U4545 ( .Y(n7290), .A0(n7293), .A1(n7294) );
  nor02 U4546 ( .Y(n7295), .A0(n7291), .A1(n7292) );
  inv01 U4547 ( .Y(n7294), .A(n7295) );
  or02 U4548 ( .Y(n7296), .A0(n7988), .A1(n7704) );
  inv02 U4549 ( .Y(n7297), .A(n7296) );
  inv02 U4550 ( .Y(n8068), .A(n7298) );
  inv01 U4551 ( .Y(n7299), .A(n8081) );
  inv01 U4552 ( .Y(n7300), .A(n8080) );
  inv01 U4553 ( .Y(n7301), .A(n8082) );
  nand02 U4554 ( .Y(n7298), .A0(n7301), .A1(n7302) );
  nand02 U4555 ( .Y(n7303), .A0(n7299), .A1(n7300) );
  inv01 U4556 ( .Y(n7302), .A(n7303) );
  inv02 U4557 ( .Y(n7793), .A(n7304) );
  nor02 U4558 ( .Y(n7305), .A0(n8097), .A1(n8098) );
  inv01 U4559 ( .Y(n7306), .A(n7704) );
  nor02 U4560 ( .Y(n7304), .A0(n7305), .A1(n7306) );
  inv02 U4561 ( .Y(n8067), .A(n7307) );
  nand02 U4562 ( .Y(n7307), .A0(n4732), .A1(n7308) );
  nand02 U4563 ( .Y(n7309), .A0(n7804), .A1(n7986) );
  inv01 U4564 ( .Y(n7308), .A(n7309) );
  buf02 U4565 ( .Y(n7310), .A(n8008) );
  buf02 U4566 ( .Y(n7311), .A(n8008) );
  inv02 U4567 ( .Y(n8034), .A(n7312) );
  nor02 U4568 ( .Y(n7313), .A0(n8083), .A1(n8084) );
  inv01 U4569 ( .Y(n7314), .A(n7704) );
  nor02 U4570 ( .Y(n7312), .A0(n7313), .A1(n7314) );
  nand02 U4571 ( .Y(n7315), .A0(fract_28_i[3]), .A1(n6966) );
  inv02 U4572 ( .Y(n7316), .A(n7315) );
  inv02 U4573 ( .Y(n8040), .A(n7317) );
  nand02 U4574 ( .Y(n7317), .A0(exp_i[5]), .A1(n7318) );
  nand02 U4575 ( .Y(n7319), .A0(n8044), .A1(exp_i[4]) );
  inv01 U4576 ( .Y(n7318), .A(n7319) );
  inv02 U4577 ( .Y(n7734), .A(n7320) );
  inv01 U4578 ( .Y(n7321), .A(n7667) );
  nor02 U4579 ( .Y(n7322), .A0(n____return2548_7_), .A1(n7321) );
  nor02 U4580 ( .Y(n7323), .A0(n7667), .A1(s_expo9_1[7]) );
  nor02 U4581 ( .Y(n7320), .A0(n7322), .A1(n7323) );
  buf02 U4582 ( .Y(n7324), .A(n7751) );
  inv02 U4583 ( .Y(n7739), .A(n7325) );
  inv01 U4584 ( .Y(n7326), .A(n7667) );
  nor02 U4585 ( .Y(n7327), .A0(n____return2548_6_), .A1(n7326) );
  nor02 U4586 ( .Y(n7328), .A0(n7667), .A1(s_expo9_1[6]) );
  nor02 U4587 ( .Y(n7325), .A0(n7327), .A1(n7328) );
  inv02 U4588 ( .Y(n7747), .A(n7329) );
  inv01 U4589 ( .Y(n7330), .A(n7667) );
  nor02 U4590 ( .Y(n7331), .A0(n____return2548_2_), .A1(n7330) );
  nor02 U4591 ( .Y(n7332), .A0(n7667), .A1(s_expo9_1[2]) );
  nor02 U4592 ( .Y(n7329), .A0(n7331), .A1(n7332) );
  inv02 U4593 ( .Y(s_expo9_2[0]), .A(n7324) );
  nand02 U4594 ( .Y(n7712), .A0(n7333), .A1(n7334) );
  inv01 U4595 ( .Y(n7335), .A(n8026) );
  inv01 U4596 ( .Y(n7336), .A(n4780) );
  inv01 U4597 ( .Y(n7337), .A(n8024) );
  inv01 U4598 ( .Y(n7338), .A(n8025) );
  nand02 U4599 ( .Y(n7339), .A0(n7335), .A1(n7336) );
  nand02 U4600 ( .Y(n7340), .A0(n7335), .A1(n7337) );
  nand02 U4601 ( .Y(n7341), .A0(n7336), .A1(n7338) );
  nand02 U4602 ( .Y(n7342), .A0(n7337), .A1(n7338) );
  nand02 U4603 ( .Y(n7343), .A0(n7339), .A1(n7340) );
  inv01 U4604 ( .Y(n7333), .A(n7343) );
  nand02 U4605 ( .Y(n7344), .A0(n7341), .A1(n7342) );
  inv01 U4606 ( .Y(n7334), .A(n7344) );
  inv02 U4607 ( .Y(n7745), .A(n7345) );
  inv01 U4608 ( .Y(n7346), .A(n7667) );
  nor02 U4609 ( .Y(n7347), .A0(n____return2548_3_), .A1(n7346) );
  nor02 U4610 ( .Y(n7348), .A0(n7667), .A1(s_expo9_1[3]) );
  nor02 U4611 ( .Y(n7345), .A0(n7347), .A1(n7348) );
  inv02 U4612 ( .Y(n7749), .A(n7349) );
  inv01 U4613 ( .Y(n7350), .A(n7667) );
  nor02 U4614 ( .Y(n7351), .A0(n____return2548_1_), .A1(n7350) );
  nor02 U4615 ( .Y(n7352), .A0(n7667), .A1(s_expo9_1[1]) );
  nor02 U4616 ( .Y(n7349), .A0(n7351), .A1(n7352) );
  inv02 U4617 ( .Y(n7708), .A(n8034) );
  inv02 U4618 ( .Y(n7707), .A(n7793) );
  inv02 U4619 ( .Y(n8033), .A(n7353) );
  nor02 U4620 ( .Y(n7354), .A0(n7550), .A1(n7544) );
  inv01 U4621 ( .Y(n7355), .A(n8051) );
  nor02 U4622 ( .Y(n7353), .A0(n7354), .A1(n7355) );
  inv02 U4623 ( .Y(n7923), .A(n7356) );
  nor02 U4624 ( .Y(n7357), .A0(n7606), .A1(n7703) );
  nor02 U4625 ( .Y(n7358), .A0(n7967), .A1(n7702) );
  inv01 U4626 ( .Y(n7359), .A(n4383) );
  nor02 U4627 ( .Y(n7356), .A0(n7359), .A1(n7360) );
  nor02 U4628 ( .Y(n7361), .A0(n7357), .A1(n7358) );
  inv01 U4629 ( .Y(n7360), .A(n7361) );
  inv02 U4630 ( .Y(n7908), .A(n7362) );
  nor02 U4631 ( .Y(n7363), .A0(n7967), .A1(n7703) );
  nor02 U4632 ( .Y(n7364), .A0(n7961), .A1(n7702) );
  inv01 U4633 ( .Y(n7365), .A(n4299) );
  nor02 U4634 ( .Y(n7362), .A0(n7365), .A1(n7366) );
  nor02 U4635 ( .Y(n7367), .A0(n7363), .A1(n7364) );
  inv01 U4636 ( .Y(n7366), .A(n7367) );
  inv02 U4637 ( .Y(n7967), .A(fract_28_i[16]) );
  inv02 U4638 ( .Y(n7818), .A(n7368) );
  nor02 U4639 ( .Y(n7369), .A0(n7957), .A1(n7699) );
  nor02 U4640 ( .Y(n7370), .A0(n7956), .A1(n7701) );
  inv01 U4641 ( .Y(n7371), .A(n4414) );
  nor02 U4642 ( .Y(n7368), .A0(n7371), .A1(n7372) );
  nor02 U4643 ( .Y(n7373), .A0(n7369), .A1(n7370) );
  inv01 U4644 ( .Y(n7372), .A(n7373) );
  inv02 U4645 ( .Y(n7855), .A(n7374) );
  nor02 U4646 ( .Y(n7375), .A0(n7980), .A1(n7698) );
  nor02 U4647 ( .Y(n7376), .A0(n7957), .A1(n7701) );
  inv01 U4648 ( .Y(n7377), .A(n7999) );
  nor02 U4649 ( .Y(n7374), .A0(n7377), .A1(n7378) );
  nor02 U4650 ( .Y(n7379), .A0(n7375), .A1(n7376) );
  inv01 U4651 ( .Y(n7378), .A(n7379) );
  inv02 U4652 ( .Y(n7849), .A(n7380) );
  nor02 U4653 ( .Y(n7381), .A0(n7974), .A1(n7699) );
  nor02 U4654 ( .Y(n7382), .A0(n7980), .A1(n7701) );
  inv01 U4655 ( .Y(n7383), .A(n4387) );
  nor02 U4656 ( .Y(n7380), .A0(n7383), .A1(n7384) );
  nor02 U4657 ( .Y(n7385), .A0(n7381), .A1(n7382) );
  inv01 U4658 ( .Y(n7384), .A(n7385) );
  inv02 U4659 ( .Y(n7980), .A(fract_28_i[13]) );
  xor2 U4660 ( .Y(n7386), .A0(exp_i[4]), .A1(n8044) );
  inv02 U4661 ( .Y(n7387), .A(n7386) );
  inv02 U4662 ( .Y(n7934), .A(n7388) );
  nor02 U4663 ( .Y(n7389), .A0(n7974), .A1(n7703) );
  nor02 U4664 ( .Y(n7390), .A0(n7606), .A1(n7702) );
  inv01 U4665 ( .Y(n7391), .A(n7975) );
  nor02 U4666 ( .Y(n7388), .A0(n7391), .A1(n7392) );
  nor02 U4667 ( .Y(n7393), .A0(n7389), .A1(n7390) );
  inv01 U4668 ( .Y(n7392), .A(n7393) );
  inv02 U4669 ( .Y(n7830), .A(n7394) );
  nor02 U4670 ( .Y(n7395), .A0(n7956), .A1(n7699) );
  nor02 U4671 ( .Y(n7396), .A0(n7875), .A1(n7701) );
  inv01 U4672 ( .Y(n7397), .A(n4367) );
  nor02 U4673 ( .Y(n7394), .A0(n7397), .A1(n7398) );
  nor02 U4674 ( .Y(n7399), .A0(n7395), .A1(n7396) );
  inv01 U4675 ( .Y(n7398), .A(n7399) );
  inv02 U4676 ( .Y(n7897), .A(n7400) );
  nor02 U4677 ( .Y(n7401), .A0(n7961), .A1(n7703) );
  nor02 U4678 ( .Y(n7402), .A0(n7949), .A1(n7702) );
  inv01 U4679 ( .Y(n7403), .A(n4391) );
  nor02 U4680 ( .Y(n7400), .A0(n7403), .A1(n7404) );
  nor02 U4681 ( .Y(n7405), .A0(n7401), .A1(n7402) );
  inv01 U4682 ( .Y(n7404), .A(n7405) );
  inv02 U4683 ( .Y(n7875), .A(fract_28_i[10]) );
  inv02 U4684 ( .Y(n7949), .A(fract_28_i[18]) );
  inv02 U4685 ( .Y(n7963), .A(n7406) );
  nor02 U4686 ( .Y(n7407), .A0(n7900), .A1(n7700) );
  nor02 U4687 ( .Y(n7408), .A0(n7902), .A1(n7701) );
  inv01 U4688 ( .Y(n7409), .A(n7995) );
  nor02 U4689 ( .Y(n7406), .A0(n7409), .A1(n7410) );
  nor02 U4690 ( .Y(n7411), .A0(n7407), .A1(n7408) );
  inv01 U4691 ( .Y(n7410), .A(n7411) );
  inv02 U4692 ( .Y(n7900), .A(fract_28_i[26]) );
  or02 U4693 ( .Y(n7412), .A0(n7799), .A1(n7800) );
  inv02 U4694 ( .Y(n7413), .A(n7412) );
  inv02 U4695 ( .Y(n7930), .A(n7414) );
  nor02 U4696 ( .Y(n7415), .A0(n7955), .A1(n7703) );
  nor02 U4697 ( .Y(n7416), .A0(n7889), .A1(n7702) );
  inv01 U4698 ( .Y(n7417), .A(n4249) );
  nor02 U4699 ( .Y(n7414), .A0(n7417), .A1(n7418) );
  nor02 U4700 ( .Y(n7419), .A0(n7415), .A1(n7416) );
  inv01 U4701 ( .Y(n7418), .A(n7419) );
  inv02 U4702 ( .Y(n7955), .A(fract_28_i[2]) );
  or02 U4703 ( .Y(n7420), .A0(n7805), .A1(s_shr1_1_) );
  inv02 U4704 ( .Y(n7421), .A(n7420) );
  inv01 U4705 ( .Y(n7422), .A(n7420) );
  inv02 U4706 ( .Y(n7725), .A(n7423) );
  nor02 U4707 ( .Y(n7424), .A0(n7755), .A1(n7730) );
  nor02 U4708 ( .Y(n7425), .A0(n7427), .A1(n7730) );
  nor02 U4709 ( .Y(n7423), .A0(n7424), .A1(n7425) );
  inv02 U4710 ( .Y(n7730), .A(n7731) );
  or02 U4711 ( .Y(n7426), .A0(n7797), .A1(n7798) );
  inv02 U4712 ( .Y(n7427), .A(n7426) );
  buf02 U4713 ( .Y(n7428), .A(n8073) );
  buf02 U4714 ( .Y(n7429), .A(n8073) );
  or02 U4715 ( .Y(n7430), .A0(n7987), .A1(n7804) );
  inv02 U4716 ( .Y(n7431), .A(n7430) );
  nor02 U4717 ( .Y(n7433), .A0(n7887), .A1(n7703) );
  nor02 U4718 ( .Y(n7434), .A0(n7873), .A1(n7702) );
  inv01 U4719 ( .Y(n7435), .A(n4313) );
  nor02 U4720 ( .Y(n7432), .A0(n7435), .A1(n7436) );
  nor02 U4721 ( .Y(n7437), .A0(n7433), .A1(n7434) );
  inv02 U4722 ( .Y(n7436), .A(n7437) );
  inv02 U4723 ( .Y(n7887), .A(fract_28_i[8]) );
  nor02 U4724 ( .Y(n7439), .A0(n7941), .A1(n7698) );
  nor02 U4725 ( .Y(n7440), .A0(n7540), .A1(n7701) );
  inv01 U4726 ( .Y(n7441), .A(n4347) );
  nor02 U4727 ( .Y(n7438), .A0(n7441), .A1(n7442) );
  nor02 U4728 ( .Y(n7443), .A0(n7439), .A1(n7440) );
  inv02 U4729 ( .Y(n7442), .A(n7443) );
  nor02 U4730 ( .Y(n7445), .A0(n7882), .A1(n7703) );
  nor02 U4731 ( .Y(n7446), .A0(n7954), .A1(n7702) );
  inv01 U4732 ( .Y(n7447), .A(n4389) );
  nor02 U4733 ( .Y(n7444), .A0(n7447), .A1(n7448) );
  nor02 U4734 ( .Y(n7449), .A0(n7445), .A1(n7446) );
  inv02 U4735 ( .Y(n7448), .A(n7449) );
  nor02 U4736 ( .Y(n7451), .A0(n7943), .A1(n7698) );
  nor02 U4737 ( .Y(n7452), .A0(n7947), .A1(n7701) );
  inv01 U4738 ( .Y(n7453), .A(n4450) );
  nor02 U4739 ( .Y(n7450), .A0(n7453), .A1(n7454) );
  nor02 U4740 ( .Y(n7455), .A0(n7451), .A1(n7452) );
  inv02 U4741 ( .Y(n7454), .A(n7455) );
  inv02 U4742 ( .Y(n8038), .A(n7456) );
  nor02 U4743 ( .Y(n7457), .A0(n8033), .A1(n8049) );
  nor02 U4744 ( .Y(n7458), .A0(n8034), .A1(n8049) );
  nor02 U4745 ( .Y(n7456), .A0(n7457), .A1(n7458) );
  nor02 U4746 ( .Y(n7460), .A0(n7954), .A1(n7703) );
  nor02 U4747 ( .Y(n7461), .A0(n7887), .A1(n7702) );
  inv01 U4748 ( .Y(n7462), .A(n4410) );
  nor02 U4749 ( .Y(n7459), .A0(n7462), .A1(n7463) );
  nor02 U4750 ( .Y(n7464), .A0(n7460), .A1(n7461) );
  inv02 U4751 ( .Y(n7463), .A(n7464) );
  inv02 U4752 ( .Y(n7892), .A(n7465) );
  nor02 U4753 ( .Y(n7466), .A0(n7980), .A1(n7703) );
  nor02 U4754 ( .Y(n7467), .A0(n7974), .A1(n7702) );
  inv01 U4755 ( .Y(n7468), .A(n4418) );
  nor02 U4756 ( .Y(n7465), .A0(n7468), .A1(n7469) );
  nor02 U4757 ( .Y(n7470), .A0(n7466), .A1(n7467) );
  inv01 U4758 ( .Y(n7469), .A(n7470) );
  inv02 U4759 ( .Y(n7974), .A(fract_28_i[14]) );
  nor02 U4760 ( .Y(n7472), .A0(n7956), .A1(n7703) );
  nor02 U4761 ( .Y(n7473), .A0(n7957), .A1(n7702) );
  inv01 U4762 ( .Y(n7474), .A(n4363) );
  nor02 U4763 ( .Y(n7471), .A0(n7474), .A1(n7475) );
  nor02 U4764 ( .Y(n7476), .A0(n7472), .A1(n7473) );
  inv02 U4765 ( .Y(n7475), .A(n7476) );
  inv02 U4766 ( .Y(n7956), .A(fract_28_i[11]) );
  inv02 U4767 ( .Y(n7823), .A(n7477) );
  nor02 U4768 ( .Y(n7478), .A0(n7967), .A1(n7700) );
  nor02 U4769 ( .Y(n7479), .A0(n7606), .A1(n7701) );
  inv01 U4770 ( .Y(n7480), .A(n4345) );
  nor02 U4771 ( .Y(n7477), .A0(n7480), .A1(n7481) );
  nor02 U4772 ( .Y(n7482), .A0(n7478), .A1(n7479) );
  inv01 U4773 ( .Y(n7481), .A(n7482) );
  nor02 U4774 ( .Y(n7484), .A0(n7607), .A1(n7700) );
  nor02 U4775 ( .Y(n7485), .A0(n7967), .A1(n7701) );
  inv01 U4776 ( .Y(n7486), .A(n4315) );
  nor02 U4777 ( .Y(n7483), .A0(n7486), .A1(n7487) );
  nor02 U4778 ( .Y(n7488), .A0(n7484), .A1(n7485) );
  inv02 U4779 ( .Y(n7487), .A(n7488) );
  inv02 U4780 ( .Y(n7913), .A(n7489) );
  nor02 U4781 ( .Y(n7490), .A0(n7957), .A1(n7703) );
  nor02 U4782 ( .Y(n7491), .A0(n7980), .A1(n7702) );
  inv01 U4783 ( .Y(n7492), .A(n7983) );
  nor02 U4784 ( .Y(n7489), .A0(n7492), .A1(n7493) );
  nor02 U4785 ( .Y(n7494), .A0(n7490), .A1(n7491) );
  inv01 U4786 ( .Y(n7493), .A(n7494) );
  inv02 U4787 ( .Y(n7957), .A(fract_28_i[12]) );
  inv02 U4788 ( .Y(n7833), .A(n7495) );
  nor02 U4789 ( .Y(n7496), .A0(n7947), .A1(n7698) );
  nor02 U4790 ( .Y(n7497), .A0(n7949), .A1(n7701) );
  inv01 U4791 ( .Y(n7498), .A(n4385) );
  nor02 U4792 ( .Y(n7495), .A0(n7498), .A1(n7499) );
  nor02 U4793 ( .Y(n7500), .A0(n7496), .A1(n7497) );
  inv01 U4794 ( .Y(n7499), .A(n7500) );
  inv02 U4795 ( .Y(n7947), .A(fract_28_i[19]) );
  buf04 U4796 ( .Y(n7698), .A(n7876) );
  nor02 U4797 ( .Y(n7502), .A0(n7873), .A1(n7703) );
  nor02 U4798 ( .Y(n7503), .A0(n7875), .A1(n7702) );
  inv01 U4799 ( .Y(n7504), .A(n4365) );
  nor02 U4800 ( .Y(n7501), .A0(n7504), .A1(n7505) );
  nor02 U4801 ( .Y(n7506), .A0(n7502), .A1(n7503) );
  inv01 U4802 ( .Y(n7505), .A(n7506) );
  nor02 U4803 ( .Y(n7508), .A0(n7932), .A1(n7699) );
  nor02 U4804 ( .Y(n7509), .A0(n7604), .A1(n7701) );
  inv01 U4805 ( .Y(n7510), .A(n4396) );
  nor02 U4806 ( .Y(n7507), .A0(n7510), .A1(n7511) );
  nor02 U4807 ( .Y(n7512), .A0(n7508), .A1(n7509) );
  inv02 U4808 ( .Y(n7511), .A(n7512) );
  inv02 U4809 ( .Y(n7873), .A(fract_28_i[9]) );
  inv02 U4810 ( .Y(n7834), .A(n7513) );
  nor02 U4811 ( .Y(n7514), .A0(n7606), .A1(n7698) );
  nor02 U4812 ( .Y(n7515), .A0(n7974), .A1(n7701) );
  inv01 U4813 ( .Y(n7516), .A(n4412) );
  nor02 U4814 ( .Y(n7513), .A0(n7516), .A1(n7517) );
  nor02 U4815 ( .Y(n7518), .A0(n7514), .A1(n7515) );
  inv01 U4816 ( .Y(n7517), .A(n7518) );
  inv02 U4817 ( .Y(n7606), .A(n7605) );
  inv02 U4818 ( .Y(n7935), .A(n7519) );
  nor02 U4819 ( .Y(n7520), .A0(n7875), .A1(n7703) );
  nor02 U4820 ( .Y(n7521), .A0(n7956), .A1(n7702) );
  inv01 U4821 ( .Y(n7522), .A(n4420) );
  nor02 U4822 ( .Y(n7519), .A0(n7522), .A1(n7523) );
  nor02 U4823 ( .Y(n7524), .A0(n7520), .A1(n7521) );
  inv01 U4824 ( .Y(n7523), .A(n7524) );
  inv02 U4825 ( .Y(n7840), .A(n7525) );
  nor02 U4826 ( .Y(n7526), .A0(n7949), .A1(n7698) );
  nor02 U4827 ( .Y(n7527), .A0(n7961), .A1(n7701) );
  inv01 U4828 ( .Y(n7528), .A(n7994) );
  nor02 U4829 ( .Y(n7525), .A0(n7528), .A1(n7529) );
  nor02 U4830 ( .Y(n7530), .A0(n7526), .A1(n7527) );
  inv01 U4831 ( .Y(n7529), .A(n7530) );
  inv02 U4832 ( .Y(n8044), .A(n7531) );
  inv01 U4833 ( .Y(n7532), .A(n8107) );
  inv01 U4834 ( .Y(n7533), .A(n8047) );
  inv01 U4835 ( .Y(n7534), .A(n8048) );
  nand02 U4836 ( .Y(n7531), .A0(n7534), .A1(n7535) );
  nand02 U4837 ( .Y(n7536), .A0(n7532), .A1(n7533) );
  inv01 U4838 ( .Y(n7535), .A(n7536) );
  inv02 U4839 ( .Y(n8017), .A(n8022) );
  inv02 U4840 ( .Y(n8072), .A(n7537) );
  nand02 U4841 ( .Y(n7537), .A0(n7429), .A1(n7538) );
  nand02 U4842 ( .Y(n7539), .A0(n6660), .A1(n7932) );
  inv01 U4843 ( .Y(n7538), .A(n7539) );
  buf02 U4844 ( .Y(n7540), .A(n7943) );
  inv02 U4845 ( .Y(n7943), .A(fract_28_i[20]) );
  or02 U4846 ( .Y(n7541), .A0(fract_28_i[27]), .A1(n4489) );
  inv02 U4847 ( .Y(n7542), .A(n7541) );
  buf02 U4848 ( .Y(n7543), .A(n8035) );
  buf02 U4849 ( .Y(n7544), .A(n8035) );
  inv02 U4850 ( .Y(n7787), .A(n7545) );
  inv01 U4851 ( .Y(n7546), .A(rmode_i[1]) );
  nor02 U4852 ( .Y(n7547), .A0(n4251), .A1(n7546) );
  nor02 U4853 ( .Y(n7548), .A0(rmode_i[1]), .A1(n7809) );
  nor02 U4854 ( .Y(n7545), .A0(n7547), .A1(n7548) );
  or02 U4855 ( .Y(n7549), .A0(fract_28_i[27]), .A1(n4257) );
  inv02 U4856 ( .Y(n7550), .A(n7549) );
  nor02 U4857 ( .Y(n7552), .A0(n7880), .A1(n7703) );
  nor02 U4858 ( .Y(n7553), .A0(n7879), .A1(n7702) );
  inv01 U4859 ( .Y(n7554), .A(n4259) );
  nor02 U4860 ( .Y(n7551), .A0(n7554), .A1(n7555) );
  nor02 U4861 ( .Y(n7556), .A0(n7552), .A1(n7553) );
  inv02 U4862 ( .Y(n7555), .A(n7556) );
  inv02 U4863 ( .Y(n7852), .A(n7557) );
  nor02 U4864 ( .Y(n7558), .A0(n7902), .A1(n7699) );
  nor02 U4865 ( .Y(n7559), .A0(n7701), .A1(n7911) );
  inv01 U4866 ( .Y(n7560), .A(n8000) );
  nor02 U4867 ( .Y(n7557), .A0(n7560), .A1(n7561) );
  nor02 U4868 ( .Y(n7562), .A0(n7558), .A1(n7559) );
  inv01 U4869 ( .Y(n7561), .A(n7562) );
  nor02 U4870 ( .Y(n7564), .A0(n7889), .A1(n7703) );
  nor02 U4871 ( .Y(n7565), .A0(n7880), .A1(n7702) );
  inv01 U4872 ( .Y(n7566), .A(n4253) );
  nor02 U4873 ( .Y(n7563), .A0(n7566), .A1(n7567) );
  nor02 U4874 ( .Y(n7568), .A0(n7564), .A1(n7565) );
  inv02 U4875 ( .Y(n7567), .A(n7568) );
  inv02 U4876 ( .Y(n7911), .A(fract_28_i[24]) );
  inv02 U4877 ( .Y(n7902), .A(fract_28_i[25]) );
  ao22 U4878 ( .Y(n7569), .A0(n2768_27_), .A1(n7788), .B0(s_fracto28_1[27]), 
        .B1(n7787) );
  inv02 U4879 ( .Y(n7570), .A(n7569) );
  nor02 U4880 ( .Y(n7572), .A0(n7879), .A1(n7703) );
  nor02 U4881 ( .Y(n7573), .A0(n7882), .A1(n7702) );
  inv01 U4882 ( .Y(n7574), .A(n4285) );
  nor02 U4883 ( .Y(n7571), .A0(n7574), .A1(n7575) );
  nor02 U4884 ( .Y(n7576), .A0(n7572), .A1(n7573) );
  inv02 U4885 ( .Y(n7575), .A(n7576) );
  inv02 U4886 ( .Y(n7882), .A(fract_28_i[6]) );
  or02 U4887 ( .Y(n7577), .A0(n7844), .A1(s_shr1_2_) );
  inv02 U4888 ( .Y(n7578), .A(n7577) );
  nor02 U4889 ( .Y(n7580), .A0(n7922), .A1(n7700) );
  nor02 U4890 ( .Y(n7581), .A0(n7932), .A1(n7701) );
  inv01 U4891 ( .Y(n7582), .A(n8013) );
  nor02 U4892 ( .Y(n7579), .A0(n7582), .A1(n7583) );
  nor02 U4893 ( .Y(n7584), .A0(n7580), .A1(n7581) );
  inv02 U4894 ( .Y(n7583), .A(n7584) );
  inv02 U4895 ( .Y(n7932), .A(fract_28_i[22]) );
  or02 U4896 ( .Y(n7585), .A0(n7866), .A1(s_shl1_2_) );
  inv02 U4897 ( .Y(n7586), .A(n7585) );
  nor02 U4898 ( .Y(n7588), .A0(n7700), .A1(n7911) );
  nor02 U4899 ( .Y(n7589), .A0(n7922), .A1(n7701) );
  inv01 U4900 ( .Y(n7590), .A(n4464) );
  nor02 U4901 ( .Y(n7587), .A0(n7590), .A1(n7591) );
  nor02 U4902 ( .Y(n7592), .A0(n7588), .A1(n7589) );
  inv02 U4903 ( .Y(n7591), .A(n7592) );
  inv02 U4904 ( .Y(n7922), .A(fract_28_i[23]) );
  and02 U4905 ( .Y(n7594), .A0(s_shr1_2_), .A1(n7844) );
  and02 U4906 ( .Y(n7593), .A0(s_shr1_2_), .A1(n7844) );
  inv02 U4907 ( .Y(n7844), .A(s_shr1_3_) );
  and02 U4908 ( .Y(n7596), .A0(s_shl1_2_), .A1(n7866) );
  and02 U4909 ( .Y(n7595), .A0(s_shl1_2_), .A1(n7866) );
  inv02 U4910 ( .Y(n7866), .A(s_shl1_3_) );
  inv02 U4911 ( .Y(n7861), .A(n7597) );
  nor02 U4912 ( .Y(n7598), .A0(n7804), .A1(n7702) );
  nor02 U4913 ( .Y(n7599), .A0(n7986), .A1(n7987) );
  nor02 U4914 ( .Y(n7597), .A0(n7598), .A1(n7599) );
  inv02 U4915 ( .Y(n7986), .A(fract_28_i[1]) );
  inv01 U4916 ( .Y(n7600), .A(n7851) );
  inv01 U4917 ( .Y(n7601), .A(n7600) );
  inv01 U4918 ( .Y(n7603), .A(n7600) );
  inv01 U4919 ( .Y(n7602), .A(n7600) );
  buf02 U4920 ( .Y(n7604), .A(n7941) );
  buf02 U4921 ( .Y(n7605), .A(fract_28_i[15]) );
  inv01 U4922 ( .Y(n7607), .A(fract_28_i[17]) );
  inv02 U4923 ( .Y(n7941), .A(fract_28_i[21]) );
  inv02 U4924 ( .Y(n7961), .A(fract_28_i[17]) );
  inv02 U4925 ( .Y(n7848), .A(n7608) );
  nor02 U4926 ( .Y(n7609), .A0(n7986), .A1(n7703) );
  nor02 U4927 ( .Y(n7610), .A0(n7955), .A1(n7702) );
  inv01 U4928 ( .Y(n7611), .A(n4263) );
  nor02 U4929 ( .Y(n7608), .A0(n7611), .A1(n7612) );
  nor02 U4930 ( .Y(n7613), .A0(n7609), .A1(n7610) );
  inv01 U4931 ( .Y(n7612), .A(n7613) );
  nand02 U4932 ( .Y(n7614), .A0(n7648), .A1(n7640) );
  nor02 U4933 ( .Y(n7617), .A0(n7704), .A1(n7699) );
  nor02 U4934 ( .Y(n7618), .A0(n7900), .A1(n7701) );
  inv01 U4935 ( .Y(n7619), .A(n4271) );
  nor02 U4936 ( .Y(n7616), .A0(n7619), .A1(n7620) );
  nor02 U4937 ( .Y(n7621), .A0(n7617), .A1(n7618) );
  inv01 U4938 ( .Y(n7620), .A(n7621) );
  nand02 U4939 ( .Y(n7622), .A0(n7626), .A1(n7649) );
  buf02 U4940 ( .Y(n7624), .A(n7845) );
  buf02 U4941 ( .Y(n7626), .A(n7845) );
  buf02 U4942 ( .Y(n7625), .A(n7845) );
  inv02 U4943 ( .Y(n7854), .A(n7627) );
  nor02 U4944 ( .Y(n7628), .A0(n7955), .A1(n7987) );
  nor02 U4945 ( .Y(n7629), .A0(n7986), .A1(n7702) );
  nor02 U4946 ( .Y(n7630), .A0(n7804), .A1(n7703) );
  nor02 U4947 ( .Y(n7627), .A0(n7630), .A1(n7631) );
  nor02 U4948 ( .Y(n7632), .A0(n7628), .A1(n7629) );
  inv01 U4949 ( .Y(n7631), .A(n7632) );
  inv02 U4950 ( .Y(n7819), .A(n7633) );
  nor02 U4951 ( .Y(n7634), .A0(n7704), .A1(n7701) );
  nor02 U4952 ( .Y(n7635), .A0(n7902), .A1(n7988) );
  nor02 U4953 ( .Y(n7636), .A0(n7881), .A1(n7900) );
  nor02 U4954 ( .Y(n7633), .A0(n7636), .A1(n7637) );
  nor02 U4955 ( .Y(n7638), .A0(n7634), .A1(n7635) );
  inv01 U4956 ( .Y(n7637), .A(n7638) );
  inv02 U4957 ( .Y(n7804), .A(fract_28_i[0]) );
  inv02 U4958 ( .Y(n7987), .A(n7695) );
  inv02 U4959 ( .Y(n7988), .A(n7690) );
  buf02 U4960 ( .Y(n7639), .A(n7921) );
  buf02 U4961 ( .Y(n7640), .A(n7921) );
  ao21 U4962 ( .Y(n7641), .A0(n7789), .A1(n7790), .B0(n7791) );
  inv01 U4963 ( .Y(n7642), .A(n7641) );
  inv02 U4964 ( .Y(n7643), .A(n7641) );
  ao21 U4965 ( .Y(n7644), .A0(n7710), .A1(n7711), .B0(n7712) );
  inv02 U4966 ( .Y(n7645), .A(n7644) );
  inv02 U4967 ( .Y(n7646), .A(n7891) );
  inv02 U4968 ( .Y(n7647), .A(n7646) );
  inv02 U4969 ( .Y(n7648), .A(n7646) );
  buf04 U4970 ( .Y(n7649), .A(n7964) );
  buf04 U4971 ( .Y(n7650), .A(n7733) );
  inv04 U4972 ( .Y(n7704), .A(fract_28_i[27]) );
  inv04 U4973 ( .Y(n7706), .A(n7705) );
  inv02 U4974 ( .Y(n7652), .A(n7939) );
  inv02 U4975 ( .Y(n7653), .A(n7652) );
  inv02 U4976 ( .Y(n7655), .A(n7652) );
  inv02 U4977 ( .Y(n7654), .A(n7652) );
  inv02 U4978 ( .Y(n7656), .A(n7820) );
  inv02 U4979 ( .Y(n7657), .A(n7656) );
  inv02 U4980 ( .Y(n7660), .A(n7656) );
  inv02 U4981 ( .Y(n7658), .A(n7656) );
  inv01 U4982 ( .Y(n7659), .A(n7656) );
  inv01 U4983 ( .Y(n7662), .A(n7792) );
  inv01 U4984 ( .Y(n7663), .A(n7413) );
  inv01 U4985 ( .Y(n7664), .A(n7427) );
  nand02 U4986 ( .Y(n7661), .A0(n7664), .A1(n7665) );
  nand02 U4987 ( .Y(n7666), .A0(n7662), .A1(n7663) );
  inv01 U4988 ( .Y(n7665), .A(n7666) );
  buf02 U4989 ( .Y(n7671), .A(n7824) );
  buf02 U4990 ( .Y(n7673), .A(n7824) );
  buf02 U4991 ( .Y(n7672), .A(n7824) );
  buf08 U4992 ( .Y(n7675), .A(n7817) );
  buf08 U4993 ( .Y(n7677), .A(n7822) );
  buf16 U4994 ( .Y(n7678), .A(n7841) );
  inv08 U4995 ( .Y(n7679), .A(n7881) );
  inv04 U4996 ( .Y(n7881), .A(n7421) );
  buf08 U4997 ( .Y(n7680), .A(n7714) );
  nand02 U4998 ( .Y(n7681), .A0(n7643), .A1(n7682) );
  nand02 U4999 ( .Y(n7683), .A0(n7570), .A1(n7788) );
  inv01 U5000 ( .Y(n7682), .A(n7683) );
  buf08 U5001 ( .Y(n7684), .A(n7717) );
  nand02 U5002 ( .Y(n7685), .A0(n7643), .A1(n7686) );
  nand02 U5003 ( .Y(n7687), .A0(n7752), .A1(n7788) );
  inv01 U5004 ( .Y(n7686), .A(n7687) );
  inv02 U5005 ( .Y(n7788), .A(n7787) );
  inv02 U5006 ( .Y(n7752), .A(n7570) );
  inv02 U5007 ( .Y(n7688), .A(n7878) );
  inv04 U5008 ( .Y(n7689), .A(n7688) );
  inv04 U5009 ( .Y(n7690), .A(n7688) );
  inv02 U5010 ( .Y(n7691), .A(n7904) );
  inv02 U5011 ( .Y(n7692), .A(n7691) );
  inv04 U5012 ( .Y(n7694), .A(n7691) );
  buf12 U5013 ( .Y(n7695), .A(n7905) );
  nand02 U5014 ( .Y(n7696), .A0(s_shr1_1_), .A1(s_shr1_0_) );
  nand02 U5015 ( .Y(n7697), .A0(s_shr1_1_), .A1(s_shr1_0_) );
  buf16 U5016 ( .Y(n7701), .A(n7874) );
  buf16 U5017 ( .Y(n7702), .A(n7901) );
  buf16 U5018 ( .Y(n7703), .A(n7903) );
  nor02 U5019 ( .Y(n7790), .A0(n7708), .A1(n4489) );
  and02 U5020 ( .Y(s_shl11786_5_), .A0(n____return1927_5_), .A1(n7645) );
  inv01 U5021 ( .Y(n8031), .A(n4712) );
  inv01 U5022 ( .Y(n8042), .A(n4712) );
  nand03 U5023 ( .Y(n8054), .A0(n8056), .A1(n8057), .A2(n8055) );
  inv01 U5024 ( .Y(n8057), .A(n8061) );
  inv01 U5025 ( .Y(n8056), .A(n8065) );
  nor02 U5026 ( .Y(n8055), .A0(n4620), .A1(n8067) );
  nor02 U5027 ( .Y(n8070), .A0(n8075), .A1(n4610) );
  inv01 U5028 ( .Y(n8069), .A(n8078) );
  inv01 U5029 ( .Y(n8084), .A(n8085) );
  nor02 U5030 ( .Y(n8085), .A0(n8064), .A1(n8066) );
  inv01 U5031 ( .Y(n8087), .A(n4610) );
  nor02 U5032 ( .Y(n8086), .A0(n8077), .A1(n8079) );
  nand02 U5033 ( .Y(n8091), .A0(n8092), .A1(n8093) );
  nor02 U5034 ( .Y(n8093), .A0(n8060), .A1(n8058) );
  nor02 U5035 ( .Y(n8092), .A0(n4620), .A1(n8067) );
  inv01 U5036 ( .Y(n8096), .A(n8076) );
  inv01 U5037 ( .Y(n8094), .A(n8059) );
  nor02 U5038 ( .Y(n8101), .A0(n8062), .A1(n8058) );
  nor02 U5039 ( .Y(n8100), .A0(n8063), .A1(n8061) );
  nor02 U5040 ( .Y(n8099), .A0(n4620), .A1(n8067) );
  inv01 U5041 ( .Y(n8097), .A(n4570) );
  ao22 U5042 ( .Y(s_shl11786_4_), .A0(n7706), .A1(n7707), .B0(
        n____return1927_4_), .B1(n7645) );
  ao22 U5043 ( .Y(s_shl11786_3_), .A0(n7706), .A1(n7542), .B0(
        n____return1927_3_), .B1(n7645) );
  ao22 U5044 ( .Y(s_shl11786_2_), .A0(n7706), .A1(n7708), .B0(
        n____return1927_2_), .B1(n7645) );
  ao22 U5045 ( .Y(s_shl11786_1_), .A0(n7706), .A1(n7550), .B0(
        n____return1927_1_), .B1(n7645) );
  ao22 U5046 ( .Y(s_shl11786_0_), .A0(n____return1927_0_), .A1(n7645), .B0(
        n7709), .B1(n7706) );
  ao221 U5047 ( .Y(s_output_o[9]), .A0(n7713), .A1(n____return2766_13_), .B0(
        n7680), .B1(s_fracto28_1[13]), .C0(n7715) );
  ao22 U5048 ( .Y(n7715), .A0(n____return2766_12_), .A1(n7716), .B0(
        s_fracto28_1[12]), .B1(n7684) );
  ao221 U5049 ( .Y(s_output_o[8]), .A0(n____return2766_12_), .A1(n7713), .B0(
        s_fracto28_1[12]), .B1(n7680), .C0(n7718) );
  ao22 U5050 ( .Y(n7718), .A0(n____return2766_11_), .A1(n7716), .B0(
        s_fracto28_1[11]), .B1(n7684) );
  ao221 U5051 ( .Y(s_output_o[7]), .A0(n7713), .A1(n____return2766_11_), .B0(
        n7680), .B1(s_fracto28_1[11]), .C0(n7719) );
  ao22 U5052 ( .Y(n7719), .A0(n____return2766_10_), .A1(n7716), .B0(
        s_fracto28_1[10]), .B1(n7684) );
  ao221 U5053 ( .Y(s_output_o[6]), .A0(n7713), .A1(n____return2766_10_), .B0(
        n7680), .B1(s_fracto28_1[10]), .C0(n7720) );
  ao22 U5054 ( .Y(n7720), .A0(n____return2766_9_), .A1(n7716), .B0(
        s_fracto28_1[9]), .B1(n7684) );
  ao221 U5055 ( .Y(s_output_o[5]), .A0(n7713), .A1(n____return2766_9_), .B0(
        n7680), .B1(s_fracto28_1[9]), .C0(n7721) );
  ao22 U5056 ( .Y(n7721), .A0(n____return2766_8_), .A1(n7716), .B0(
        s_fracto28_1[8]), .B1(n7684) );
  ao221 U5057 ( .Y(s_output_o[4]), .A0(n7713), .A1(n____return2766_8_), .B0(
        n7680), .B1(s_fracto28_1[8]), .C0(n7722) );
  ao22 U5058 ( .Y(n7722), .A0(n____return2766_7_), .A1(n7716), .B0(
        s_fracto28_1[7]), .B1(n7684) );
  ao221 U5059 ( .Y(s_output_o[3]), .A0(n7713), .A1(n____return2766_7_), .B0(
        n7680), .B1(s_fracto28_1[7]), .C0(n7723) );
  ao22 U5060 ( .Y(n7723), .A0(n____return2766_6_), .A1(n7716), .B0(
        s_fracto28_1[6]), .B1(n7684) );
  nor02 U5061 ( .Y(n7727), .A0(n7725), .A1(n7726) );
  and03 U5062 ( .Y(n7726), .A0(n7427), .A1(n4708), .A2(n7730) );
  inv01 U5063 ( .Y(n7732), .A(n____return2864_7_) );
  ao221 U5064 ( .Y(s_output_o[2]), .A0(n7713), .A1(n____return2766_6_), .B0(
        n7680), .B1(s_fracto28_1[6]), .C0(n7737) );
  ao22 U5065 ( .Y(n7737), .A0(n____return2766_5_), .A1(n7716), .B0(
        s_fracto28_1[5]), .B1(n7684) );
  inv01 U5066 ( .Y(n7738), .A(n____return2864_6_) );
  inv01 U5067 ( .Y(n7746), .A(n____return2864_2_) );
  inv01 U5068 ( .Y(n7748), .A(n____return2864_1_) );
  nand02 U5069 ( .Y(n7735), .A0(n7643), .A1(n7570) );
  nand02 U5070 ( .Y(n7733), .A0(n7643), .A1(n7752) );
  nand03 U5071 ( .Y(s_output_o[22]), .A0(n7725), .A1(n7753), .A2(n7754) );
  nand02 U5072 ( .Y(n7753), .A0(s_fracto28_1[26]), .A1(n7680) );
  nand04 U5073 ( .Y(n7757), .A0(n4524), .A1(n7758), .A2(n7759), .A3(n7760) );
  nand04 U5074 ( .Y(n7756), .A0(n7761), .A1(n7762), .A2(n7763), .A3(n7764) );
  ao21 U5075 ( .Y(n7755), .A0(n7413), .A1(n4651), .B0(n4708) );
  nand04 U5076 ( .Y(n7729), .A0(n7765), .A1(n7766), .A2(n7767), .A3(n7768) );
  or03 U5077 ( .Y(n7769), .A0(opb_i[9]), .A1(opb_i[8]), .A2(opb_i[7]) );
  or03 U5078 ( .Y(n7770), .A0(opb_i[3]), .A1(opb_i[21]), .A2(opb_i[22]) );
  or03 U5079 ( .Y(n7771), .A0(opb_i[14]), .A1(opb_i[15]), .A2(opb_i[17]) );
  or02 U5080 ( .Y(n7772), .A0(opb_i[13]), .A1(opb_i[12]) );
  ao221 U5081 ( .Y(s_output_o[21]), .A0(n7713), .A1(n____return2766_25_), .B0(
        n7680), .B1(s_fracto28_1[25]), .C0(n7773) );
  ao22 U5082 ( .Y(n7773), .A0(n____return2766_24_), .A1(n7716), .B0(
        s_fracto28_1[24]), .B1(n7684) );
  ao221 U5083 ( .Y(s_output_o[20]), .A0(n7713), .A1(n____return2766_24_), .B0(
        n7680), .B1(s_fracto28_1[24]), .C0(n7774) );
  ao22 U5084 ( .Y(n7774), .A0(n____return2766_23_), .A1(n7716), .B0(
        s_fracto28_1[23]), .B1(n7684) );
  ao221 U5085 ( .Y(s_output_o[1]), .A0(n7713), .A1(n____return2766_5_), .B0(
        n7680), .B1(s_fracto28_1[5]), .C0(n7775) );
  ao22 U5086 ( .Y(n7775), .A0(n____return2766_4_), .A1(n7716), .B0(
        s_fracto28_1[4]), .B1(n7684) );
  ao221 U5087 ( .Y(s_output_o[19]), .A0(n7713), .A1(n____return2766_23_), .B0(
        n7680), .B1(s_fracto28_1[23]), .C0(n7776) );
  ao22 U5088 ( .Y(n7776), .A0(n____return2766_22_), .A1(n7716), .B0(
        s_fracto28_1[22]), .B1(n7684) );
  ao221 U5089 ( .Y(s_output_o[18]), .A0(n7713), .A1(n____return2766_22_), .B0(
        n7680), .B1(s_fracto28_1[22]), .C0(n7777) );
  ao22 U5090 ( .Y(n7777), .A0(n____return2766_21_), .A1(n7716), .B0(
        s_fracto28_1[21]), .B1(n7684) );
  ao221 U5091 ( .Y(s_output_o[17]), .A0(n7713), .A1(n____return2766_21_), .B0(
        n7680), .B1(s_fracto28_1[21]), .C0(n7778) );
  ao22 U5092 ( .Y(n7778), .A0(n____return2766_20_), .A1(n7716), .B0(
        s_fracto28_1[20]), .B1(n7684) );
  ao221 U5093 ( .Y(s_output_o[16]), .A0(n7713), .A1(n____return2766_20_), .B0(
        n7680), .B1(s_fracto28_1[20]), .C0(n7779) );
  ao22 U5094 ( .Y(n7779), .A0(n____return2766_19_), .A1(n7716), .B0(
        s_fracto28_1[19]), .B1(n7684) );
  ao221 U5095 ( .Y(s_output_o[15]), .A0(n7713), .A1(n____return2766_19_), .B0(
        n7680), .B1(s_fracto28_1[19]), .C0(n7780) );
  ao22 U5096 ( .Y(n7780), .A0(n____return2766_18_), .A1(n7716), .B0(
        s_fracto28_1[18]), .B1(n7684) );
  ao221 U5097 ( .Y(s_output_o[14]), .A0(n7713), .A1(n____return2766_18_), .B0(
        n7680), .B1(s_fracto28_1[18]), .C0(n7781) );
  ao22 U5098 ( .Y(n7781), .A0(n____return2766_17_), .A1(n7716), .B0(
        s_fracto28_1[17]), .B1(n7684) );
  ao221 U5099 ( .Y(s_output_o[13]), .A0(n7713), .A1(n____return2766_17_), .B0(
        n7680), .B1(s_fracto28_1[17]), .C0(n7782) );
  ao22 U5100 ( .Y(n7782), .A0(n____return2766_16_), .A1(n7716), .B0(
        s_fracto28_1[16]), .B1(n7684) );
  ao221 U5101 ( .Y(s_output_o[12]), .A0(n7713), .A1(n____return2766_16_), .B0(
        n7680), .B1(s_fracto28_1[16]), .C0(n7783) );
  ao22 U5102 ( .Y(n7783), .A0(n____return2766_15_), .A1(n7716), .B0(
        s_fracto28_1[15]), .B1(n7684) );
  ao221 U5103 ( .Y(s_output_o[11]), .A0(n7713), .A1(n____return2766_15_), .B0(
        n7680), .B1(s_fracto28_1[15]), .C0(n7784) );
  ao22 U5104 ( .Y(n7784), .A0(n____return2766_14_), .A1(n7716), .B0(
        s_fracto28_1[14]), .B1(n7684) );
  ao221 U5105 ( .Y(s_output_o[10]), .A0(n7713), .A1(n____return2766_14_), .B0(
        n7680), .B1(s_fracto28_1[14]), .C0(n7785) );
  ao22 U5106 ( .Y(n7785), .A0(n____return2766_13_), .A1(n7716), .B0(
        s_fracto28_1[13]), .B1(n7684) );
  ao221 U5107 ( .Y(s_output_o[0]), .A0(n7713), .A1(n____return2766_4_), .B0(
        n7680), .B1(s_fracto28_1[4]), .C0(n7786) );
  ao22 U5108 ( .Y(n7786), .A0(n____return2766_3_), .A1(n7716), .B0(
        s_fracto28_1[3]), .B1(n7684) );
  and03 U5109 ( .Y(n7717), .A0(n7570), .A1(n7787), .A2(n7642) );
  and03 U5110 ( .Y(n7714), .A0(n7787), .A1(n7752), .A2(n7642) );
  inv01 U5111 ( .Y(n7791), .A(n7736) );
  inv01 U5112 ( .Y(n7792), .A(n7802) );
  inv01 U5113 ( .Y(n7742), .A(n____return2864_4_) );
  inv01 U5114 ( .Y(n7744), .A(n____return2864_3_) );
  inv01 U5115 ( .Y(n7740), .A(n____return2864_5_) );
  nand02 U5116 ( .Y(n7803), .A0(n____return2864_7_), .A1(n____return2864_6_)
         );
  inv01 U5117 ( .Y(n7750), .A(n____return2864_0_) );
  nor02 U5118 ( .Y(n7801), .A0(n7804), .A1(n7805) );
  and02 U5119 ( .Y(n7807), .A0(n7752), .A1(s_fracto28_1[3]) );
  and02 U5120 ( .Y(n7808), .A0(n7752), .A1(n____return2766_3_) );
  inv01 U5121 ( .Y(n7810), .A(n7812) );
  nor02 U5122 ( .Y(n7813), .A0(s_fracto28_1[3]), .A1(n7812) );
  ao21 U5123 ( .Y(n7812), .A0(fract_28_i[0]), .A1(fract_28_i[27]), .B0(n7814)
         );
  or02 U5124 ( .Y(n7814), .A0(s_fracto28_1[0]), .A1(s_fracto28_1[1]) );
  inv01 U5125 ( .Y(n7811), .A(s_fracto28_1[2]) );
  nand02 U5126 ( .Y(s_fracto28_12090_9_), .A0(n7815), .A1(n7816) );
  nand02 U5127 ( .Y(s_fracto28_12090_8_), .A0(n7828), .A1(n7829) );
  nand03 U5128 ( .Y(s_fracto28_12090_7_), .A0(n7836), .A1(n7837), .A2(n7838)
         );
  nand04 U5129 ( .Y(s_fracto28_12090_6_), .A0(n4574), .A1(n4584), .A2(n4624), 
        .A3(n4659) );
  nand03 U5130 ( .Y(s_fracto28_12090_4_), .A0(n4497), .A1(n7863), .A2(n7864)
         );
  and02 U5131 ( .Y(n7850), .A0(n7594), .A1(n7626) );
  nand02 U5132 ( .Y(s_fracto28_12090_3_), .A0(n7869), .A1(n7870) );
  nand02 U5133 ( .Y(s_fracto28_12090_2_), .A0(n7883), .A1(n7884) );
  ao221 U5134 ( .Y(s_fracto28_12090_27_), .A0(n7890), .A1(n7647), .B0(n7892), 
        .B1(n7674), .C0(n7894) );
  inv01 U5135 ( .Y(n7894), .A(n7895) );
  nand02 U5136 ( .Y(s_fracto28_12090_26_), .A0(n7906), .A1(n7907) );
  nand02 U5137 ( .Y(s_fracto28_12090_25_), .A0(n7914), .A1(n7915) );
  nand02 U5138 ( .Y(s_fracto28_12090_24_), .A0(n7925), .A1(n7926) );
  nand03 U5139 ( .Y(s_fracto28_12090_23_), .A0(n4494), .A1(n7936), .A2(n7937)
         );
  nand04 U5140 ( .Y(s_fracto28_12090_22_), .A0(n4568), .A1(n4607), .A2(n4616), 
        .A3(n7942) );
  nand04 U5141 ( .Y(s_fracto28_12090_21_), .A0(n4576), .A1(n7945), .A2(n4618), 
        .A3(n7946) );
  and02 U5142 ( .Y(n7940), .A0(n7648), .A1(n7596) );
  nand03 U5143 ( .Y(s_fracto28_12090_20_), .A0(n4485), .A1(n4864), .A2(n7948)
         );
  nand02 U5144 ( .Y(s_fracto28_12090_1_), .A0(n7951), .A1(n7952) );
  nand02 U5145 ( .Y(s_fracto28_12090_19_), .A0(n7959), .A1(n7960) );
  nand02 U5146 ( .Y(s_fracto28_12090_18_), .A0(n7965), .A1(n7966) );
  nand02 U5147 ( .Y(s_fracto28_12090_17_), .A0(n7969), .A1(n7970) );
  nand02 U5148 ( .Y(s_fracto28_12090_16_), .A0(n7972), .A1(n7973) );
  nor02 U5149 ( .Y(n7891), .A0(n7976), .A1(n4608) );
  inv01 U5150 ( .Y(n7976), .A(s_shl1_4_) );
  nand03 U5151 ( .Y(s_fracto28_12090_15_), .A0(n4511), .A1(n4885), .A2(n7979)
         );
  mux21 U5152 ( .Y(n7981), .A0(n7963), .A1(n7297), .S0(s_shr1_2_) );
  nand04 U5153 ( .Y(s_fracto28_12090_14_), .A0(n7982), .A1(n4592), .A2(n4612), 
        .A3(n4647) );
  and02 U5154 ( .Y(n7896), .A0(n7657), .A1(n7586) );
  and03 U5155 ( .Y(n7893), .A0(s_shl1_2_), .A1(s_shl1_3_), .A2(n7658) );
  nand03 U5156 ( .Y(s_fracto28_12090_12_), .A0(n4487), .A1(n7989), .A2(n7990)
         );
  mux21 U5157 ( .Y(n7991), .A0(n7930), .A1(n7431), .S0(s_shl1_2_) );
  and02 U5158 ( .Y(n7847), .A0(n7660), .A1(n7919) );
  nand02 U5159 ( .Y(s_fracto28_12090_11_), .A0(n7992), .A1(n7993) );
  inv01 U5160 ( .Y(n7890), .A(n7996) );
  nand02 U5161 ( .Y(s_fracto28_12090_10_), .A0(n7997), .A1(n7998) );
  and02 U5162 ( .Y(n7817), .A0(n7655), .A1(n7649) );
  and02 U5163 ( .Y(n7919), .A0(s_shl1_2_), .A1(n7866) );
  nor02 U5164 ( .Y(n7904), .A0(n8002), .A1(n8003) );
  nand02 U5165 ( .Y(n7903), .A0(s_shl1_1_), .A1(n8003) );
  inv01 U5166 ( .Y(n8003), .A(s_shl1_0_) );
  nand02 U5167 ( .Y(n7901), .A0(s_shl1_0_), .A1(n8002) );
  inv01 U5168 ( .Y(n8002), .A(s_shl1_1_) );
  nand02 U5169 ( .Y(s_fracto28_12090_0_), .A0(n8004), .A1(n8005) );
  nor02 U5170 ( .Y(n7905), .A0(s_shl1_1_), .A1(s_shl1_0_) );
  and02 U5171 ( .Y(n7841), .A0(n7659), .A1(n7639) );
  nor02 U5172 ( .Y(n7921), .A0(s_shl1_3_), .A1(s_shl1_2_) );
  nor02 U5173 ( .Y(n7820), .A0(n4608), .A1(s_shl1_4_) );
  nand04 U5174 ( .Y(n7977), .A0(n7689), .A1(n7310), .A2(n8114), .A3(n8009) );
  inv01 U5175 ( .Y(n8009), .A(s_shr1_5_) );
  and02 U5176 ( .Y(n7822), .A0(n7867), .A1(n7653) );
  and02 U5177 ( .Y(n7826), .A0(n7578), .A1(n7655) );
  and03 U5178 ( .Y(n7824), .A0(s_shr1_2_), .A1(n7654), .A2(s_shr1_3_) );
  nor02 U5179 ( .Y(n7939), .A0(n8011), .A1(s_shr1_4_) );
  and02 U5180 ( .Y(n7867), .A0(s_shr1_2_), .A1(n7844) );
  nand02 U5181 ( .Y(n7876), .A0(s_shr1_1_), .A1(s_shr1_0_) );
  nand02 U5182 ( .Y(n7874), .A0(s_shr1_1_), .A1(n7805) );
  and02 U5183 ( .Y(n7845), .A0(s_shr1_4_), .A1(n8007) );
  inv01 U5184 ( .Y(n8007), .A(n8011) );
  ao21 U5185 ( .Y(n8011), .A0(n7690), .A1(n7311), .B0(s_shr1_5_) );
  nor02 U5186 ( .Y(n8008), .A0(n8014), .A1(s_shr1_4_) );
  inv01 U5187 ( .Y(n8014), .A(n7649) );
  nor02 U5188 ( .Y(n7964), .A0(s_shr1_3_), .A1(s_shr1_2_) );
  nor02 U5189 ( .Y(n7878), .A0(s_shr1_1_), .A1(s_shr1_0_) );
  inv01 U5190 ( .Y(s_expo9_2[7]), .A(n7734) );
  inv01 U5191 ( .Y(s_expo9_2[6]), .A(n7739) );
  inv01 U5192 ( .Y(s_expo9_2[3]), .A(n7745) );
  inv01 U5193 ( .Y(s_expo9_2[2]), .A(n7747) );
  inv01 U5194 ( .Y(s_expo9_2[1]), .A(n7749) );
  mux21 U5195 ( .Y(n7751), .A0(s_expo9_1[0]), .A1(n____return2548_0_), .S0(
        n7667) );
  nor02 U5196 ( .Y(n8016), .A0(s_fracto28_1[27]), .A1(s_fracto28_1[26]) );
  ao21 U5197 ( .Y(s_expo9_11794_6_), .A0(n7706), .A1(n4748), .B0(n8017) );
  ao21 U5198 ( .Y(s_expo9_11794_5_), .A0(n7706), .A1(n8018), .B0(n8017) );
  ao21 U5199 ( .Y(s_expo9_11794_4_), .A0(n7706), .A1(n8019), .B0(n8017) );
  ao21 U5200 ( .Y(s_expo9_11794_3_), .A0(n7706), .A1(n4771), .B0(n8017) );
  ao21 U5201 ( .Y(s_expo9_11794_2_), .A0(n7706), .A1(n8020), .B0(n8017) );
  ao21 U5202 ( .Y(s_expo9_11794_1_), .A0(n7706), .A1(n4730), .B0(n8017) );
  nand02 U5203 ( .Y(n7705), .A0(n7712), .A1(n8022) );
  nand03 U5204 ( .Y(s_expo9_11794_0_), .A0(n8023), .A1(n4778), .A2(n7712) );
  xor2 U5205 ( .Y(n8019), .A0(n8027), .A1(n7387) );
  xor2 U5206 ( .Y(n8018), .A0(n8030), .A1(n8031) );
  xor2 U5207 ( .Y(n8020), .A0(n8033), .A1(n4716) );
  xnor2 U5208 ( .Y(n8021), .A0(n7543), .A1(n8036) );
  xor2 U5209 ( .Y(n8036), .A0(n4720), .A1(n7550) );
  xor2 U5210 ( .Y(n8039), .A0(n7082), .A1(n7542) );
  and02 U5211 ( .Y(n8024), .A0(n7188), .A1(n7190) );
  inv01 U5212 ( .Y(n8041), .A(n8042) );
  nand02 U5213 ( .Y(n8043), .A0(n8044), .A1(exp_i[4]) );
  ao21 U5214 ( .Y(n8045), .A0(n7707), .A1(n7387), .B0(n8029) );
  inv01 U5215 ( .Y(n8029), .A(n8028) );
  ao21 U5216 ( .Y(n8046), .A0(n7542), .A1(n8038), .B0(n7082) );
  inv01 U5217 ( .Y(n8049), .A(n8050) );
  ao21 U5218 ( .Y(n8051), .A0(n7550), .A1(n7544), .B0(n4720) );
  xor2 U5219 ( .Y(n8037), .A0(n8052), .A1(exp_i[1]) );
  nand02 U5220 ( .Y(n8052), .A0(exp_i[0]), .A1(fract_28_i[27]) );
  nor02 U5221 ( .Y(n7794), .A0(n8053), .A1(n8054) );
  nand04 U5222 ( .Y(n8053), .A0(n8068), .A1(n8069), .A2(n8070), .A3(n8071) );
  inv01 U5223 ( .Y(n8074), .A(n6660) );
  nand04 U5224 ( .Y(n8083), .A0(n8068), .A1(n8086), .A2(n8087), .A3(n8088) );
  inv01 U5225 ( .Y(n8089), .A(n7245) );
  nand04 U5226 ( .Y(n8090), .A0(n8094), .A1(n4758), .A2(n8095), .A3(n8096) );
  nand04 U5227 ( .Y(n8098), .A0(n8101), .A1(n4769), .A2(n8100), .A3(n8099) );
  and02 U5228 ( .Y(n8062), .A0(fract_28_i[10]), .A1(n4895) );
  and02 U5229 ( .Y(n8061), .A0(fract_28_i[8]), .A1(n8102) );
  and03 U5230 ( .Y(n8066), .A0(n4513), .A1(n7954), .A2(fract_28_i[6]) );
  and03 U5231 ( .Y(n8076), .A0(n6967), .A1(n7889), .A2(fract_28_i[2]) );
  and02 U5232 ( .Y(n8075), .A0(fract_28_i[16]), .A1(n8105) );
  and02 U5233 ( .Y(n8079), .A0(fract_28_i[14]), .A1(n8106) );
  and03 U5234 ( .Y(n8081), .A0(n4893), .A1(n7980), .A2(fract_28_i[12]) );
  and02 U5235 ( .Y(n8059), .A0(fract_28_i[18]), .A1(n4746) );
  nand03 U5236 ( .Y(n8022), .A0(n8040), .A1(exp_i[6]), .A2(exp_i[7]) );
  inv01 U5237 ( .Y(n8107), .A(exp_i[3]) );
  inv01 U5238 ( .Y(n8047), .A(exp_i[2]) );
  inv01 U5239 ( .Y(n8023), .A(n8032) );
  ao21 U5240 ( .Y(n8032), .A0(n4750), .A1(n8108), .B0(n7544) );
  nor02 U5241 ( .Y(n8035), .A0(n8108), .A1(n4750) );
  inv01 U5242 ( .Y(n8108), .A(n7709) );
  nor02 U5243 ( .Y(n7709), .A0(fract_28_i[27]), .A1(n7795) );
  and04 U5244 ( .Y(n7795), .A0(n8109), .A1(n8110), .A2(n8111), .A3(n8112) );
  and03 U5245 ( .Y(n8063), .A0(n4895), .A1(n7875), .A2(fract_28_i[9]) );
  and02 U5246 ( .Y(n8065), .A0(fract_28_i[7]), .A1(n4513) );
  and02 U5247 ( .Y(n8064), .A0(fract_28_i[5]), .A1(n8104) );
  and03 U5248 ( .Y(n8060), .A0(n4746), .A1(n7949), .A2(fract_28_i[17]) );
  and02 U5249 ( .Y(n8058), .A0(fract_28_i[1]), .A1(n4732) );
  and03 U5250 ( .Y(n8080), .A0(n8072), .A1(n7245), .A2(fract_28_i[19]) );
  and03 U5251 ( .Y(n8103), .A0(n7880), .A1(n7879), .A2(n8104) );
  and03 U5252 ( .Y(n8102), .A0(n7875), .A1(n7873), .A2(n4895) );
  and03 U5253 ( .Y(n8078), .A0(n8105), .A1(n7967), .A2(fract_28_i[15]) );
  and02 U5254 ( .Y(n8077), .A0(fract_28_i[13]), .A1(n4893) );
  and02 U5255 ( .Y(n8082), .A0(fract_28_i[11]), .A1(n8113) );
  and03 U5256 ( .Y(n8113), .A0(n7957), .A1(n7980), .A2(n4893) );
  and03 U5257 ( .Y(n8106), .A0(n7606), .A1(n7967), .A2(n8105) );
  nor02 U5258 ( .Y(n8073), .A0(fract_28_i[26]), .A1(fract_28_i[25]) );
  post_norm_addsub_DW01_inc_9_0 add_188_plus_plus ( .A(s_expo9_2), .SUM({
        n2866_8_, n____return2864_7_, n____return2864_6_, n____return2864_5_, 
        n____return2864_4_, n____return2864_3_, n____return2864_2_, 
        n____return2864_1_, n____return2864_0_}) );
  post_norm_addsub_DW01_add_28_0 add_182_plus_plus ( .A(s_fracto28_1), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b1, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({n2768_27_, 
        n____return2766_26_, n____return2766_25_, n____return2766_24_, 
        n____return2766_23_, n____return2766_22_, n____return2766_21_, 
        n____return2766_20_, n____return2766_19_, n____return2766_18_, 
        n____return2766_17_, n____return2766_16_, n____return2766_15_, 
        n____return2766_14_, n____return2766_13_, n____return2766_12_, 
        n____return2766_11_, n____return2766_10_, n____return2766_9_, 
        n____return2766_8_, n____return2766_7_, n____return2766_6_, 
        n____return2766_5_, n____return2766_4_, n____return2766_3_, 
        n____return2766_2_, n____return2766_1_, n____return2766_0_}) );
  post_norm_addsub_DW01_dec_9_0 sub_172_minus_minus ( .A(s_expo9_1), .SUM({
        n2550_8_, n____return2548_7_, n____return2548_6_, n____return2548_5_, 
        n____return2548_4_, n____return2548_3_, n____return2548_2_, 
        n____return2548_1_, n____return2548_0_}) );
  post_norm_addsub_DW01_dec_6_0 sub_140_minus_minus ( .A(exp_i[5:0]), .SUM({
        n____return1927_5_, n____return1927_4_, n____return1927_3_, 
        n____return1927_2_, n____return1927_1_, n____return1927_0_}) );
endmodule


module pre_norm_mul_DW01_add_10_0 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   carry_7_, carry_6_, carry_5_, carry_4_, carry_3_, carry_2_, n174, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173;

  buf02 U4 ( .Y(n1), .A(A[7]) );
  inv02 U5 ( .Y(n2), .A(n1) );
  or02 U6 ( .Y(n3), .A0(B[1]), .A1(A[1]) );
  inv01 U7 ( .Y(n4), .A(n3) );
  or02 U8 ( .Y(n5), .A0(B[6]), .A1(A[6]) );
  inv01 U9 ( .Y(n6), .A(n5) );
  or02 U10 ( .Y(n7), .A0(B[3]), .A1(A[3]) );
  inv01 U11 ( .Y(n8), .A(n7) );
  or02 U12 ( .Y(n9), .A0(B[5]), .A1(A[5]) );
  inv01 U13 ( .Y(n10), .A(n9) );
  or02 U14 ( .Y(n11), .A0(B[2]), .A1(A[2]) );
  inv01 U15 ( .Y(n12), .A(n11) );
  or02 U16 ( .Y(n13), .A0(A[1]), .A1(n29) );
  inv01 U17 ( .Y(n14), .A(n13) );
  or02 U18 ( .Y(n15), .A0(B[7]), .A1(A[7]) );
  inv01 U19 ( .Y(n16), .A(n15) );
  or02 U20 ( .Y(n17), .A0(A[6]), .A1(carry_6_) );
  inv01 U21 ( .Y(n18), .A(n17) );
  or02 U22 ( .Y(n19), .A0(A[3]), .A1(carry_3_) );
  inv01 U23 ( .Y(n20), .A(n19) );
  or02 U24 ( .Y(n21), .A0(A[2]), .A1(carry_2_) );
  inv01 U25 ( .Y(n22), .A(n21) );
  or02 U26 ( .Y(n23), .A0(A[5]), .A1(n125) );
  inv01 U27 ( .Y(n24), .A(n23) );
  or02 U28 ( .Y(n25), .A0(A[7]), .A1(carry_7_) );
  inv01 U29 ( .Y(n26), .A(n25) );
  buf02 U30 ( .Y(SUM[0]), .A(n174) );
  nand02 U31 ( .Y(n28), .A0(A[0]), .A1(B[0]) );
  inv02 U32 ( .Y(n29), .A(n28) );
  inv01 U33 ( .Y(SUM[7]), .A(n30) );
  inv02 U34 ( .Y(SUM[8]), .A(n31) );
  inv02 U35 ( .Y(n32), .A(B[7]) );
  inv02 U36 ( .Y(n33), .A(carry_7_) );
  nor02 U37 ( .Y(n34), .A0(n32), .A1(n35) );
  nor02 U38 ( .Y(n36), .A0(n2), .A1(n37) );
  nor02 U39 ( .Y(n38), .A0(n33), .A1(n39) );
  nor02 U40 ( .Y(n40), .A0(n33), .A1(n41) );
  nor02 U41 ( .Y(n30), .A0(n42), .A1(n43) );
  nor02 U42 ( .Y(n44), .A0(n2), .A1(n33) );
  nor02 U43 ( .Y(n45), .A0(n32), .A1(n33) );
  nor02 U44 ( .Y(n46), .A0(n32), .A1(n2) );
  nor02 U45 ( .Y(n31), .A0(n46), .A1(n47) );
  inv01 U46 ( .Y(n35), .A(n26) );
  nor02 U47 ( .Y(n48), .A0(B[7]), .A1(carry_7_) );
  inv01 U48 ( .Y(n37), .A(n48) );
  inv01 U49 ( .Y(n39), .A(n16) );
  nor02 U50 ( .Y(n49), .A0(n32), .A1(n2) );
  inv01 U51 ( .Y(n41), .A(n49) );
  nor02 U52 ( .Y(n50), .A0(n34), .A1(n36) );
  inv01 U53 ( .Y(n42), .A(n50) );
  nor02 U54 ( .Y(n51), .A0(n38), .A1(n40) );
  inv01 U55 ( .Y(n43), .A(n51) );
  nor02 U56 ( .Y(n52), .A0(n44), .A1(n45) );
  inv01 U57 ( .Y(n47), .A(n52) );
  inv02 U58 ( .Y(SUM[3]), .A(n53) );
  inv02 U59 ( .Y(carry_4_), .A(n54) );
  inv02 U60 ( .Y(n55), .A(B[3]) );
  inv02 U61 ( .Y(n56), .A(A[3]) );
  inv02 U62 ( .Y(n57), .A(carry_3_) );
  nor02 U63 ( .Y(n58), .A0(n55), .A1(n59) );
  nor02 U64 ( .Y(n60), .A0(n56), .A1(n61) );
  nor02 U65 ( .Y(n62), .A0(n57), .A1(n63) );
  nor02 U66 ( .Y(n64), .A0(n57), .A1(n65) );
  nor02 U67 ( .Y(n53), .A0(n66), .A1(n67) );
  nor02 U68 ( .Y(n68), .A0(n56), .A1(n57) );
  nor02 U69 ( .Y(n69), .A0(n55), .A1(n57) );
  nor02 U70 ( .Y(n70), .A0(n55), .A1(n56) );
  nor02 U71 ( .Y(n54), .A0(n70), .A1(n71) );
  inv01 U72 ( .Y(n59), .A(n20) );
  nor02 U73 ( .Y(n72), .A0(B[3]), .A1(carry_3_) );
  inv01 U74 ( .Y(n61), .A(n72) );
  inv01 U75 ( .Y(n63), .A(n8) );
  nor02 U76 ( .Y(n73), .A0(n55), .A1(n56) );
  inv01 U77 ( .Y(n65), .A(n73) );
  nor02 U78 ( .Y(n74), .A0(n58), .A1(n60) );
  inv01 U79 ( .Y(n66), .A(n74) );
  nor02 U80 ( .Y(n75), .A0(n62), .A1(n64) );
  inv01 U81 ( .Y(n67), .A(n75) );
  nor02 U82 ( .Y(n76), .A0(n68), .A1(n69) );
  inv01 U83 ( .Y(n71), .A(n76) );
  inv02 U84 ( .Y(SUM[2]), .A(n77) );
  inv02 U85 ( .Y(carry_3_), .A(n78) );
  inv02 U86 ( .Y(n79), .A(B[2]) );
  inv02 U87 ( .Y(n80), .A(A[2]) );
  inv02 U88 ( .Y(n81), .A(carry_2_) );
  nor02 U89 ( .Y(n82), .A0(n79), .A1(n83) );
  nor02 U90 ( .Y(n84), .A0(n80), .A1(n85) );
  nor02 U91 ( .Y(n86), .A0(n81), .A1(n87) );
  nor02 U92 ( .Y(n88), .A0(n81), .A1(n89) );
  nor02 U93 ( .Y(n77), .A0(n90), .A1(n91) );
  nor02 U94 ( .Y(n92), .A0(n80), .A1(n81) );
  nor02 U95 ( .Y(n93), .A0(n79), .A1(n81) );
  nor02 U96 ( .Y(n94), .A0(n79), .A1(n80) );
  nor02 U97 ( .Y(n78), .A0(n94), .A1(n95) );
  inv01 U98 ( .Y(n83), .A(n22) );
  nor02 U99 ( .Y(n96), .A0(B[2]), .A1(carry_2_) );
  inv01 U100 ( .Y(n85), .A(n96) );
  inv01 U101 ( .Y(n87), .A(n12) );
  nor02 U102 ( .Y(n97), .A0(n79), .A1(n80) );
  inv01 U103 ( .Y(n89), .A(n97) );
  nor02 U104 ( .Y(n98), .A0(n82), .A1(n84) );
  inv01 U105 ( .Y(n90), .A(n98) );
  nor02 U106 ( .Y(n99), .A0(n86), .A1(n88) );
  inv01 U107 ( .Y(n91), .A(n99) );
  nor02 U108 ( .Y(n100), .A0(n92), .A1(n93) );
  inv01 U109 ( .Y(n95), .A(n100) );
  inv02 U110 ( .Y(SUM[6]), .A(n101) );
  inv02 U111 ( .Y(carry_7_), .A(n102) );
  inv02 U112 ( .Y(n103), .A(B[6]) );
  inv02 U113 ( .Y(n104), .A(A[6]) );
  inv02 U114 ( .Y(n105), .A(carry_6_) );
  nor02 U115 ( .Y(n106), .A0(n103), .A1(n107) );
  nor02 U116 ( .Y(n108), .A0(n104), .A1(n109) );
  nor02 U117 ( .Y(n110), .A0(n105), .A1(n111) );
  nor02 U118 ( .Y(n112), .A0(n105), .A1(n113) );
  nor02 U119 ( .Y(n101), .A0(n114), .A1(n115) );
  nor02 U120 ( .Y(n116), .A0(n104), .A1(n105) );
  nor02 U121 ( .Y(n117), .A0(n103), .A1(n105) );
  nor02 U122 ( .Y(n118), .A0(n103), .A1(n104) );
  nor02 U123 ( .Y(n102), .A0(n118), .A1(n119) );
  inv01 U124 ( .Y(n107), .A(n18) );
  nor02 U125 ( .Y(n120), .A0(B[6]), .A1(carry_6_) );
  inv01 U126 ( .Y(n109), .A(n120) );
  inv01 U127 ( .Y(n111), .A(n6) );
  nor02 U128 ( .Y(n121), .A0(n103), .A1(n104) );
  inv01 U129 ( .Y(n113), .A(n121) );
  nor02 U130 ( .Y(n122), .A0(n106), .A1(n108) );
  inv01 U131 ( .Y(n114), .A(n122) );
  nor02 U132 ( .Y(n123), .A0(n110), .A1(n112) );
  inv01 U133 ( .Y(n115), .A(n123) );
  nor02 U134 ( .Y(n124), .A0(n116), .A1(n117) );
  inv01 U135 ( .Y(n119), .A(n124) );
  buf02 U136 ( .Y(n125), .A(carry_5_) );
  inv02 U137 ( .Y(SUM[1]), .A(n126) );
  inv02 U138 ( .Y(carry_2_), .A(n127) );
  inv02 U139 ( .Y(n128), .A(B[1]) );
  inv02 U140 ( .Y(n129), .A(A[1]) );
  inv02 U141 ( .Y(n130), .A(n29) );
  nor02 U142 ( .Y(n131), .A0(n128), .A1(n132) );
  nor02 U143 ( .Y(n133), .A0(n129), .A1(n134) );
  nor02 U144 ( .Y(n135), .A0(n130), .A1(n136) );
  nor02 U145 ( .Y(n137), .A0(n130), .A1(n138) );
  nor02 U146 ( .Y(n126), .A0(n139), .A1(n140) );
  nor02 U147 ( .Y(n141), .A0(n129), .A1(n130) );
  nor02 U148 ( .Y(n142), .A0(n128), .A1(n130) );
  nor02 U149 ( .Y(n143), .A0(n128), .A1(n129) );
  nor02 U150 ( .Y(n127), .A0(n143), .A1(n144) );
  inv01 U151 ( .Y(n132), .A(n14) );
  nor02 U152 ( .Y(n145), .A0(B[1]), .A1(n29) );
  inv01 U153 ( .Y(n134), .A(n145) );
  inv01 U154 ( .Y(n136), .A(n4) );
  nor02 U155 ( .Y(n146), .A0(n128), .A1(n129) );
  inv01 U156 ( .Y(n138), .A(n146) );
  nor02 U157 ( .Y(n147), .A0(n131), .A1(n133) );
  inv01 U158 ( .Y(n139), .A(n147) );
  nor02 U159 ( .Y(n148), .A0(n135), .A1(n137) );
  inv01 U160 ( .Y(n140), .A(n148) );
  nor02 U161 ( .Y(n149), .A0(n141), .A1(n142) );
  inv01 U162 ( .Y(n144), .A(n149) );
  inv02 U163 ( .Y(SUM[5]), .A(n150) );
  inv02 U164 ( .Y(carry_6_), .A(n151) );
  inv02 U165 ( .Y(n152), .A(B[5]) );
  inv02 U166 ( .Y(n153), .A(A[5]) );
  inv02 U167 ( .Y(n154), .A(n125) );
  nor02 U168 ( .Y(n155), .A0(n152), .A1(n156) );
  nor02 U169 ( .Y(n157), .A0(n153), .A1(n158) );
  nor02 U170 ( .Y(n159), .A0(n154), .A1(n160) );
  nor02 U171 ( .Y(n161), .A0(n154), .A1(n162) );
  nor02 U172 ( .Y(n150), .A0(n163), .A1(n164) );
  nor02 U173 ( .Y(n165), .A0(n153), .A1(n154) );
  nor02 U174 ( .Y(n166), .A0(n152), .A1(n154) );
  nor02 U175 ( .Y(n167), .A0(n152), .A1(n153) );
  nor02 U176 ( .Y(n151), .A0(n167), .A1(n168) );
  inv01 U177 ( .Y(n156), .A(n24) );
  nor02 U178 ( .Y(n169), .A0(B[5]), .A1(n125) );
  inv01 U179 ( .Y(n158), .A(n169) );
  inv01 U180 ( .Y(n160), .A(n10) );
  nor02 U181 ( .Y(n170), .A0(n152), .A1(n153) );
  inv01 U182 ( .Y(n162), .A(n170) );
  nor02 U183 ( .Y(n171), .A0(n155), .A1(n157) );
  inv01 U184 ( .Y(n163), .A(n171) );
  nor02 U185 ( .Y(n172), .A0(n159), .A1(n161) );
  inv01 U186 ( .Y(n164), .A(n172) );
  nor02 U187 ( .Y(n173), .A0(n165), .A1(n166) );
  inv01 U188 ( .Y(n168), .A(n173) );
  xor2 U189 ( .Y(n174), .A0(B[0]), .A1(A[0]) );
  fadd1 U1_4 ( .S(SUM[4]), .CO(carry_5_), .A(A[4]), .B(B[4]), .CI(carry_4_) );
endmodule


module pre_norm_mul ( clk_i, opa_i, opb_i, exp_10_o, fracta_24_o, fractb_24_o
 );
  input [31:0] opa_i;
  input [31:0] opb_i;
  output [9:0] exp_10_o;
  output [23:0] fracta_24_o;
  output [23:0] fractb_24_o;
  input clk_i;
  wire   opa_i_22_, opa_i_21_, opa_i_20_, opa_i_19_, opa_i_18_, opa_i_17_,
         opa_i_16_, opa_i_15_, opa_i_14_, opa_i_13_, opa_i_12_, opa_i_11_,
         opa_i_10_, opa_i_9_, opa_i_8_, opa_i_7_, opa_i_6_, opa_i_5_, opa_i_4_,
         opa_i_3_, opa_i_2_, opa_i_1_, opa_i_0_, opb_i_22_, opb_i_21_,
         opb_i_20_, opb_i_19_, opb_i_18_, opb_i_17_, opb_i_16_, opb_i_15_,
         opb_i_14_, opb_i_13_, opb_i_12_, opb_i_11_, opb_i_10_, opb_i_9_,
         opb_i_8_, opb_i_7_, opb_i_6_, opb_i_5_, opb_i_4_, opb_i_3_, opb_i_2_,
         opb_i_1_, opb_i_0_, s_exp_10_o_9_, s_exp_10_o_7_, s_exp_10_o_5_,
         s_exp_10_o_0_, n386, n387, s_expa_in_0_, s_expb_in_0_,
         n____return225_8_, n____return225_7_, n____return225_6_,
         n____return225_5_, n____return225_4_, n____return225_3_,
         n____return225_2_, n____return225_1_, n____return225_0_, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n361, n363, n364, n365, n366, n367, n368, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, SYNOPSYS_UNCONNECTED_1;
  assign fracta_24_o[22] = opa_i_22_;
  assign opa_i_22_ = opa_i[22];
  assign fracta_24_o[21] = opa_i_21_;
  assign opa_i_21_ = opa_i[21];
  assign fracta_24_o[20] = opa_i_20_;
  assign opa_i_20_ = opa_i[20];
  assign fracta_24_o[19] = opa_i_19_;
  assign opa_i_19_ = opa_i[19];
  assign fracta_24_o[18] = opa_i_18_;
  assign opa_i_18_ = opa_i[18];
  assign fracta_24_o[17] = opa_i_17_;
  assign opa_i_17_ = opa_i[17];
  assign fracta_24_o[16] = opa_i_16_;
  assign opa_i_16_ = opa_i[16];
  assign fracta_24_o[15] = opa_i_15_;
  assign opa_i_15_ = opa_i[15];
  assign fracta_24_o[14] = opa_i_14_;
  assign opa_i_14_ = opa_i[14];
  assign fracta_24_o[13] = opa_i_13_;
  assign opa_i_13_ = opa_i[13];
  assign fracta_24_o[12] = opa_i_12_;
  assign opa_i_12_ = opa_i[12];
  assign fracta_24_o[11] = opa_i_11_;
  assign opa_i_11_ = opa_i[11];
  assign fracta_24_o[10] = opa_i_10_;
  assign opa_i_10_ = opa_i[10];
  assign fracta_24_o[9] = opa_i_9_;
  assign opa_i_9_ = opa_i[9];
  assign fracta_24_o[8] = opa_i_8_;
  assign opa_i_8_ = opa_i[8];
  assign fracta_24_o[7] = opa_i_7_;
  assign opa_i_7_ = opa_i[7];
  assign fracta_24_o[6] = opa_i_6_;
  assign opa_i_6_ = opa_i[6];
  assign fracta_24_o[5] = opa_i_5_;
  assign opa_i_5_ = opa_i[5];
  assign fracta_24_o[4] = opa_i_4_;
  assign opa_i_4_ = opa_i[4];
  assign fracta_24_o[3] = opa_i_3_;
  assign opa_i_3_ = opa_i[3];
  assign fracta_24_o[2] = opa_i_2_;
  assign opa_i_2_ = opa_i[2];
  assign fracta_24_o[1] = opa_i_1_;
  assign opa_i_1_ = opa_i[1];
  assign fracta_24_o[0] = opa_i_0_;
  assign opa_i_0_ = opa_i[0];
  assign fractb_24_o[22] = opb_i_22_;
  assign opb_i_22_ = opb_i[22];
  assign fractb_24_o[21] = opb_i_21_;
  assign opb_i_21_ = opb_i[21];
  assign fractb_24_o[20] = opb_i_20_;
  assign opb_i_20_ = opb_i[20];
  assign fractb_24_o[19] = opb_i_19_;
  assign opb_i_19_ = opb_i[19];
  assign fractb_24_o[18] = opb_i_18_;
  assign opb_i_18_ = opb_i[18];
  assign fractb_24_o[17] = opb_i_17_;
  assign opb_i_17_ = opb_i[17];
  assign fractb_24_o[16] = opb_i_16_;
  assign opb_i_16_ = opb_i[16];
  assign fractb_24_o[15] = opb_i_15_;
  assign opb_i_15_ = opb_i[15];
  assign fractb_24_o[14] = opb_i_14_;
  assign opb_i_14_ = opb_i[14];
  assign fractb_24_o[13] = opb_i_13_;
  assign opb_i_13_ = opb_i[13];
  assign fractb_24_o[12] = opb_i_12_;
  assign opb_i_12_ = opb_i[12];
  assign fractb_24_o[11] = opb_i_11_;
  assign opb_i_11_ = opb_i[11];
  assign fractb_24_o[10] = opb_i_10_;
  assign opb_i_10_ = opb_i[10];
  assign fractb_24_o[9] = opb_i_9_;
  assign opb_i_9_ = opb_i[9];
  assign fractb_24_o[8] = opb_i_8_;
  assign opb_i_8_ = opb_i[8];
  assign fractb_24_o[7] = opb_i_7_;
  assign opb_i_7_ = opb_i[7];
  assign fractb_24_o[6] = opb_i_6_;
  assign opb_i_6_ = opb_i[6];
  assign fractb_24_o[5] = opb_i_5_;
  assign opb_i_5_ = opb_i[5];
  assign fractb_24_o[4] = opb_i_4_;
  assign opb_i_4_ = opb_i[4];
  assign fractb_24_o[3] = opb_i_3_;
  assign opb_i_3_ = opb_i[3];
  assign fractb_24_o[2] = opb_i_2_;
  assign opb_i_2_ = opb_i[2];
  assign fractb_24_o[1] = opb_i_1_;
  assign opb_i_1_ = opb_i[1];
  assign fractb_24_o[0] = opb_i_0_;
  assign opb_i_0_ = opb_i[0];

  dff exp_10_o_reg_9_ ( .Q(exp_10_o[9]), .D(s_exp_10_o_9_), .CLK(clk_i) );
  dff exp_10_o_reg_8_ ( .Q(exp_10_o[8]), .D(n310), .CLK(clk_i) );
  dff exp_10_o_reg_7_ ( .Q(exp_10_o[7]), .D(s_exp_10_o_7_), .CLK(clk_i) );
  dff exp_10_o_reg_6_ ( .Q(exp_10_o[6]), .D(n314), .CLK(clk_i) );
  dff exp_10_o_reg_5_ ( .Q(exp_10_o[5]), .D(s_exp_10_o_5_), .CLK(clk_i) );
  dff exp_10_o_reg_4_ ( .Q(exp_10_o[4]), .D(n316), .CLK(clk_i) );
  dff exp_10_o_reg_3_ ( .Q(exp_10_o[3]), .D(n306), .CLK(clk_i) );
  dff exp_10_o_reg_2_ ( .Q(exp_10_o[2]), .D(n308), .CLK(clk_i) );
  dff exp_10_o_reg_1_ ( .Q(exp_10_o[1]), .D(n312), .CLK(clk_i) );
  dff exp_10_o_reg_0_ ( .Q(exp_10_o[0]), .D(s_exp_10_o_0_), .CLK(clk_i) );
  buf02 U42 ( .Y(n301), .A(s_expb_in_0_) );
  buf02 U43 ( .Y(n302), .A(s_expa_in_0_) );
  or02 U44 ( .Y(n303), .A0(n379), .A1(n378) );
  inv01 U45 ( .Y(n304), .A(n303) );
  xor2 U46 ( .Y(n305), .A0(n____return225_3_), .A1(n379) );
  inv01 U47 ( .Y(n306), .A(n305) );
  xor2 U48 ( .Y(n307), .A0(n____return225_2_), .A1(n381) );
  inv01 U49 ( .Y(n308), .A(n307) );
  xor2 U50 ( .Y(n309), .A0(n____return225_8_), .A1(n373) );
  inv01 U51 ( .Y(n310), .A(n309) );
  xor2 U52 ( .Y(n311), .A0(s_exp_10_o_0_), .A1(n____return225_1_) );
  inv01 U53 ( .Y(n312), .A(n311) );
  xor2 U54 ( .Y(n313), .A0(n____return225_6_), .A1(n377) );
  inv01 U55 ( .Y(n314), .A(n313) );
  xor2 U56 ( .Y(n315), .A0(n304), .A1(n380) );
  inv01 U57 ( .Y(n316), .A(n315) );
  inv01 U58 ( .Y(n317), .A(n373) );
  inv02 U59 ( .Y(n373), .A(n374) );
  inv01 U60 ( .Y(n382), .A(n318) );
  inv01 U61 ( .Y(n319), .A(opb_i[23]) );
  inv01 U62 ( .Y(n320), .A(opb_i[24]) );
  inv01 U63 ( .Y(n321), .A(opb_i[25]) );
  inv01 U64 ( .Y(n322), .A(opb_i[26]) );
  nand02 U65 ( .Y(n318), .A0(n323), .A1(n324) );
  nand02 U66 ( .Y(n325), .A0(n319), .A1(n320) );
  inv01 U67 ( .Y(n323), .A(n325) );
  nand02 U68 ( .Y(n326), .A0(n321), .A1(n322) );
  inv01 U69 ( .Y(n324), .A(n326) );
  inv01 U70 ( .Y(n383), .A(n327) );
  inv01 U71 ( .Y(n328), .A(opb_i[27]) );
  inv01 U72 ( .Y(n329), .A(opb_i[28]) );
  inv01 U73 ( .Y(n330), .A(opb_i[29]) );
  inv01 U74 ( .Y(n331), .A(opb_i[30]) );
  nand02 U75 ( .Y(n327), .A0(n332), .A1(n333) );
  nand02 U76 ( .Y(n334), .A0(n328), .A1(n329) );
  inv01 U77 ( .Y(n332), .A(n334) );
  nand02 U78 ( .Y(n335), .A0(n330), .A1(n331) );
  inv01 U79 ( .Y(n333), .A(n335) );
  inv02 U80 ( .Y(n379), .A(n336) );
  inv01 U81 ( .Y(n337), .A(n____return225_2_) );
  inv01 U82 ( .Y(n338), .A(n____return225_0_) );
  inv01 U83 ( .Y(n339), .A(n____return225_1_) );
  nor02 U84 ( .Y(n336), .A0(n339), .A1(n340) );
  nor02 U85 ( .Y(n341), .A0(n337), .A1(n338) );
  inv01 U86 ( .Y(n340), .A(n341) );
  inv02 U87 ( .Y(s_exp_10_o_0_), .A(n____return225_0_) );
  inv01 U88 ( .Y(n385), .A(n342) );
  inv01 U89 ( .Y(n343), .A(opa_i[27]) );
  inv01 U90 ( .Y(n344), .A(opa_i[28]) );
  inv01 U91 ( .Y(n345), .A(opa_i[29]) );
  inv01 U92 ( .Y(n346), .A(opa_i[30]) );
  nand02 U93 ( .Y(n342), .A0(n347), .A1(n348) );
  nand02 U94 ( .Y(n349), .A0(n343), .A1(n344) );
  inv01 U95 ( .Y(n347), .A(n349) );
  nand02 U96 ( .Y(n350), .A0(n345), .A1(n346) );
  inv01 U97 ( .Y(n348), .A(n350) );
  inv01 U98 ( .Y(n384), .A(n351) );
  inv01 U99 ( .Y(n352), .A(opa_i[23]) );
  inv01 U100 ( .Y(n353), .A(opa_i[24]) );
  inv01 U101 ( .Y(n354), .A(opa_i[25]) );
  inv01 U102 ( .Y(n355), .A(opa_i[26]) );
  nand02 U103 ( .Y(n351), .A0(n356), .A1(n357) );
  nand02 U104 ( .Y(n358), .A0(n352), .A1(n353) );
  inv01 U105 ( .Y(n356), .A(n358) );
  nand02 U106 ( .Y(n359), .A0(n354), .A1(n355) );
  inv01 U107 ( .Y(n357), .A(n359) );
  buf02 U108 ( .Y(fractb_24_o[23]), .A(n387) );
  buf02 U109 ( .Y(n361), .A(n387) );
  buf02 U110 ( .Y(fracta_24_o[23]), .A(n386) );
  inv02 U111 ( .Y(n376), .A(n363) );
  inv01 U112 ( .Y(n364), .A(n380) );
  inv01 U113 ( .Y(n365), .A(n379) );
  inv01 U114 ( .Y(n366), .A(n378) );
  nand02 U115 ( .Y(n363), .A0(n366), .A1(n367) );
  nand02 U116 ( .Y(n368), .A0(n364), .A1(n365) );
  inv01 U117 ( .Y(n367), .A(n368) );
  inv02 U118 ( .Y(n380), .A(n____return225_4_) );
  inv01 U119 ( .Y(s_exp_10_o_9_), .A(n372) );
  nand02 U120 ( .Y(s_expb_in_0_), .A0(n361), .A1(n370) );
  inv01 U121 ( .Y(n370), .A(opb_i[23]) );
  nand02 U123 ( .Y(s_expa_in_0_), .A0(fracta_24_o[23]), .A1(n371) );
  inv01 U124 ( .Y(n371), .A(opa_i[23]) );
  or02 U125 ( .Y(n372), .A0(n373), .A1(n____return225_8_) );
  ao21 U126 ( .Y(s_exp_10_o_7_), .A0(n____return225_7_), .A1(n375), .B0(n317)
         );
  nor02 U127 ( .Y(n374), .A0(n____return225_7_), .A1(n375) );
  and03 U128 ( .Y(n375), .A0(n____return225_5_), .A1(n376), .A2(
        n____return225_6_) );
  nand02 U129 ( .Y(n377), .A0(n____return225_5_), .A1(n376) );
  xor2 U130 ( .Y(s_exp_10_o_5_), .A0(n376), .A1(n____return225_5_) );
  inv01 U131 ( .Y(n378), .A(n____return225_3_) );
  nand02 U132 ( .Y(n381), .A0(n____return225_1_), .A1(n____return225_0_) );
  nand02 U133 ( .Y(n387), .A0(n382), .A1(n383) );
  nand02 U134 ( .Y(n386), .A0(n384), .A1(n385) );
  pre_norm_mul_DW01_add_10_0 add_1_root_sub_101_minus_minus ( .A({1'b0, 1'b0, 
        opa_i[30:24], n302}), .B({1'b0, 1'b0, opb_i[30:24], n301}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED_1, n____return225_8_, n____return225_7_, 
        n____return225_6_, n____return225_5_, n____return225_4_, 
        n____return225_3_, n____return225_2_, n____return225_1_, 
        n____return225_0_}) );
endmodule


module post_norm_mul_DW01_inc_9_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;
  wire   carry_8_, carry_7_, carry_6_, carry_5_, carry_4_, carry_3_, carry_2_;

  inv01 U5 ( .Y(SUM[0]), .A(A[0]) );
  xor2 U6 ( .Y(SUM[8]), .A0(carry_8_), .A1(A[8]) );
  hadd1 U1_1_1 ( .S(SUM[1]), .CO(carry_2_), .A(A[1]), .B(A[0]) );
  hadd1 U1_1_2 ( .S(SUM[2]), .CO(carry_3_), .A(A[2]), .B(carry_2_) );
  hadd1 U1_1_3 ( .S(SUM[3]), .CO(carry_4_), .A(A[3]), .B(carry_3_) );
  hadd1 U1_1_4 ( .S(SUM[4]), .CO(carry_5_), .A(A[4]), .B(carry_4_) );
  hadd1 U1_1_5 ( .S(SUM[5]), .CO(carry_6_), .A(A[5]), .B(carry_5_) );
  hadd1 U1_1_6 ( .S(SUM[6]), .CO(carry_7_), .A(A[6]), .B(carry_6_) );
  hadd1 U1_1_7 ( .S(SUM[7]), .CO(carry_8_), .A(A[7]), .B(carry_7_) );
endmodule


module post_norm_mul_DW01_inc_25_0 ( A, SUM );
  input [24:0] A;
  output [24:0] SUM;
  wire   carry_24_, carry_23_, carry_22_, carry_21_, carry_20_, carry_19_,
         carry_18_, carry_17_, carry_16_, carry_15_, carry_14_, carry_13_,
         carry_12_, carry_11_, carry_10_, carry_9_, carry_8_, carry_7_,
         carry_6_, carry_5_, carry_4_, carry_3_, carry_2_;

  inv04 U5 ( .Y(SUM[0]), .A(A[0]) );
  xor2 U6 ( .Y(SUM[24]), .A0(carry_24_), .A1(A[24]) );
  hadd1 U1_1_1 ( .S(SUM[1]), .CO(carry_2_), .A(A[1]), .B(A[0]) );
  hadd1 U1_1_2 ( .S(SUM[2]), .CO(carry_3_), .A(A[2]), .B(carry_2_) );
  hadd1 U1_1_3 ( .S(SUM[3]), .CO(carry_4_), .A(A[3]), .B(carry_3_) );
  hadd1 U1_1_4 ( .S(SUM[4]), .CO(carry_5_), .A(A[4]), .B(carry_4_) );
  hadd1 U1_1_5 ( .S(SUM[5]), .CO(carry_6_), .A(A[5]), .B(carry_5_) );
  hadd1 U1_1_6 ( .S(SUM[6]), .CO(carry_7_), .A(A[6]), .B(carry_6_) );
  hadd1 U1_1_7 ( .S(SUM[7]), .CO(carry_8_), .A(A[7]), .B(carry_7_) );
  hadd1 U1_1_8 ( .S(SUM[8]), .CO(carry_9_), .A(A[8]), .B(carry_8_) );
  hadd1 U1_1_9 ( .S(SUM[9]), .CO(carry_10_), .A(A[9]), .B(carry_9_) );
  hadd1 U1_1_10 ( .S(SUM[10]), .CO(carry_11_), .A(A[10]), .B(carry_10_) );
  hadd1 U1_1_11 ( .S(SUM[11]), .CO(carry_12_), .A(A[11]), .B(carry_11_) );
  hadd1 U1_1_12 ( .S(SUM[12]), .CO(carry_13_), .A(A[12]), .B(carry_12_) );
  hadd1 U1_1_13 ( .S(SUM[13]), .CO(carry_14_), .A(A[13]), .B(carry_13_) );
  hadd1 U1_1_14 ( .S(SUM[14]), .CO(carry_15_), .A(A[14]), .B(carry_14_) );
  hadd1 U1_1_15 ( .S(SUM[15]), .CO(carry_16_), .A(A[15]), .B(carry_15_) );
  hadd1 U1_1_16 ( .S(SUM[16]), .CO(carry_17_), .A(A[16]), .B(carry_16_) );
  hadd1 U1_1_17 ( .S(SUM[17]), .CO(carry_18_), .A(A[17]), .B(carry_17_) );
  hadd1 U1_1_18 ( .S(SUM[18]), .CO(carry_19_), .A(A[18]), .B(carry_18_) );
  hadd1 U1_1_19 ( .S(SUM[19]), .CO(carry_20_), .A(A[19]), .B(carry_19_) );
  hadd1 U1_1_20 ( .S(SUM[20]), .CO(carry_21_), .A(A[20]), .B(carry_20_) );
  hadd1 U1_1_21 ( .S(SUM[21]), .CO(carry_22_), .A(A[21]), .B(carry_21_) );
  hadd1 U1_1_22 ( .S(SUM[22]), .CO(carry_23_), .A(A[22]), .B(carry_22_) );
  hadd1 U1_1_23 ( .S(SUM[23]), .CO(carry_24_), .A(A[23]), .B(carry_23_) );
endmodule


module post_norm_mul_DW01_dec_9_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;
  wire   carry_8_, carry_7_, carry_6_, carry_5_, carry_4_, carry_3_, carry_2_,
         n5, n7, n9, n11, n13, n15, n17, n19, n21, n22, n23, n24, n25, n26;

  xor2 U6 ( .Y(n5), .A0(A[1]), .A1(A[0]) );
  inv01 U7 ( .Y(SUM[1]), .A(n5) );
  xor2 U8 ( .Y(n7), .A0(A[5]), .A1(n26) );
  inv01 U9 ( .Y(SUM[5]), .A(n7) );
  xor2 U10 ( .Y(n9), .A0(A[4]), .A1(n25) );
  inv01 U11 ( .Y(SUM[4]), .A(n9) );
  xor2 U12 ( .Y(n11), .A0(A[6]), .A1(n21) );
  inv01 U13 ( .Y(SUM[6]), .A(n11) );
  xor2 U14 ( .Y(n13), .A0(A[7]), .A1(n23) );
  inv01 U15 ( .Y(SUM[7]), .A(n13) );
  xor2 U16 ( .Y(n15), .A0(carry_8_), .A1(A[8]) );
  inv01 U17 ( .Y(SUM[8]), .A(n15) );
  xor2 U18 ( .Y(n17), .A0(A[2]), .A1(n22) );
  inv01 U19 ( .Y(SUM[2]), .A(n17) );
  xor2 U20 ( .Y(n19), .A0(A[3]), .A1(n24) );
  inv01 U21 ( .Y(SUM[3]), .A(n19) );
  buf02 U22 ( .Y(n21), .A(carry_6_) );
  buf02 U23 ( .Y(n22), .A(carry_2_) );
  buf02 U24 ( .Y(n23), .A(carry_7_) );
  buf02 U25 ( .Y(n24), .A(carry_3_) );
  buf02 U26 ( .Y(n25), .A(carry_4_) );
  buf02 U27 ( .Y(n26), .A(carry_5_) );
  inv01 U28 ( .Y(SUM[0]), .A(A[0]) );
  or02 U1_B_1 ( .Y(carry_2_), .A0(A[1]), .A1(A[0]) );
  or02 U1_B_2 ( .Y(carry_3_), .A0(A[2]), .A1(n22) );
  or02 U1_B_3 ( .Y(carry_4_), .A0(A[3]), .A1(n24) );
  or02 U1_B_4 ( .Y(carry_5_), .A0(A[4]), .A1(n25) );
  or02 U1_B_5 ( .Y(carry_6_), .A0(A[5]), .A1(n26) );
  or02 U1_B_6 ( .Y(carry_7_), .A0(A[6]), .A1(n21) );
  or02 U1_B_7 ( .Y(carry_8_), .A0(A[7]), .A1(n23) );
endmodule


module post_norm_mul_DW01_sub_7_0 ( A, B, CI, DIFF, CO );
  input [6:0] A;
  input [6:0] B;
  output [6:0] DIFF;
  input CI;
  output CO;
  wire   carry_6_, carry_5_, carry_4_, carry_3_, carry_2_, carry_1_, n135, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134;
  wire   [6:0] B_not;

  inv02 U6 ( .Y(DIFF[2]), .A(n57) );
  inv02 U7 ( .Y(B_not[6]), .A(B[6]) );
  nand02 U8 ( .Y(DIFF[5]), .A0(n5), .A1(n6) );
  nand02 U9 ( .Y(carry_6_), .A0(n7), .A1(n8) );
  inv01 U10 ( .Y(n9), .A(carry_5_) );
  inv01 U11 ( .Y(n10), .A(A[5]) );
  inv01 U12 ( .Y(n11), .A(B_not[5]) );
  nand02 U13 ( .Y(n12), .A0(n10), .A1(n13) );
  nand02 U14 ( .Y(n14), .A0(n11), .A1(n15) );
  nand02 U15 ( .Y(n16), .A0(n11), .A1(n17) );
  nand02 U16 ( .Y(n18), .A0(carry_5_), .A1(n19) );
  nand02 U17 ( .Y(n20), .A0(A[5]), .A1(carry_5_) );
  nand02 U18 ( .Y(n21), .A0(B_not[5]), .A1(carry_5_) );
  nand02 U19 ( .Y(n7), .A0(B_not[5]), .A1(A[5]) );
  nand02 U20 ( .Y(n22), .A0(B_not[5]), .A1(n9) );
  inv01 U21 ( .Y(n13), .A(n22) );
  nand02 U22 ( .Y(n23), .A0(A[5]), .A1(n9) );
  inv01 U23 ( .Y(n15), .A(n23) );
  nand02 U24 ( .Y(n24), .A0(carry_5_), .A1(n10) );
  inv01 U25 ( .Y(n17), .A(n24) );
  nand02 U26 ( .Y(n25), .A0(B_not[5]), .A1(A[5]) );
  inv01 U27 ( .Y(n19), .A(n25) );
  nand02 U28 ( .Y(n26), .A0(n12), .A1(n14) );
  inv01 U29 ( .Y(n5), .A(n26) );
  nand02 U30 ( .Y(n27), .A0(n16), .A1(n18) );
  inv01 U31 ( .Y(n6), .A(n27) );
  nand02 U32 ( .Y(n28), .A0(n20), .A1(n21) );
  inv01 U33 ( .Y(n8), .A(n28) );
  inv02 U34 ( .Y(B_not[5]), .A(B[5]) );
  buf02 U35 ( .Y(DIFF[0]), .A(n135) );
  inv01 U36 ( .Y(DIFF[4]), .A(n30) );
  inv02 U37 ( .Y(carry_5_), .A(n31) );
  inv02 U38 ( .Y(n32), .A(B_not[4]) );
  inv02 U39 ( .Y(n33), .A(A[4]) );
  inv02 U40 ( .Y(n34), .A(carry_4_) );
  nor02 U41 ( .Y(n35), .A0(n32), .A1(n36) );
  nor02 U42 ( .Y(n37), .A0(n33), .A1(n38) );
  nor02 U43 ( .Y(n39), .A0(n34), .A1(n40) );
  nor02 U44 ( .Y(n41), .A0(n34), .A1(n42) );
  nor02 U45 ( .Y(n30), .A0(n43), .A1(n44) );
  nor02 U46 ( .Y(n45), .A0(n33), .A1(n34) );
  nor02 U47 ( .Y(n46), .A0(n32), .A1(n34) );
  nor02 U48 ( .Y(n47), .A0(n32), .A1(n33) );
  nor02 U49 ( .Y(n31), .A0(n47), .A1(n48) );
  nor02 U50 ( .Y(n49), .A0(A[4]), .A1(carry_4_) );
  inv01 U51 ( .Y(n36), .A(n49) );
  nor02 U52 ( .Y(n50), .A0(B_not[4]), .A1(carry_4_) );
  inv01 U53 ( .Y(n38), .A(n50) );
  nor02 U54 ( .Y(n51), .A0(B_not[4]), .A1(A[4]) );
  inv01 U55 ( .Y(n40), .A(n51) );
  nor02 U56 ( .Y(n52), .A0(n32), .A1(n33) );
  inv01 U57 ( .Y(n42), .A(n52) );
  nor02 U58 ( .Y(n53), .A0(n35), .A1(n37) );
  inv01 U59 ( .Y(n43), .A(n53) );
  nor02 U60 ( .Y(n54), .A0(n39), .A1(n41) );
  inv01 U61 ( .Y(n44), .A(n54) );
  nor02 U62 ( .Y(n55), .A0(n45), .A1(n46) );
  inv01 U63 ( .Y(n48), .A(n55) );
  inv02 U64 ( .Y(B_not[4]), .A(B[4]) );
  inv02 U65 ( .Y(n56), .A(n113) );
  inv02 U66 ( .Y(carry_3_), .A(n58) );
  inv02 U67 ( .Y(n59), .A(B_not[2]) );
  inv02 U68 ( .Y(n60), .A(A[2]) );
  inv02 U69 ( .Y(n61), .A(carry_2_) );
  nor02 U70 ( .Y(n62), .A0(n59), .A1(n63) );
  nor02 U71 ( .Y(n64), .A0(n60), .A1(n65) );
  nor02 U72 ( .Y(n66), .A0(n61), .A1(n67) );
  nor02 U73 ( .Y(n68), .A0(n61), .A1(n69) );
  nor02 U74 ( .Y(n57), .A0(n70), .A1(n71) );
  nor02 U75 ( .Y(n72), .A0(n60), .A1(n61) );
  nor02 U76 ( .Y(n73), .A0(n59), .A1(n61) );
  nor02 U77 ( .Y(n74), .A0(n59), .A1(n60) );
  nor02 U78 ( .Y(n58), .A0(n74), .A1(n75) );
  nor02 U79 ( .Y(n76), .A0(A[2]), .A1(carry_2_) );
  inv01 U80 ( .Y(n63), .A(n76) );
  nor02 U81 ( .Y(n77), .A0(B_not[2]), .A1(carry_2_) );
  inv01 U82 ( .Y(n65), .A(n77) );
  nor02 U83 ( .Y(n78), .A0(B_not[2]), .A1(A[2]) );
  inv01 U84 ( .Y(n67), .A(n78) );
  nor02 U85 ( .Y(n79), .A0(n59), .A1(n60) );
  inv01 U86 ( .Y(n69), .A(n79) );
  nor02 U87 ( .Y(n80), .A0(n62), .A1(n64) );
  inv01 U88 ( .Y(n70), .A(n80) );
  nor02 U89 ( .Y(n81), .A0(n66), .A1(n68) );
  inv01 U90 ( .Y(n71), .A(n81) );
  nor02 U91 ( .Y(n82), .A0(n72), .A1(n73) );
  inv01 U92 ( .Y(n75), .A(n82) );
  inv02 U93 ( .Y(DIFF[3]), .A(n83) );
  inv02 U94 ( .Y(carry_4_), .A(n84) );
  inv02 U95 ( .Y(n85), .A(B_not[3]) );
  inv02 U96 ( .Y(n86), .A(A[3]) );
  inv02 U97 ( .Y(n87), .A(carry_3_) );
  nor02 U98 ( .Y(n88), .A0(n85), .A1(n89) );
  nor02 U99 ( .Y(n90), .A0(n86), .A1(n91) );
  nor02 U100 ( .Y(n92), .A0(n87), .A1(n93) );
  nor02 U101 ( .Y(n94), .A0(n87), .A1(n95) );
  nor02 U102 ( .Y(n83), .A0(n96), .A1(n97) );
  nor02 U103 ( .Y(n98), .A0(n86), .A1(n87) );
  nor02 U104 ( .Y(n99), .A0(n85), .A1(n87) );
  nor02 U105 ( .Y(n100), .A0(n85), .A1(n86) );
  nor02 U106 ( .Y(n84), .A0(n100), .A1(n101) );
  nor02 U107 ( .Y(n102), .A0(A[3]), .A1(carry_3_) );
  inv01 U108 ( .Y(n89), .A(n102) );
  nor02 U109 ( .Y(n103), .A0(B_not[3]), .A1(carry_3_) );
  inv01 U110 ( .Y(n91), .A(n103) );
  nor02 U111 ( .Y(n104), .A0(B_not[3]), .A1(A[3]) );
  inv01 U112 ( .Y(n93), .A(n104) );
  nor02 U113 ( .Y(n105), .A0(n85), .A1(n86) );
  inv01 U114 ( .Y(n95), .A(n105) );
  nor02 U115 ( .Y(n106), .A0(n88), .A1(n90) );
  inv02 U116 ( .Y(n96), .A(n106) );
  nor02 U117 ( .Y(n107), .A0(n92), .A1(n94) );
  inv01 U118 ( .Y(n97), .A(n107) );
  nor02 U119 ( .Y(n108), .A0(n98), .A1(n99) );
  inv01 U120 ( .Y(n101), .A(n108) );
  inv02 U121 ( .Y(DIFF[1]), .A(n109) );
  inv02 U122 ( .Y(carry_2_), .A(n110) );
  inv02 U123 ( .Y(n111), .A(B_not[1]) );
  inv02 U124 ( .Y(n112), .A(A[1]) );
  inv02 U125 ( .Y(n113), .A(carry_1_) );
  nor02 U126 ( .Y(n114), .A0(n111), .A1(n115) );
  nor02 U127 ( .Y(n116), .A0(n112), .A1(n117) );
  nor02 U128 ( .Y(n118), .A0(n113), .A1(n119) );
  nor02 U129 ( .Y(n120), .A0(n113), .A1(n121) );
  nor02 U130 ( .Y(n109), .A0(n122), .A1(n123) );
  nor02 U131 ( .Y(n124), .A0(n112), .A1(n113) );
  nor02 U132 ( .Y(n125), .A0(n111), .A1(n113) );
  nor02 U133 ( .Y(n126), .A0(n111), .A1(n112) );
  nor02 U134 ( .Y(n110), .A0(n126), .A1(n127) );
  nor02 U135 ( .Y(n128), .A0(A[1]), .A1(carry_1_) );
  inv02 U136 ( .Y(n115), .A(n128) );
  nor02 U137 ( .Y(n129), .A0(B_not[1]), .A1(n56) );
  inv01 U138 ( .Y(n117), .A(n129) );
  nor02 U139 ( .Y(n130), .A0(B_not[1]), .A1(A[1]) );
  inv01 U140 ( .Y(n119), .A(n130) );
  nor02 U141 ( .Y(n131), .A0(n111), .A1(n112) );
  inv01 U142 ( .Y(n121), .A(n131) );
  nor02 U143 ( .Y(n132), .A0(n114), .A1(n116) );
  inv02 U144 ( .Y(n122), .A(n132) );
  nor02 U145 ( .Y(n133), .A0(n118), .A1(n120) );
  inv01 U146 ( .Y(n123), .A(n133) );
  nor02 U147 ( .Y(n134), .A0(n124), .A1(n125) );
  inv01 U148 ( .Y(n127), .A(n134) );
  inv02 U149 ( .Y(B_not[0]), .A(B[0]) );
  inv02 U150 ( .Y(B_not[2]), .A(B[2]) );
  inv02 U151 ( .Y(B_not[3]), .A(B[3]) );
  inv02 U152 ( .Y(B_not[1]), .A(B[1]) );
  xor2 U153 ( .Y(DIFF[6]), .A0(B_not[6]), .A1(carry_6_) );
  or02 U154 ( .Y(carry_1_), .A0(B_not[0]), .A1(A[0]) );
  xnor2 U155 ( .Y(n135), .A0(B_not[0]), .A1(A[0]) );
endmodule


module post_norm_mul_DW01_sub_10_0 ( A, B, CI, DIFF, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] DIFF;
  input CI;
  output CO;
  wire   carry_8_, carry_6_, carry_5_, carry_4_, carry_3_, carry_2_, B_not_5_,
         B_not_4_, B_not_3_, B_not_2_, B_not_1_, B_not_0_, n5, n6, n7, n9, n11,
         n12, n13, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99;

  nor02 U6 ( .Y(n5), .A0(A[8]), .A1(n18) );
  inv02 U7 ( .Y(n6), .A(n5) );
  xor2 U8 ( .Y(n7), .A0(B_not_0_), .A1(A[0]) );
  inv01 U9 ( .Y(DIFF[0]), .A(n7) );
  xor2 U10 ( .Y(n9), .A0(A[6]), .A1(n98) );
  inv01 U11 ( .Y(DIFF[6]), .A(n9) );
  nor02 U12 ( .Y(n11), .A0(B_not_0_), .A1(A[0]) );
  inv02 U13 ( .Y(n12), .A(n11) );
  xor2 U14 ( .Y(n13), .A0(A[7]), .A1(n16) );
  inv01 U15 ( .Y(DIFF[7]), .A(n13) );
  nor02 U16 ( .Y(n15), .A0(A[6]), .A1(n98) );
  inv02 U17 ( .Y(n16), .A(n15) );
  buf02 U18 ( .Y(n17), .A(carry_8_) );
  buf02 U19 ( .Y(n18), .A(carry_8_) );
  inv01 U20 ( .Y(DIFF[4]), .A(n19) );
  inv02 U21 ( .Y(carry_5_), .A(n20) );
  inv02 U22 ( .Y(n21), .A(B_not_4_) );
  inv02 U23 ( .Y(n22), .A(A[4]) );
  inv02 U24 ( .Y(n23), .A(carry_4_) );
  nor02 U25 ( .Y(n24), .A0(n21), .A1(n25) );
  nor02 U26 ( .Y(n26), .A0(n22), .A1(n27) );
  nor02 U27 ( .Y(n28), .A0(n23), .A1(n29) );
  nor02 U28 ( .Y(n30), .A0(n23), .A1(n31) );
  nor02 U29 ( .Y(n19), .A0(n32), .A1(n33) );
  nor02 U30 ( .Y(n34), .A0(n22), .A1(n23) );
  nor02 U31 ( .Y(n35), .A0(n21), .A1(n23) );
  nor02 U32 ( .Y(n36), .A0(n21), .A1(n22) );
  nor02 U33 ( .Y(n20), .A0(n36), .A1(n37) );
  nor02 U34 ( .Y(n38), .A0(A[4]), .A1(carry_4_) );
  inv01 U35 ( .Y(n25), .A(n38) );
  nor02 U36 ( .Y(n39), .A0(B_not_4_), .A1(carry_4_) );
  inv01 U37 ( .Y(n27), .A(n39) );
  nor02 U38 ( .Y(n40), .A0(B_not_4_), .A1(A[4]) );
  inv01 U39 ( .Y(n29), .A(n40) );
  nor02 U40 ( .Y(n41), .A0(n21), .A1(n22) );
  inv01 U41 ( .Y(n31), .A(n41) );
  nor02 U42 ( .Y(n42), .A0(n24), .A1(n26) );
  inv01 U43 ( .Y(n32), .A(n42) );
  nor02 U44 ( .Y(n43), .A0(n28), .A1(n30) );
  inv01 U45 ( .Y(n33), .A(n43) );
  nor02 U46 ( .Y(n44), .A0(n34), .A1(n35) );
  inv01 U47 ( .Y(n37), .A(n44) );
  inv02 U48 ( .Y(B_not_4_), .A(B[4]) );
  inv01 U49 ( .Y(DIFF[3]), .A(n45) );
  inv02 U50 ( .Y(carry_4_), .A(n46) );
  inv02 U51 ( .Y(n47), .A(B_not_3_) );
  inv02 U52 ( .Y(n48), .A(A[3]) );
  inv02 U53 ( .Y(n49), .A(carry_3_) );
  nor02 U54 ( .Y(n50), .A0(n47), .A1(n51) );
  nor02 U55 ( .Y(n52), .A0(n48), .A1(n53) );
  nor02 U56 ( .Y(n54), .A0(n49), .A1(n55) );
  nor02 U57 ( .Y(n56), .A0(n49), .A1(n57) );
  nor02 U58 ( .Y(n45), .A0(n58), .A1(n59) );
  nor02 U59 ( .Y(n60), .A0(n48), .A1(n49) );
  nor02 U60 ( .Y(n61), .A0(n47), .A1(n49) );
  nor02 U61 ( .Y(n62), .A0(n47), .A1(n48) );
  nor02 U62 ( .Y(n46), .A0(n62), .A1(n63) );
  nor02 U63 ( .Y(n64), .A0(A[3]), .A1(carry_3_) );
  inv01 U64 ( .Y(n51), .A(n64) );
  nor02 U65 ( .Y(n65), .A0(B_not_3_), .A1(carry_3_) );
  inv01 U66 ( .Y(n53), .A(n65) );
  nor02 U67 ( .Y(n66), .A0(B_not_3_), .A1(A[3]) );
  inv01 U68 ( .Y(n55), .A(n66) );
  nor02 U69 ( .Y(n67), .A0(n47), .A1(n48) );
  inv01 U70 ( .Y(n57), .A(n67) );
  nor02 U71 ( .Y(n68), .A0(n50), .A1(n52) );
  inv01 U72 ( .Y(n58), .A(n68) );
  nor02 U73 ( .Y(n69), .A0(n54), .A1(n56) );
  inv01 U74 ( .Y(n59), .A(n69) );
  nor02 U75 ( .Y(n70), .A0(n60), .A1(n61) );
  inv01 U76 ( .Y(n63), .A(n70) );
  inv02 U77 ( .Y(B_not_3_), .A(B[3]) );
  inv01 U78 ( .Y(DIFF[2]), .A(n71) );
  inv02 U79 ( .Y(carry_3_), .A(n72) );
  inv02 U80 ( .Y(n73), .A(B_not_2_) );
  inv02 U81 ( .Y(n74), .A(A[2]) );
  inv02 U82 ( .Y(n75), .A(n97) );
  nor02 U83 ( .Y(n76), .A0(n73), .A1(n77) );
  nor02 U84 ( .Y(n78), .A0(n74), .A1(n79) );
  nor02 U85 ( .Y(n80), .A0(n75), .A1(n81) );
  nor02 U86 ( .Y(n82), .A0(n75), .A1(n83) );
  nor02 U87 ( .Y(n71), .A0(n84), .A1(n85) );
  nor02 U88 ( .Y(n86), .A0(n74), .A1(n75) );
  nor02 U89 ( .Y(n87), .A0(n73), .A1(n75) );
  nor02 U90 ( .Y(n88), .A0(n73), .A1(n74) );
  nor02 U91 ( .Y(n72), .A0(n88), .A1(n89) );
  nor02 U92 ( .Y(n90), .A0(A[2]), .A1(n97) );
  inv01 U93 ( .Y(n77), .A(n90) );
  nor02 U94 ( .Y(n91), .A0(B_not_2_), .A1(n97) );
  inv01 U95 ( .Y(n79), .A(n91) );
  nor02 U96 ( .Y(n92), .A0(B_not_2_), .A1(A[2]) );
  inv01 U97 ( .Y(n81), .A(n92) );
  nor02 U98 ( .Y(n93), .A0(n73), .A1(n74) );
  inv01 U99 ( .Y(n83), .A(n93) );
  nor02 U100 ( .Y(n94), .A0(n76), .A1(n78) );
  inv01 U101 ( .Y(n84), .A(n94) );
  nor02 U102 ( .Y(n95), .A0(n80), .A1(n82) );
  inv01 U103 ( .Y(n85), .A(n95) );
  nor02 U104 ( .Y(n96), .A0(n86), .A1(n87) );
  inv01 U105 ( .Y(n89), .A(n96) );
  inv02 U106 ( .Y(B_not_2_), .A(B[2]) );
  buf02 U107 ( .Y(n97), .A(carry_2_) );
  buf02 U108 ( .Y(n98), .A(carry_6_) );
  xor2 U109 ( .Y(n99), .A0(A[8]), .A1(n17) );
  inv02 U110 ( .Y(DIFF[8]), .A(n99) );
  xnor2 U111 ( .Y(DIFF[9]), .A0(A[9]), .A1(n6) );
  or02 U112 ( .Y(carry_8_), .A0(A[7]), .A1(n16) );
  inv04 U113 ( .Y(B_not_5_), .A(B[5]) );
  inv04 U114 ( .Y(B_not_1_), .A(B[1]) );
  inv04 U115 ( .Y(B_not_0_), .A(B[0]) );
  fadd1 U2_1 ( .S(DIFF[1]), .CO(carry_2_), .A(A[1]), .B(B_not_1_), .CI(n12) );
  fadd1 U2_5 ( .S(DIFF[5]), .CO(carry_6_), .A(A[5]), .B(B_not_5_), .CI(
        carry_5_) );
endmodule


module post_norm_mul_DW01_cmp2_6_0 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [5:0] A;
  input [5:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42;

  buf02 U6 ( .Y(n15), .A(n29) );
  inv02 U7 ( .Y(n30), .A(B[5]) );
  inv01 U8 ( .Y(n42), .A(B[0]) );
  inv01 U9 ( .Y(n31), .A(n16) );
  nor02 U10 ( .Y(n17), .A0(B[4]), .A1(n33) );
  nor02 U11 ( .Y(n18), .A0(B[3]), .A1(n34) );
  inv01 U12 ( .Y(n19), .A(n35) );
  nor02 U13 ( .Y(n16), .A0(n19), .A1(n20) );
  nor02 U14 ( .Y(n21), .A0(n17), .A1(n18) );
  inv01 U15 ( .Y(n20), .A(n21) );
  inv02 U16 ( .Y(n34), .A(A[3]) );
  inv02 U17 ( .Y(n33), .A(A[4]) );
  inv01 U18 ( .Y(n38), .A(n22) );
  nor02 U19 ( .Y(n23), .A0(B[2]), .A1(n36) );
  nor02 U20 ( .Y(n24), .A0(n39), .A1(n40) );
  inv01 U21 ( .Y(n25), .A(n41) );
  nor02 U22 ( .Y(n22), .A0(n25), .A1(n26) );
  nor02 U23 ( .Y(n27), .A0(n23), .A1(n24) );
  inv01 U24 ( .Y(n26), .A(n27) );
  inv01 U25 ( .Y(n37), .A(n38) );
  inv02 U26 ( .Y(n40), .A(A[1]) );
  inv02 U27 ( .Y(n36), .A(A[2]) );
  inv04 U28 ( .Y(n28), .A(A[5]) );
  ao21 U29 ( .Y(LT_LE), .A0(B[5]), .A1(n28), .B0(n15) );
  aoi22 U30 ( .Y(n29), .A0(A[5]), .A1(n30), .B0(n31), .B1(n32) );
  nand02 U31 ( .Y(n32), .A0(B[4]), .A1(n33) );
  ao221 U32 ( .Y(n35), .A0(n36), .A1(B[2]), .B0(n34), .B1(B[3]), .C0(n37) );
  ao21 U33 ( .Y(n41), .A0(n39), .A1(n40), .B0(B[1]) );
  nor02 U34 ( .Y(n39), .A0(n42), .A1(A[0]) );
endmodule


module post_norm_mul ( clk_i, opa_i, opb_i, exp_10_i, fract_48_i, sign_i, 
        rmode_i, output_o, ine_o );
  input [31:0] opa_i;
  input [31:0] opb_i;
  input [9:0] exp_10_i;
  input [47:0] fract_48_i;
  input [1:0] rmode_i;
  output [31:0] output_o;
  input clk_i, sign_i;
  output ine_o;
  wire   s_output_o_30_, s_output_o_29_, s_output_o_28_, s_output_o_27_,
         s_output_o_26_, s_output_o_25_, s_output_o_24_, s_output_o_23_,
         s_output_o_22_, s_output_o_21_, s_output_o_20_, s_output_o_19_,
         s_output_o_18_, s_output_o_17_, s_output_o_16_, s_output_o_15_,
         s_output_o_14_, s_output_o_13_, s_output_o_12_, s_output_o_11_,
         s_output_o_10_, s_output_o_9_, s_output_o_8_, s_output_o_7_,
         s_output_o_6_, s_output_o_5_, s_output_o_4_, s_output_o_3_,
         s_output_o_2_, s_output_o_1_, s_output_o_0_, v_shl15711_5_,
         v_shl15711_4_, v_shl15711_3_, v_shl15711_2_, v_shl15711_1_,
         v_shl15711_0_, s_frac2a_47_, s_frac2a_46_, s_frac2a_45_, s_frac2a_44_,
         s_frac2a_43_, s_frac2a_42_, s_frac2a_41_, s_frac2a_40_, s_frac2a_39_,
         s_frac2a_38_, s_frac2a_37_, s_frac2a_36_, s_frac2a_35_, s_frac2a_34_,
         s_frac2a_33_, s_frac2a_32_, s_frac2a_31_, s_frac2a_30_, s_frac2a_29_,
         s_frac2a_28_, s_frac2a_27_, s_frac2a_26_, s_frac2a_25_, s_frac2a_24_,
         s_frac2a_23_, s_frac2a_20_, s_frac2a_19_, s_frac2a_15_, s_frac2a_14_,
         s_frac2a_13_, s_frac2a_10_, s_frac2a_6_, s_frac2a_5_, s_frac2a_4_,
         s_frac2a_1_, s_frac2a_0_, s_round, s_sign_i, s_frac_rnd_23_,
         s_frac_rnd_22_, s_frac_rnd_1_, s_shr3, s_opa_i_30_, s_opa_i_29_,
         s_opa_i_28_, s_opa_i_25_, s_opa_i_24_, s_opa_i_23_, s_opa_i_21_,
         s_opa_i_20_, s_opa_i_16_, s_opa_i_15_, s_opa_i_14_, s_opa_i_11_,
         s_opa_i_10_, s_opa_i_6_, s_opa_i_5_, s_opa_i_4_, s_opa_i_1_,
         s_opa_i_0_, s_opb_i_30_, s_opb_i_29_, s_opb_i_28_, s_opb_i_25_,
         s_opb_i_24_, s_opb_i_23_, s_opb_i_21_, s_opb_i_20_, s_opb_i_16_,
         s_opb_i_15_, s_opb_i_14_, s_opb_i_11_, s_opb_i_10_, s_opb_i_6_,
         s_opb_i_5_, s_opb_i_4_, s_opb_i_1_, s_opb_i_0_, s_exp_10_i_8_,
         s_exp_10_i_7_, s_exp_10_i_6_, s_exp_10_i_5_, s_exp_10_i_4_,
         s_exp_10_i_3_, s_exp_10_i_2_, s_exp_10_i_1_, s_exp_10_i_0_,
         s_rmode_i_1_, s_rmode_i_0_, s_zeros1047_0_, v_count3287_5_,
         v_count3287_4_, v_count3287_3_, v_count3287_2_, v_count3287_1_,
         v_count3287_0_, s_r_zeros_5_, s_r_zeros_4_, s_r_zeros_3_,
         s_r_zeros_2_, s_r_zeros_1_, s_r_zeros_0_, s_exp_10a_9_, s_exp_10a_8_,
         s_exp_10a_7_, s_exp_10a_6_, s_exp_10a_4_, s_expo15773_7_,
         s_expo15773_6_, s_expo15773_5_, s_expo15773_4_, s_expo15773_3_,
         s_expo15773_2_, s_expo15773_1_, s_expo15773_0_, s_shr25775_5_,
         s_shr25775_4_, s_shr25775_3_, s_shr25775_2_, s_shr25775_1_,
         s_shr25775_0_, s_shr2_5_, s_shr2_4_, s_shr2_3_, s_shr2_2_, s_shr2_1_,
         s_shr2_0_, s_shl2_5_, s_shl2_4_, s_shl2_3_, s_shl2_2_, s_shl2_1_,
         s_shl2_0_, n____return5956_5_, n____return5956_4_, n____return5956_3_,
         n____return5956_2_, n____return5956_1_, n____return5956_0_,
         n____return6004_6_, s_frac2a6207_47_, s_frac2a6207_46_,
         s_frac2a6207_45_, s_frac2a6207_44_, s_frac2a6207_43_,
         s_frac2a6207_42_, s_frac2a6207_41_, s_frac2a6207_40_,
         s_frac2a6207_39_, s_frac2a6207_38_, s_frac2a6207_37_,
         s_frac2a6207_36_, s_frac2a6207_35_, s_frac2a6207_34_,
         s_frac2a6207_33_, s_frac2a6207_32_, s_frac2a6207_31_,
         s_frac2a6207_30_, s_frac2a6207_29_, s_frac2a6207_28_,
         s_frac2a6207_27_, s_frac2a6207_26_, s_frac2a6207_25_,
         s_frac2a6207_24_, s_frac2a6207_23_, s_frac2a6207_22_,
         s_frac2a6207_21_, s_frac2a6207_20_, s_frac2a6207_19_,
         s_frac2a6207_18_, s_frac2a6207_17_, s_frac2a6207_16_,
         s_frac2a6207_15_, s_frac2a6207_14_, s_frac2a6207_13_,
         s_frac2a6207_12_, s_frac2a6207_11_, s_frac2a6207_10_, s_frac2a6207_9_,
         s_frac2a6207_8_, s_frac2a6207_7_, s_frac2a6207_6_, s_frac2a6207_5_,
         s_frac2a6207_4_, s_frac2a6207_3_, s_frac2a6207_2_, s_frac2a6207_1_,
         s_frac2a6207_0_, n6653_8_, n____return6651_7_, n____return6651_6_,
         n____return6651_5_, n____return6651_4_, n____return6651_3_,
         n____return6651_2_, n____return6651_1_, n____return6651_0_,
         n____return6760, n____return6722_5_, n____return6722_3_,
         n____return6722_1_, s_frac_rnd7043_24_, s_frac_rnd7043_23_,
         s_frac_rnd7043_22_, s_frac_rnd7043_21_, s_frac_rnd7043_20_,
         s_frac_rnd7043_19_, s_frac_rnd7043_18_, s_frac_rnd7043_17_,
         s_frac_rnd7043_16_, s_frac_rnd7043_15_, s_frac_rnd7043_14_,
         s_frac_rnd7043_13_, s_frac_rnd7043_12_, s_frac_rnd7043_11_,
         s_frac_rnd7043_10_, s_frac_rnd7043_9_, s_frac_rnd7043_8_,
         s_frac_rnd7043_7_, s_frac_rnd7043_6_, s_frac_rnd7043_5_,
         s_frac_rnd7043_4_, s_frac_rnd7043_3_, s_frac_rnd7043_2_,
         s_frac_rnd7043_1_, s_frac_rnd7043_0_, n7072_23_, n____return7070_24_,
         n____return7070_22_, n____return7070_21_, n____return7070_20_,
         n____return7070_19_, n____return7070_18_, n____return7070_17_,
         n____return7070_16_, n____return7070_15_, n____return7070_14_,
         n____return7070_13_, n____return7070_12_, n____return7070_11_,
         n____return7070_10_, n____return7070_9_, n____return7070_8_,
         n____return7070_7_, n____return7070_6_, n____return7070_5_,
         n____return7070_4_, n____return7070_3_, n____return7070_2_,
         n____return7070_1_, n____return7070_0_, n7170_8_, n____return7168_7_,
         n____return7168_6_, n____return7168_5_, n____return7168_4_,
         n____return7168_3_, n____return7168_2_, n____return7168_1_,
         n____return7168_0_, U1086_U4_Z_6, U1086_U3_Z_0, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500;
  wire   [47:0] s_fract_48_i;
  wire   [5:0] s_zeros;
  wire   [9:0] s_exp_10b;
  wire   [8:0] s_expo1;
  wire   [8:0] s_expo2b;

  dff s_expo1_reg_8_ ( .Q(s_expo1[8]), .D(1'b0), .CLK(clk_i) );
  dff s_expa_reg_7_ ( .QB(n14460), .D(opa_i[30]), .CLK(clk_i) );
  dff s_expa_reg_6_ ( .QB(n14459), .D(opa_i[29]), .CLK(clk_i) );
  dff s_expa_reg_5_ ( .QB(n14458), .D(opa_i[28]), .CLK(clk_i) );
  dff s_expa_reg_4_ ( .QB(n14457), .D(opa_i[27]), .CLK(clk_i) );
  dff s_expa_reg_3_ ( .QB(n14464), .D(opa_i[26]), .CLK(clk_i) );
  dff s_expa_reg_2_ ( .QB(n14463), .D(opa_i[25]), .CLK(clk_i) );
  dff s_expa_reg_1_ ( .QB(n14462), .D(opa_i[24]), .CLK(clk_i) );
  dff s_expa_reg_0_ ( .QB(n14461), .D(opa_i[23]), .CLK(clk_i) );
  dff s_expb_reg_7_ ( .QB(n14452), .D(opb_i[30]), .CLK(clk_i) );
  dff s_expb_reg_6_ ( .QB(n14451), .D(opb_i[29]), .CLK(clk_i) );
  dff s_expb_reg_5_ ( .QB(n14450), .D(opb_i[28]), .CLK(clk_i) );
  dff s_expb_reg_4_ ( .QB(n14449), .D(opb_i[27]), .CLK(clk_i) );
  dff s_expb_reg_3_ ( .QB(n14456), .D(opb_i[26]), .CLK(clk_i) );
  dff s_expb_reg_2_ ( .QB(n14455), .D(opb_i[25]), .CLK(clk_i) );
  dff s_expb_reg_1_ ( .QB(n14454), .D(opb_i[24]), .CLK(clk_i) );
  dff s_expb_reg_0_ ( .QB(n14453), .D(opb_i[23]), .CLK(clk_i) );
  dff s_exp_10_i_reg_9_ ( .QB(n14500), .D(exp_10_i[9]), .CLK(clk_i) );
  dff s_exp_10_i_reg_8_ ( .Q(s_exp_10_i_8_), .D(exp_10_i[8]), .CLK(clk_i) );
  dff s_exp_10_i_reg_7_ ( .Q(s_exp_10_i_7_), .D(exp_10_i[7]), .CLK(clk_i) );
  dff s_exp_10_i_reg_6_ ( .Q(s_exp_10_i_6_), .D(exp_10_i[6]), .CLK(clk_i) );
  dff s_exp_10_i_reg_5_ ( .Q(s_exp_10_i_5_), .D(exp_10_i[5]), .CLK(clk_i) );
  dff s_exp_10_i_reg_4_ ( .Q(s_exp_10_i_4_), .D(exp_10_i[4]), .CLK(clk_i) );
  dff s_exp_10_i_reg_3_ ( .Q(s_exp_10_i_3_), .D(exp_10_i[3]), .CLK(clk_i) );
  dff s_exp_10_i_reg_2_ ( .Q(s_exp_10_i_2_), .D(exp_10_i[2]), .CLK(clk_i) );
  dff s_exp_10_i_reg_1_ ( .Q(s_exp_10_i_1_), .D(exp_10_i[1]), .CLK(clk_i) );
  dff s_exp_10_i_reg_0_ ( .Q(s_exp_10_i_0_), .D(exp_10_i[0]), .CLK(clk_i) );
  dff s_fract_48_i_reg_47_ ( .Q(s_fract_48_i[47]), .D(fract_48_i[47]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_46_ ( .Q(s_fract_48_i[46]), .D(fract_48_i[46]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_45_ ( .Q(s_fract_48_i[45]), .D(fract_48_i[45]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_44_ ( .Q(s_fract_48_i[44]), .D(fract_48_i[44]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_43_ ( .Q(s_fract_48_i[43]), .D(fract_48_i[43]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_42_ ( .Q(s_fract_48_i[42]), .D(fract_48_i[42]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_41_ ( .Q(s_fract_48_i[41]), .D(fract_48_i[41]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_40_ ( .Q(s_fract_48_i[40]), .D(fract_48_i[40]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_39_ ( .Q(s_fract_48_i[39]), .D(fract_48_i[39]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_38_ ( .Q(s_fract_48_i[38]), .D(fract_48_i[38]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_37_ ( .Q(s_fract_48_i[37]), .D(fract_48_i[37]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_36_ ( .Q(s_fract_48_i[36]), .D(fract_48_i[36]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_35_ ( .Q(s_fract_48_i[35]), .D(fract_48_i[35]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_34_ ( .Q(s_fract_48_i[34]), .D(fract_48_i[34]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_33_ ( .Q(s_fract_48_i[33]), .D(fract_48_i[33]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_32_ ( .Q(s_fract_48_i[32]), .D(fract_48_i[32]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_31_ ( .Q(s_fract_48_i[31]), .D(fract_48_i[31]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_30_ ( .Q(s_fract_48_i[30]), .D(fract_48_i[30]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_29_ ( .Q(s_fract_48_i[29]), .D(fract_48_i[29]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_28_ ( .Q(s_fract_48_i[28]), .D(fract_48_i[28]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_27_ ( .Q(s_fract_48_i[27]), .D(fract_48_i[27]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_26_ ( .Q(s_fract_48_i[26]), .D(fract_48_i[26]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_25_ ( .Q(s_fract_48_i[25]), .D(fract_48_i[25]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_24_ ( .Q(s_fract_48_i[24]), .D(fract_48_i[24]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_23_ ( .Q(s_fract_48_i[23]), .D(fract_48_i[23]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_22_ ( .Q(s_fract_48_i[22]), .D(fract_48_i[22]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_21_ ( .Q(s_fract_48_i[21]), .D(fract_48_i[21]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_20_ ( .Q(s_fract_48_i[20]), .D(fract_48_i[20]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_19_ ( .Q(s_fract_48_i[19]), .D(fract_48_i[19]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_18_ ( .Q(s_fract_48_i[18]), .D(fract_48_i[18]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_17_ ( .Q(s_fract_48_i[17]), .D(fract_48_i[17]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_16_ ( .Q(s_fract_48_i[16]), .D(fract_48_i[16]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_15_ ( .Q(s_fract_48_i[15]), .D(fract_48_i[15]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_14_ ( .Q(s_fract_48_i[14]), .D(fract_48_i[14]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_13_ ( .Q(s_fract_48_i[13]), .D(fract_48_i[13]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_12_ ( .Q(s_fract_48_i[12]), .D(fract_48_i[12]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_11_ ( .Q(s_fract_48_i[11]), .D(fract_48_i[11]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_10_ ( .Q(s_fract_48_i[10]), .D(fract_48_i[10]), .CLK(
        clk_i) );
  dff s_fract_48_i_reg_9_ ( .Q(s_fract_48_i[9]), .D(fract_48_i[9]), .CLK(clk_i) );
  dff s_fract_48_i_reg_8_ ( .Q(s_fract_48_i[8]), .D(fract_48_i[8]), .CLK(clk_i) );
  dff s_fract_48_i_reg_7_ ( .Q(s_fract_48_i[7]), .D(fract_48_i[7]), .CLK(clk_i) );
  dff s_fract_48_i_reg_6_ ( .Q(s_fract_48_i[6]), .D(fract_48_i[6]), .CLK(clk_i) );
  dff s_fract_48_i_reg_5_ ( .Q(s_fract_48_i[5]), .D(fract_48_i[5]), .CLK(clk_i) );
  dff s_fract_48_i_reg_4_ ( .Q(s_fract_48_i[4]), .D(fract_48_i[4]), .CLK(clk_i) );
  dff s_fract_48_i_reg_3_ ( .Q(s_fract_48_i[3]), .D(fract_48_i[3]), .CLK(clk_i) );
  dff s_fract_48_i_reg_2_ ( .Q(s_fract_48_i[2]), .D(fract_48_i[2]), .CLK(clk_i) );
  dff s_fract_48_i_reg_1_ ( .Q(s_fract_48_i[1]), .D(fract_48_i[1]), .CLK(clk_i) );
  dff s_fract_48_i_reg_0_ ( .Q(s_fract_48_i[0]), .D(fract_48_i[0]), .CLK(clk_i) );
  dff s_rmode_i_reg_1_ ( .Q(s_rmode_i_1_), .D(rmode_i[1]), .CLK(clk_i) );
  dff s_rmode_i_reg_0_ ( .Q(s_rmode_i_0_), .D(rmode_i[0]), .CLK(clk_i) );
  dff output_o_reg_31_ ( .Q(output_o[31]), .D(s_sign_i), .CLK(clk_i) );
  dff output_o_reg_30_ ( .Q(output_o[30]), .D(s_output_o_30_), .CLK(clk_i) );
  dff output_o_reg_29_ ( .Q(output_o[29]), .D(s_output_o_29_), .CLK(clk_i) );
  dff output_o_reg_28_ ( .Q(output_o[28]), .D(s_output_o_28_), .CLK(clk_i) );
  dff output_o_reg_27_ ( .Q(output_o[27]), .D(s_output_o_27_), .CLK(clk_i) );
  dff output_o_reg_26_ ( .Q(output_o[26]), .D(s_output_o_26_), .CLK(clk_i) );
  dff output_o_reg_25_ ( .Q(output_o[25]), .D(s_output_o_25_), .CLK(clk_i) );
  dff output_o_reg_24_ ( .Q(output_o[24]), .D(s_output_o_24_), .CLK(clk_i) );
  dff output_o_reg_23_ ( .Q(output_o[23]), .D(s_output_o_23_), .CLK(clk_i) );
  dff output_o_reg_22_ ( .Q(output_o[22]), .D(s_output_o_22_), .CLK(clk_i) );
  dff output_o_reg_21_ ( .Q(output_o[21]), .D(s_output_o_21_), .CLK(clk_i) );
  dff output_o_reg_20_ ( .Q(output_o[20]), .D(s_output_o_20_), .CLK(clk_i) );
  dff output_o_reg_19_ ( .Q(output_o[19]), .D(s_output_o_19_), .CLK(clk_i) );
  dff output_o_reg_18_ ( .Q(output_o[18]), .D(s_output_o_18_), .CLK(clk_i) );
  dff output_o_reg_17_ ( .Q(output_o[17]), .D(s_output_o_17_), .CLK(clk_i) );
  dff output_o_reg_16_ ( .Q(output_o[16]), .D(s_output_o_16_), .CLK(clk_i) );
  dff output_o_reg_15_ ( .Q(output_o[15]), .D(s_output_o_15_), .CLK(clk_i) );
  dff output_o_reg_14_ ( .Q(output_o[14]), .D(s_output_o_14_), .CLK(clk_i) );
  dff output_o_reg_13_ ( .Q(output_o[13]), .D(s_output_o_13_), .CLK(clk_i) );
  dff output_o_reg_12_ ( .Q(output_o[12]), .D(s_output_o_12_), .CLK(clk_i) );
  dff output_o_reg_11_ ( .Q(output_o[11]), .D(s_output_o_11_), .CLK(clk_i) );
  dff output_o_reg_10_ ( .Q(output_o[10]), .D(s_output_o_10_), .CLK(clk_i) );
  dff output_o_reg_9_ ( .Q(output_o[9]), .D(s_output_o_9_), .CLK(clk_i) );
  dff output_o_reg_8_ ( .Q(output_o[8]), .D(s_output_o_8_), .CLK(clk_i) );
  dff output_o_reg_7_ ( .Q(output_o[7]), .D(s_output_o_7_), .CLK(clk_i) );
  dff output_o_reg_6_ ( .Q(output_o[6]), .D(s_output_o_6_), .CLK(clk_i) );
  dff output_o_reg_5_ ( .Q(output_o[5]), .D(s_output_o_5_), .CLK(clk_i) );
  dff output_o_reg_4_ ( .Q(output_o[4]), .D(s_output_o_4_), .CLK(clk_i) );
  dff output_o_reg_3_ ( .Q(output_o[3]), .D(s_output_o_3_), .CLK(clk_i) );
  dff output_o_reg_2_ ( .Q(output_o[2]), .D(s_output_o_2_), .CLK(clk_i) );
  dff output_o_reg_1_ ( .Q(output_o[1]), .D(s_output_o_1_), .CLK(clk_i) );
  dff output_o_reg_0_ ( .Q(output_o[0]), .D(s_output_o_0_), .CLK(clk_i) );
  dff s_zeros_reg_5_ ( .Q(s_zeros[5]), .D(n9778), .CLK(clk_i) );
  dff s_zeros_reg_4_ ( .Q(s_zeros[4]), .D(n9900), .CLK(clk_i) );
  dff s_zeros_reg_3_ ( .Q(s_zeros[3]), .D(n9776), .CLK(clk_i) );
  dff s_zeros_reg_2_ ( .Q(s_zeros[2]), .D(n9762), .CLK(clk_i) );
  dff s_zeros_reg_1_ ( .Q(s_zeros[1]), .D(n9764), .CLK(clk_i) );
  dff s_zeros_reg_0_ ( .Q(s_zeros[0]), .D(s_zeros1047_0_), .CLK(clk_i) );
  dff s_r_zeros_reg_5_ ( .Q(s_r_zeros_5_), .QB(n14421), .D(v_count3287_5_), 
        .CLK(clk_i) );
  dff s_r_zeros_reg_4_ ( .Q(s_r_zeros_4_), .QB(n14422), .D(v_count3287_4_), 
        .CLK(clk_i) );
  dff s_r_zeros_reg_3_ ( .Q(s_r_zeros_3_), .D(v_count3287_3_), .CLK(clk_i) );
  dff s_r_zeros_reg_2_ ( .Q(s_r_zeros_2_), .D(v_count3287_2_), .CLK(clk_i) );
  dff s_r_zeros_reg_1_ ( .Q(s_r_zeros_1_), .D(v_count3287_1_), .CLK(clk_i) );
  dff s_r_zeros_reg_0_ ( .Q(s_r_zeros_0_), .D(n10198), .CLK(clk_i) );
  dff s_expo1_reg_7_ ( .Q(s_expo1[7]), .D(s_expo15773_7_), .CLK(clk_i) );
  dff s_expo1_reg_6_ ( .Q(s_expo1[6]), .D(s_expo15773_6_), .CLK(clk_i) );
  dff s_expo1_reg_5_ ( .Q(s_expo1[5]), .D(s_expo15773_5_), .CLK(clk_i) );
  dff s_expo1_reg_4_ ( .Q(s_expo1[4]), .D(s_expo15773_4_), .CLK(clk_i) );
  dff s_expo1_reg_3_ ( .Q(s_expo1[3]), .D(s_expo15773_3_), .CLK(clk_i) );
  dff s_expo1_reg_2_ ( .Q(s_expo1[2]), .D(s_expo15773_2_), .CLK(clk_i) );
  dff s_expo1_reg_1_ ( .Q(s_expo1[1]), .D(s_expo15773_1_), .CLK(clk_i) );
  dff s_expo1_reg_0_ ( .Q(s_expo1[0]), .D(s_expo15773_0_), .CLK(clk_i) );
  dff s_shr2_reg_5_ ( .Q(s_shr2_5_), .D(s_shr25775_5_), .CLK(clk_i) );
  dff s_shr2_reg_4_ ( .Q(s_shr2_4_), .D(s_shr25775_4_), .CLK(clk_i) );
  dff s_shr2_reg_3_ ( .Q(s_shr2_3_), .D(s_shr25775_3_), .CLK(clk_i) );
  dff s_shr2_reg_2_ ( .Q(s_shr2_2_), .D(s_shr25775_2_), .CLK(clk_i) );
  dff s_shr2_reg_1_ ( .Q(s_shr2_1_), .D(s_shr25775_1_), .CLK(clk_i) );
  dff s_shr2_reg_0_ ( .Q(s_shr2_0_), .QB(n10280), .D(s_shr25775_0_), .CLK(
        clk_i) );
  dff s_shl2_reg_5_ ( .Q(s_shl2_5_), .D(v_shl15711_5_), .CLK(clk_i) );
  dff s_shl2_reg_4_ ( .Q(s_shl2_4_), .D(v_shl15711_4_), .CLK(clk_i) );
  dff s_shl2_reg_3_ ( .Q(s_shl2_3_), .D(v_shl15711_3_), .CLK(clk_i) );
  dff s_shl2_reg_2_ ( .Q(s_shl2_2_), .D(v_shl15711_2_), .CLK(clk_i) );
  dff s_shl2_reg_1_ ( .Q(s_shl2_1_), .D(v_shl15711_1_), .CLK(clk_i) );
  dff s_shl2_reg_0_ ( .Q(s_shl2_0_), .D(v_shl15711_0_), .CLK(clk_i) );
  dff s_frac2a_reg_47_ ( .Q(s_frac2a_47_), .QB(n14473), .D(s_frac2a6207_47_), 
        .CLK(clk_i) );
  dff s_frac2a_reg_46_ ( .Q(s_frac2a_46_), .QB(n13519), .D(s_frac2a6207_46_), 
        .CLK(clk_i) );
  dff s_frac2a_reg_45_ ( .Q(s_frac2a_45_), .QB(n14474), .D(s_frac2a6207_45_), 
        .CLK(clk_i) );
  dff s_frac2a_reg_44_ ( .Q(s_frac2a_44_), .QB(n14475), .D(s_frac2a6207_44_), 
        .CLK(clk_i) );
  dff s_frac2a_reg_43_ ( .Q(s_frac2a_43_), .QB(n14476), .D(s_frac2a6207_43_), 
        .CLK(clk_i) );
  dff s_frac2a_reg_42_ ( .Q(s_frac2a_42_), .QB(n14478), .D(s_frac2a6207_42_), 
        .CLK(clk_i) );
  dff s_frac2a_reg_41_ ( .Q(s_frac2a_41_), .QB(n14479), .D(s_frac2a6207_41_), 
        .CLK(clk_i) );
  dff s_frac2a_reg_40_ ( .Q(s_frac2a_40_), .QB(n14480), .D(s_frac2a6207_40_), 
        .CLK(clk_i) );
  dff s_frac2a_reg_39_ ( .Q(s_frac2a_39_), .QB(n14481), .D(s_frac2a6207_39_), 
        .CLK(clk_i) );
  dff s_frac2a_reg_38_ ( .Q(s_frac2a_38_), .QB(n14482), .D(s_frac2a6207_38_), 
        .CLK(clk_i) );
  dff s_frac2a_reg_37_ ( .Q(s_frac2a_37_), .QB(n14483), .D(s_frac2a6207_37_), 
        .CLK(clk_i) );
  dff s_frac2a_reg_36_ ( .Q(s_frac2a_36_), .QB(n14484), .D(s_frac2a6207_36_), 
        .CLK(clk_i) );
  dff s_frac2a_reg_35_ ( .Q(s_frac2a_35_), .QB(n14485), .D(s_frac2a6207_35_), 
        .CLK(clk_i) );
  dff s_frac2a_reg_34_ ( .Q(s_frac2a_34_), .QB(n14486), .D(s_frac2a6207_34_), 
        .CLK(clk_i) );
  dff s_frac2a_reg_33_ ( .Q(s_frac2a_33_), .QB(n14487), .D(s_frac2a6207_33_), 
        .CLK(clk_i) );
  dff s_frac2a_reg_32_ ( .Q(s_frac2a_32_), .QB(n14465), .D(s_frac2a6207_32_), 
        .CLK(clk_i) );
  dff s_frac2a_reg_31_ ( .Q(s_frac2a_31_), .QB(n14466), .D(s_frac2a6207_31_), 
        .CLK(clk_i) );
  dff s_frac2a_reg_30_ ( .Q(s_frac2a_30_), .QB(n14467), .D(s_frac2a6207_30_), 
        .CLK(clk_i) );
  dff s_frac2a_reg_29_ ( .Q(s_frac2a_29_), .QB(n14468), .D(s_frac2a6207_29_), 
        .CLK(clk_i) );
  dff s_frac2a_reg_28_ ( .Q(s_frac2a_28_), .QB(n14469), .D(s_frac2a6207_28_), 
        .CLK(clk_i) );
  dff s_frac2a_reg_27_ ( .Q(s_frac2a_27_), .QB(n14470), .D(s_frac2a6207_27_), 
        .CLK(clk_i) );
  dff s_frac2a_reg_26_ ( .Q(s_frac2a_26_), .QB(n14471), .D(s_frac2a6207_26_), 
        .CLK(clk_i) );
  dff s_frac2a_reg_25_ ( .Q(s_frac2a_25_), .QB(n14472), .D(s_frac2a6207_25_), 
        .CLK(clk_i) );
  dff s_frac2a_reg_24_ ( .Q(s_frac2a_24_), .QB(n14477), .D(s_frac2a6207_24_), 
        .CLK(clk_i) );
  dff s_frac2a_reg_23_ ( .Q(s_frac2a_23_), .D(s_frac2a6207_23_), .CLK(clk_i)
         );
  dff s_frac2a_reg_22_ ( .Q(n14489), .D(s_frac2a6207_22_), .CLK(clk_i) );
  dff s_frac2a_reg_21_ ( .Q(s_round), .D(s_frac2a6207_21_), .CLK(clk_i) );
  dff s_frac2a_reg_20_ ( .Q(s_frac2a_20_), .D(s_frac2a6207_20_), .CLK(clk_i)
         );
  dff s_frac2a_reg_19_ ( .Q(s_frac2a_19_), .D(s_frac2a6207_19_), .CLK(clk_i)
         );
  dff s_frac2a_reg_18_ ( .QB(n14497), .D(s_frac2a6207_18_), .CLK(clk_i) );
  dff s_frac2a_reg_17_ ( .QB(n14496), .D(s_frac2a6207_17_), .CLK(clk_i) );
  dff s_frac2a_reg_16_ ( .QB(n14495), .D(s_frac2a6207_16_), .CLK(clk_i) );
  dff s_frac2a_reg_15_ ( .Q(s_frac2a_15_), .D(s_frac2a6207_15_), .CLK(clk_i)
         );
  dff s_frac2a_reg_14_ ( .Q(s_frac2a_14_), .D(s_frac2a6207_14_), .CLK(clk_i)
         );
  dff s_frac2a_reg_13_ ( .Q(s_frac2a_13_), .D(s_frac2a6207_13_), .CLK(clk_i)
         );
  dff s_frac2a_reg_12_ ( .QB(n14499), .D(s_frac2a6207_12_), .CLK(clk_i) );
  dff s_frac2a_reg_11_ ( .QB(n14498), .D(s_frac2a6207_11_), .CLK(clk_i) );
  dff s_frac2a_reg_10_ ( .Q(s_frac2a_10_), .D(s_frac2a6207_10_), .CLK(clk_i)
         );
  dff s_frac2a_reg_9_ ( .QB(n14492), .D(s_frac2a6207_9_), .CLK(clk_i) );
  dff s_frac2a_reg_8_ ( .QB(n14491), .D(s_frac2a6207_8_), .CLK(clk_i) );
  dff s_frac2a_reg_7_ ( .QB(n14490), .D(s_frac2a6207_7_), .CLK(clk_i) );
  dff s_frac2a_reg_6_ ( .Q(s_frac2a_6_), .D(s_frac2a6207_6_), .CLK(clk_i) );
  dff s_frac2a_reg_5_ ( .Q(s_frac2a_5_), .D(s_frac2a6207_5_), .CLK(clk_i) );
  dff s_frac2a_reg_4_ ( .Q(s_frac2a_4_), .D(s_frac2a6207_4_), .CLK(clk_i) );
  dff s_frac2a_reg_3_ ( .QB(n14494), .D(s_frac2a6207_3_), .CLK(clk_i) );
  dff s_frac2a_reg_2_ ( .QB(n14493), .D(s_frac2a6207_2_), .CLK(clk_i) );
  dff s_frac2a_reg_1_ ( .Q(s_frac2a_1_), .D(s_frac2a6207_1_), .CLK(clk_i) );
  dff s_frac2a_reg_0_ ( .Q(s_frac2a_0_), .D(s_frac2a6207_0_), .CLK(clk_i) );
  dff s_frac_rnd_reg_24_ ( .Q(s_shr3), .D(n10226), .CLK(clk_i) );
  dff s_frac_rnd_reg_23_ ( .Q(s_frac_rnd_23_), .D(s_frac_rnd7043_23_), .CLK(
        clk_i) );
  dff s_frac_rnd_reg_22_ ( .Q(s_frac_rnd_22_), .D(n10227), .CLK(clk_i) );
  dff s_frac_rnd_reg_21_ ( .Q(n14407), .D(n10216), .CLK(clk_i) );
  dff s_frac_rnd_reg_20_ ( .Q(n14409), .D(n10211), .CLK(clk_i) );
  dff s_frac_rnd_reg_19_ ( .Q(n14410), .D(n10210), .CLK(clk_i) );
  dff s_frac_rnd_reg_18_ ( .Q(n14411), .D(n10228), .CLK(clk_i) );
  dff s_frac_rnd_reg_17_ ( .Q(n14412), .D(n10219), .CLK(clk_i) );
  dff s_frac_rnd_reg_16_ ( .Q(n14413), .D(n10214), .CLK(clk_i) );
  dff s_frac_rnd_reg_15_ ( .Q(n14414), .D(n10217), .CLK(clk_i) );
  dff s_frac_rnd_reg_14_ ( .Q(n14415), .D(n10225), .CLK(clk_i) );
  dff s_frac_rnd_reg_13_ ( .Q(n14416), .D(n10222), .CLK(clk_i) );
  dff s_frac_rnd_reg_12_ ( .Q(n14417), .D(n10207), .CLK(clk_i) );
  dff s_frac_rnd_reg_11_ ( .Q(n14419), .D(n10212), .CLK(clk_i) );
  dff s_frac_rnd_reg_10_ ( .Q(n14418), .D(n10208), .CLK(clk_i) );
  dff s_frac_rnd_reg_9_ ( .Q(n14400), .D(n10209), .CLK(clk_i) );
  dff s_frac_rnd_reg_8_ ( .Q(n14401), .D(n10224), .CLK(clk_i) );
  dff s_frac_rnd_reg_7_ ( .Q(n14402), .D(n10215), .CLK(clk_i) );
  dff s_frac_rnd_reg_6_ ( .Q(n14403), .D(n10220), .CLK(clk_i) );
  dff s_frac_rnd_reg_5_ ( .Q(n14404), .D(n10218), .CLK(clk_i) );
  dff s_frac_rnd_reg_4_ ( .Q(n14405), .D(n10221), .CLK(clk_i) );
  dff s_frac_rnd_reg_3_ ( .Q(n14406), .D(n10213), .CLK(clk_i) );
  dff s_frac_rnd_reg_2_ ( .Q(n14408), .D(n10223), .CLK(clk_i) );
  dff s_frac_rnd_reg_1_ ( .Q(s_frac_rnd_1_), .D(n10229), .CLK(clk_i) );
  dff s_frac_rnd_reg_0_ ( .QB(n14420), .D(s_frac_rnd7043_0_), .CLK(clk_i) );
  dff s_opa_i_reg_30_ ( .Q(s_opa_i_30_), .D(opa_i[30]), .CLK(clk_i) );
  dff s_opa_i_reg_29_ ( .Q(s_opa_i_29_), .D(opa_i[29]), .CLK(clk_i) );
  dff s_opa_i_reg_28_ ( .Q(s_opa_i_28_), .D(opa_i[28]), .CLK(clk_i) );
  dff s_opa_i_reg_27_ ( .QB(n14448), .D(opa_i[27]), .CLK(clk_i) );
  dff s_opa_i_reg_26_ ( .QB(n14447), .D(opa_i[26]), .CLK(clk_i) );
  dff s_opa_i_reg_25_ ( .Q(s_opa_i_25_), .D(opa_i[25]), .CLK(clk_i) );
  dff s_opa_i_reg_24_ ( .Q(s_opa_i_24_), .D(opa_i[24]), .CLK(clk_i) );
  dff s_opa_i_reg_23_ ( .Q(s_opa_i_23_), .D(opa_i[23]), .CLK(clk_i) );
  dff s_opa_i_reg_22_ ( .QB(n14439), .D(opa_i[22]), .CLK(clk_i) );
  dff s_opa_i_reg_21_ ( .Q(s_opa_i_21_), .D(opa_i[21]), .CLK(clk_i) );
  dff s_opa_i_reg_20_ ( .Q(s_opa_i_20_), .D(opa_i[20]), .CLK(clk_i) );
  dff s_opa_i_reg_19_ ( .QB(n14444), .D(opa_i[19]), .CLK(clk_i) );
  dff s_opa_i_reg_18_ ( .QB(n14443), .D(opa_i[18]), .CLK(clk_i) );
  dff s_opa_i_reg_17_ ( .QB(n14442), .D(opa_i[17]), .CLK(clk_i) );
  dff s_opa_i_reg_16_ ( .Q(s_opa_i_16_), .D(opa_i[16]), .CLK(clk_i) );
  dff s_opa_i_reg_15_ ( .Q(s_opa_i_15_), .D(opa_i[15]), .CLK(clk_i) );
  dff s_opa_i_reg_14_ ( .Q(s_opa_i_14_), .D(opa_i[14]), .CLK(clk_i) );
  dff s_opa_i_reg_13_ ( .QB(n14446), .D(opa_i[13]), .CLK(clk_i) );
  dff s_opa_i_reg_12_ ( .QB(n14445), .D(opa_i[12]), .CLK(clk_i) );
  dff s_opa_i_reg_11_ ( .Q(s_opa_i_11_), .D(opa_i[11]), .CLK(clk_i) );
  dff s_opa_i_reg_10_ ( .Q(s_opa_i_10_), .D(opa_i[10]), .CLK(clk_i) );
  dff s_opa_i_reg_9_ ( .QB(n14438), .D(opa_i[9]), .CLK(clk_i) );
  dff s_opa_i_reg_8_ ( .QB(n14437), .D(opa_i[8]), .CLK(clk_i) );
  dff s_opa_i_reg_7_ ( .QB(n14436), .D(opa_i[7]), .CLK(clk_i) );
  dff s_opa_i_reg_6_ ( .Q(s_opa_i_6_), .D(opa_i[6]), .CLK(clk_i) );
  dff s_opa_i_reg_5_ ( .Q(s_opa_i_5_), .D(opa_i[5]), .CLK(clk_i) );
  dff s_opa_i_reg_4_ ( .Q(s_opa_i_4_), .D(opa_i[4]), .CLK(clk_i) );
  dff s_opa_i_reg_3_ ( .QB(n14441), .D(opa_i[3]), .CLK(clk_i) );
  dff s_opa_i_reg_2_ ( .QB(n14440), .D(opa_i[2]), .CLK(clk_i) );
  dff s_opa_i_reg_1_ ( .Q(s_opa_i_1_), .D(opa_i[1]), .CLK(clk_i) );
  dff s_opa_i_reg_0_ ( .Q(s_opa_i_0_), .D(opa_i[0]), .CLK(clk_i) );
  dff s_opb_i_reg_30_ ( .Q(s_opb_i_30_), .D(opb_i[30]), .CLK(clk_i) );
  dff s_opb_i_reg_29_ ( .Q(s_opb_i_29_), .D(opb_i[29]), .CLK(clk_i) );
  dff s_opb_i_reg_28_ ( .Q(s_opb_i_28_), .D(opb_i[28]), .CLK(clk_i) );
  dff s_opb_i_reg_27_ ( .QB(n14435), .D(opb_i[27]), .CLK(clk_i) );
  dff s_opb_i_reg_26_ ( .QB(n14434), .D(opb_i[26]), .CLK(clk_i) );
  dff s_opb_i_reg_25_ ( .Q(s_opb_i_25_), .D(opb_i[25]), .CLK(clk_i) );
  dff s_opb_i_reg_24_ ( .Q(s_opb_i_24_), .D(opb_i[24]), .CLK(clk_i) );
  dff s_opb_i_reg_23_ ( .Q(s_opb_i_23_), .D(opb_i[23]), .CLK(clk_i) );
  dff s_opb_i_reg_22_ ( .QB(n14426), .D(opb_i[22]), .CLK(clk_i) );
  dff s_opb_i_reg_21_ ( .Q(s_opb_i_21_), .D(opb_i[21]), .CLK(clk_i) );
  dff s_opb_i_reg_20_ ( .Q(s_opb_i_20_), .D(opb_i[20]), .CLK(clk_i) );
  dff s_opb_i_reg_19_ ( .QB(n14431), .D(opb_i[19]), .CLK(clk_i) );
  dff s_opb_i_reg_18_ ( .QB(n14430), .D(opb_i[18]), .CLK(clk_i) );
  dff s_opb_i_reg_17_ ( .QB(n14429), .D(opb_i[17]), .CLK(clk_i) );
  dff s_opb_i_reg_16_ ( .Q(s_opb_i_16_), .D(opb_i[16]), .CLK(clk_i) );
  dff s_opb_i_reg_15_ ( .Q(s_opb_i_15_), .D(opb_i[15]), .CLK(clk_i) );
  dff s_opb_i_reg_14_ ( .Q(s_opb_i_14_), .D(opb_i[14]), .CLK(clk_i) );
  dff s_opb_i_reg_13_ ( .QB(n14433), .D(opb_i[13]), .CLK(clk_i) );
  dff s_opb_i_reg_12_ ( .QB(n14432), .D(opb_i[12]), .CLK(clk_i) );
  dff s_opb_i_reg_11_ ( .Q(s_opb_i_11_), .D(opb_i[11]), .CLK(clk_i) );
  dff s_opb_i_reg_10_ ( .Q(s_opb_i_10_), .D(opb_i[10]), .CLK(clk_i) );
  dff s_opb_i_reg_9_ ( .QB(n14425), .D(opb_i[9]), .CLK(clk_i) );
  dff s_opb_i_reg_8_ ( .QB(n14424), .D(opb_i[8]), .CLK(clk_i) );
  dff s_opb_i_reg_7_ ( .QB(n14423), .D(opb_i[7]), .CLK(clk_i) );
  dff s_opb_i_reg_6_ ( .Q(s_opb_i_6_), .D(opb_i[6]), .CLK(clk_i) );
  dff s_opb_i_reg_5_ ( .Q(s_opb_i_5_), .D(opb_i[5]), .CLK(clk_i) );
  dff s_opb_i_reg_4_ ( .Q(s_opb_i_4_), .D(opb_i[4]), .CLK(clk_i) );
  dff s_opb_i_reg_3_ ( .QB(n14428), .D(opb_i[3]), .CLK(clk_i) );
  dff s_opb_i_reg_2_ ( .QB(n14427), .D(opb_i[2]), .CLK(clk_i) );
  dff s_opb_i_reg_1_ ( .Q(s_opb_i_1_), .D(opb_i[1]), .CLK(clk_i) );
  dff s_opb_i_reg_0_ ( .Q(s_opb_i_0_), .D(opb_i[0]), .CLK(clk_i) );
  dff s_sign_i_reg ( .Q(s_sign_i), .QB(n14488), .D(sign_i), .CLK(clk_i) );
  dff ine_o_reg ( .Q(ine_o), .D(n10388), .CLK(clk_i) );
  inv02 U2545 ( .Y(n14352), .A(s_shr2_3_) );
  nor02 U2546 ( .Y(n9627), .A0(n14365), .A1(s_shl2_5_) );
  inv01 U2547 ( .Y(n9628), .A(n13580) );
  inv01 U2548 ( .Y(n9629), .A(n13580) );
  inv01 U2549 ( .Y(n9630), .A(n13580) );
  buf16 U2550 ( .Y(n13580), .A(n14106) );
  or03 U2551 ( .Y(n9631), .A0(n12408), .A1(n12350), .A2(n12462) );
  inv01 U2552 ( .Y(n9632), .A(n9631) );
  inv02 U2553 ( .Y(n13895), .A(n13830) );
  xor2 U2554 ( .Y(n9633), .A0(n12415), .A1(n13611) );
  inv01 U2555 ( .Y(n9634), .A(n9633) );
  xor2 U2556 ( .Y(n9635), .A0(n12449), .A1(n13607) );
  inv01 U2557 ( .Y(n9636), .A(n9635) );
  inv02 U2558 ( .Y(n13639), .A(n13736) );
  ao22 U2559 ( .Y(n9637), .A0(n13592), .A1(n10506), .B0(n13579), .B1(
        s_fract_48_i[44]) );
  inv01 U2560 ( .Y(n9638), .A(n9637) );
  ao22 U2561 ( .Y(n9639), .A0(n13593), .A1(n10290), .B0(n13590), .B1(n10885)
         );
  inv01 U2562 ( .Y(n9640), .A(n9639) );
  ao22 U2563 ( .Y(n9641), .A0(n13592), .A1(n10726), .B0(n13579), .B1(
        s_fract_48_i[22]) );
  inv01 U2564 ( .Y(n9642), .A(n9641) );
  ao22 U2565 ( .Y(n9643), .A0(n13593), .A1(n10506), .B0(n13588), .B1(
        s_fract_48_i[46]) );
  inv01 U2566 ( .Y(n9644), .A(n9643) );
  ao22 U2567 ( .Y(n9645), .A0(n13592), .A1(n12257), .B0(n13579), .B1(n10831)
         );
  inv01 U2568 ( .Y(n9646), .A(n9645) );
  ao22 U2569 ( .Y(n9647), .A0(n13593), .A1(n10286), .B0(n13586), .B1(
        s_fract_48_i[10]) );
  inv01 U2570 ( .Y(n9648), .A(n9647) );
  ao22 U2571 ( .Y(n9649), .A0(n13592), .A1(n10722), .B0(n13579), .B1(n12420)
         );
  inv01 U2572 ( .Y(n9650), .A(n9649) );
  ao22 U2573 ( .Y(n9651), .A0(n13593), .A1(n10575), .B0(n13586), .B1(
        s_fract_48_i[30]) );
  inv01 U2574 ( .Y(n9652), .A(n9651) );
  ao22 U2575 ( .Y(n9653), .A0(n13592), .A1(n10568), .B0(n13579), .B1(
        s_fract_48_i[17]) );
  inv01 U2576 ( .Y(n9654), .A(n9653) );
  ao22 U2577 ( .Y(n9655), .A0(n13592), .A1(n10288), .B0(n13579), .B1(n12925)
         );
  inv01 U2578 ( .Y(n9656), .A(n9655) );
  ao22 U2579 ( .Y(n9657), .A0(n13592), .A1(n10503), .B0(n13579), .B1(
        s_fract_48_i[14]) );
  inv01 U2580 ( .Y(n9658), .A(n9657) );
  ao22 U2581 ( .Y(n9659), .A0(n13592), .A1(n10292), .B0(n13579), .B1(
        s_fract_48_i[30]) );
  inv01 U2582 ( .Y(n9660), .A(n9659) );
  ao22 U2583 ( .Y(n9661), .A0(n13592), .A1(n10378), .B0(n13579), .B1(
        s_fract_48_i[6]) );
  inv01 U2584 ( .Y(n9662), .A(n9661) );
  ao22 U2585 ( .Y(n9663), .A0(n13592), .A1(n10882), .B0(n13579), .B1(
        s_fract_48_i[33]) );
  inv01 U2586 ( .Y(n9664), .A(n9663) );
  ao22 U2587 ( .Y(n9665), .A0(n13593), .A1(n10416), .B0(n13590), .B1(
        s_fract_48_i[14]) );
  inv01 U2588 ( .Y(n9666), .A(n9665) );
  ao22 U2589 ( .Y(n9667), .A0(n13593), .A1(n10377), .B0(n13590), .B1(n12923)
         );
  inv01 U2590 ( .Y(n9668), .A(n9667) );
  ao22 U2591 ( .Y(n9669), .A0(n13593), .A1(n10723), .B0(n13586), .B1(n12461)
         );
  inv01 U2592 ( .Y(n9670), .A(n9669) );
  ao22 U2593 ( .Y(n9671), .A0(n13592), .A1(n12889), .B0(n13579), .B1(
        s_fract_48_i[10]) );
  inv01 U2594 ( .Y(n9672), .A(n9671) );
  ao22 U2595 ( .Y(n9673), .A0(n13593), .A1(n12350), .B0(n13590), .B1(n10291)
         );
  inv01 U2596 ( .Y(n9674), .A(n9673) );
  ao22 U2597 ( .Y(n9675), .A0(n13592), .A1(n12252), .B0(n13579), .B1(n10293)
         );
  inv01 U2598 ( .Y(n9676), .A(n9675) );
  ao22 U2599 ( .Y(n9677), .A0(n13592), .A1(n10419), .B0(n13579), .B1(
        s_fract_48_i[12]) );
  inv01 U2600 ( .Y(n9678), .A(n9677) );
  ao22 U2601 ( .Y(n9679), .A0(n13592), .A1(n10819), .B0(n13579), .B1(n12254)
         );
  inv01 U2602 ( .Y(n9680), .A(n9679) );
  ao22 U2603 ( .Y(n9681), .A0(n13592), .A1(n12410), .B0(n13579), .B1(n12351)
         );
  inv01 U2604 ( .Y(n9682), .A(n9681) );
  ao22 U2605 ( .Y(n9683), .A0(n13593), .A1(n10501), .B0(n13588), .B1(n10571)
         );
  inv01 U2606 ( .Y(n9684), .A(n9683) );
  ao22 U2607 ( .Y(n9685), .A0(n13592), .A1(n10397), .B0(n13579), .B1(
        s_fract_48_i[43]) );
  inv01 U2608 ( .Y(n9686), .A(n9685) );
  ao22 U2609 ( .Y(n9687), .A0(n13592), .A1(n12348), .B0(n13579), .B1(n10572)
         );
  inv01 U2610 ( .Y(n9688), .A(n9687) );
  ao22 U2611 ( .Y(n9689), .A0(n13592), .A1(n10832), .B0(n13579), .B1(
        s_fract_48_i[38]) );
  inv01 U2612 ( .Y(n9690), .A(n9689) );
  ao22 U2613 ( .Y(n9691), .A0(n13592), .A1(n12420), .B0(n13579), .B1(n10725)
         );
  inv01 U2614 ( .Y(n9692), .A(n9691) );
  ao22 U2615 ( .Y(n9693), .A0(n13593), .A1(n10885), .B0(n13590), .B1(n10819)
         );
  inv01 U2616 ( .Y(n9694), .A(n9693) );
  nand02 U2617 ( .Y(n14314), .A0(n9695), .A1(n9696) );
  inv01 U2618 ( .Y(n9697), .A(n10719) );
  inv01 U2619 ( .Y(n9698), .A(n10571) );
  inv01 U2620 ( .Y(n9699), .A(n13593) );
  inv01 U2621 ( .Y(n9700), .A(n13588) );
  nand02 U2622 ( .Y(n9701), .A0(n9697), .A1(n9698) );
  nand02 U2623 ( .Y(n9702), .A0(n9697), .A1(n9699) );
  nand02 U2624 ( .Y(n9703), .A0(n9698), .A1(n9700) );
  nand02 U2625 ( .Y(n9704), .A0(n9699), .A1(n9700) );
  nand02 U2626 ( .Y(n9705), .A0(n9701), .A1(n9702) );
  inv01 U2627 ( .Y(n9695), .A(n9705) );
  nand02 U2628 ( .Y(n9706), .A0(n9703), .A1(n9704) );
  inv01 U2629 ( .Y(n9696), .A(n9706) );
  ao22 U2630 ( .Y(n9707), .A0(n13593), .A1(n10719), .B0(n13588), .B1(
        s_fract_48_i[22]) );
  inv01 U2631 ( .Y(n9708), .A(n9707) );
  ao22 U2632 ( .Y(n9709), .A0(n13593), .A1(n12462), .B0(n13586), .B1(n10574)
         );
  inv01 U2633 ( .Y(n9710), .A(n9709) );
  ao22 U2634 ( .Y(n9711), .A0(n13592), .A1(n10572), .B0(n13579), .B1(n12253)
         );
  inv01 U2635 ( .Y(n9712), .A(n9711) );
  ao22 U2636 ( .Y(n9713), .A0(n13592), .A1(n12461), .B0(n13579), .B1(n12410)
         );
  inv01 U2637 ( .Y(n9714), .A(n9713) );
  ao22 U2638 ( .Y(n9715), .A0(n13593), .A1(n10371), .B0(n13586), .B1(
        s_fract_48_i[15]) );
  inv01 U2639 ( .Y(n9716), .A(n9715) );
  ao22 U2640 ( .Y(n9717), .A0(n13593), .A1(n12250), .B0(n13588), .B1(
        s_fract_48_i[31]) );
  inv01 U2641 ( .Y(n9718), .A(n9717) );
  ao22 U2642 ( .Y(n9719), .A0(n13593), .A1(n12256), .B0(n13586), .B1(
        s_fract_48_i[39]) );
  inv01 U2643 ( .Y(n9720), .A(n9719) );
  ao22 U2644 ( .Y(n9721), .A0(n13593), .A1(n12411), .B0(n13588), .B1(n12252)
         );
  inv01 U2645 ( .Y(n9722), .A(n9721) );
  ao22 U2646 ( .Y(n9723), .A0(n13593), .A1(n10369), .B0(n13590), .B1(n10501)
         );
  inv01 U2647 ( .Y(n9724), .A(n9723) );
  nand02 U2648 ( .Y(n14219), .A0(n9725), .A1(n9726) );
  inv01 U2649 ( .Y(n9727), .A(n10287) );
  inv01 U2650 ( .Y(n9728), .A(n10370) );
  inv01 U2651 ( .Y(n9729), .A(n13592) );
  inv01 U2652 ( .Y(n9730), .A(n13579) );
  nand02 U2653 ( .Y(n9731), .A0(n9727), .A1(n9728) );
  nand02 U2654 ( .Y(n9732), .A0(n9727), .A1(n9729) );
  nand02 U2655 ( .Y(n9733), .A0(n9728), .A1(n9730) );
  nand02 U2656 ( .Y(n9734), .A0(n9729), .A1(n9730) );
  nand02 U2657 ( .Y(n9735), .A0(n9731), .A1(n9732) );
  inv01 U2658 ( .Y(n9725), .A(n9735) );
  nand02 U2659 ( .Y(n9736), .A0(n9733), .A1(n9734) );
  inv01 U2660 ( .Y(n9726), .A(n9736) );
  ao22 U2661 ( .Y(n9737), .A0(n13593), .A1(n10370), .B0(n13586), .B1(n12889)
         );
  inv01 U2662 ( .Y(n9738), .A(n9737) );
  ao22 U2663 ( .Y(n9739), .A0(n13592), .A1(n10371), .B0(n13579), .B1(n10504)
         );
  inv01 U2664 ( .Y(n9740), .A(n9739) );
  ao22 U2665 ( .Y(n9741), .A0(n13593), .A1(n12419), .B0(n13590), .B1(
        s_fract_48_i[23]) );
  inv01 U2666 ( .Y(n9742), .A(n9741) );
  ao22 U2667 ( .Y(n9743), .A0(n13593), .A1(n10398), .B0(n13586), .B1(
        s_fract_48_i[45]) );
  inv01 U2668 ( .Y(n9744), .A(n9743) );
  ao22 U2669 ( .Y(n9745), .A0(n13592), .A1(n10369), .B0(n13579), .B1(n10419)
         );
  inv01 U2670 ( .Y(n9746), .A(n9745) );
  ao22 U2671 ( .Y(n9747), .A0(n13592), .A1(n12922), .B0(n13579), .B1(n12888)
         );
  inv01 U2672 ( .Y(n9748), .A(n9747) );
  ao22 U2673 ( .Y(n9749), .A0(n13593), .A1(n12924), .B0(n13590), .B1(n10418)
         );
  inv01 U2674 ( .Y(n9750), .A(n9749) );
  ao22 U2675 ( .Y(n9751), .A0(n13593), .A1(n12887), .B0(n13586), .B1(
        s_fract_48_i[12]) );
  inv01 U2676 ( .Y(n9752), .A(n9751) );
  ao22 U2677 ( .Y(n9753), .A0(n13556), .A1(n14288), .B0(n13557), .B1(n14289)
         );
  inv01 U2678 ( .Y(n9754), .A(n9753) );
  xor2 U2679 ( .Y(n9755), .A0(n13605), .A1(n10401) );
  inv01 U2680 ( .Y(n9756), .A(n9755) );
  xor2 U2681 ( .Y(n9757), .A0(n____return5956_3_), .A1(n10161) );
  inv01 U2682 ( .Y(n9758), .A(n9757) );
  xor2 U2683 ( .Y(n9759), .A0(n____return5956_1_), .A1(n10099) );
  inv01 U2684 ( .Y(n9760), .A(n9759) );
  or02 U2685 ( .Y(n9761), .A0(n13514), .A1(n13885) );
  inv01 U2686 ( .Y(n9762), .A(n9761) );
  or02 U2687 ( .Y(n9763), .A0(n13514), .A1(n13903) );
  inv01 U2688 ( .Y(n9764), .A(n9763) );
  ao22 U2689 ( .Y(n9765), .A0(n13593), .A1(n10829), .B0(n13588), .B1(
        s_fract_48_i[40]) );
  inv01 U2690 ( .Y(n9766), .A(n9765) );
  ao22 U2691 ( .Y(n9767), .A0(n13593), .A1(n10821), .B0(n13590), .B1(
        s_fract_48_i[38]) );
  inv01 U2692 ( .Y(n9768), .A(n9767) );
  inv01 U2693 ( .Y(n13954), .A(n9769) );
  nor02 U2694 ( .Y(n9770), .A0(s_fract_48_i[46]), .A1(n10283) );
  nor02 U2695 ( .Y(n9771), .A0(n13938), .A1(n13745) );
  nor02 U2696 ( .Y(n9769), .A0(n9770), .A1(n9771) );
  ao22 U2697 ( .Y(n9772), .A0(n13564), .A1(n12809), .B0(n13573), .B1(n14069)
         );
  inv01 U2698 ( .Y(n9773), .A(n9772) );
  buf02 U2699 ( .Y(n9774), .A(n13443) );
  or02 U2700 ( .Y(n9775), .A0(n13513), .A1(n13869) );
  inv01 U2701 ( .Y(n9776), .A(n9775) );
  or02 U2702 ( .Y(n9777), .A0(n13513), .A1(n10848) );
  inv01 U2703 ( .Y(n9778), .A(n9777) );
  ao22 U2704 ( .Y(n9779), .A0(n13560), .A1(n14225), .B0(n13542), .B1(n14250)
         );
  inv01 U2705 ( .Y(n9780), .A(n9779) );
  xor2 U2706 ( .Y(n9781), .A0(s_rmode_i_0_), .A1(n14488) );
  inv01 U2707 ( .Y(n9782), .A(n9781) );
  ao22 U2708 ( .Y(n9783), .A0(n13560), .A1(n14216), .B0(n13542), .B1(n14237)
         );
  inv01 U2709 ( .Y(n9784), .A(n9783) );
  ao22 U2710 ( .Y(n9785), .A0(n13560), .A1(n14211), .B0(n13542), .B1(n14235)
         );
  inv01 U2711 ( .Y(n9786), .A(n9785) );
  ao22 U2712 ( .Y(n9787), .A0(n13560), .A1(n14229), .B0(n13542), .B1(n14267)
         );
  inv01 U2713 ( .Y(n9788), .A(n9787) );
  ao22 U2714 ( .Y(n9789), .A0(n13560), .A1(n14235), .B0(n13542), .B1(n14280)
         );
  inv01 U2715 ( .Y(n9790), .A(n9789) );
  ao22 U2716 ( .Y(n9791), .A0(n13560), .A1(n14237), .B0(n13542), .B1(n14291)
         );
  inv01 U2717 ( .Y(n9792), .A(n9791) );
  ao22 U2718 ( .Y(n9793), .A0(n13560), .A1(n14189), .B0(n13542), .B1(n14216)
         );
  inv01 U2719 ( .Y(n9794), .A(n9793) );
  ao22 U2720 ( .Y(n9795), .A0(n13560), .A1(n14183), .B0(n13542), .B1(n14211)
         );
  inv01 U2721 ( .Y(n9796), .A(n9795) );
  ao22 U2722 ( .Y(n9797), .A0(n13560), .A1(n14203), .B0(n13542), .B1(n14229)
         );
  inv01 U2723 ( .Y(n9798), .A(n9797) );
  ao22 U2724 ( .Y(n9799), .A0(n13964), .A1(n13513), .B0(n13965), .B1(n13769)
         );
  inv01 U2725 ( .Y(n9800), .A(n9799) );
  ao22 U2726 ( .Y(n9801), .A0(n13560), .A1(n14194), .B0(n13542), .B1(n14225)
         );
  inv01 U2727 ( .Y(n9802), .A(n9801) );
  ao22 U2728 ( .Y(n9803), .A0(n13576), .A1(n14248), .B0(n13556), .B1(n14124)
         );
  inv01 U2729 ( .Y(n9804), .A(n9803) );
  ao22 U2730 ( .Y(n9805), .A0(n13576), .A1(n14278), .B0(n13556), .B1(n14318)
         );
  inv01 U2731 ( .Y(n9806), .A(n9805) );
  ao22 U2732 ( .Y(n9807), .A0(n13542), .A1(n14240), .B0(n13560), .B1(n14250)
         );
  inv01 U2733 ( .Y(n9808), .A(n9807) );
  ao22 U2734 ( .Y(n9809), .A0(s_shr2_1_), .A1(n14398), .B0(n13579), .B1(s_shr3) );
  inv01 U2735 ( .Y(n9810), .A(n9809) );
  nand02 U2736 ( .Y(n14331), .A0(n9811), .A1(n9812) );
  inv01 U2737 ( .Y(n9813), .A(n14267) );
  inv01 U2738 ( .Y(n9814), .A(n14256) );
  inv01 U2739 ( .Y(n9815), .A(n13560) );
  inv01 U2740 ( .Y(n9816), .A(n13566) );
  nand02 U2741 ( .Y(n9817), .A0(n9813), .A1(n9814) );
  nand02 U2742 ( .Y(n9818), .A0(n9813), .A1(n9815) );
  nand02 U2743 ( .Y(n9819), .A0(n9814), .A1(n9816) );
  nand02 U2744 ( .Y(n9820), .A0(n9815), .A1(n9816) );
  nand02 U2745 ( .Y(n9821), .A0(n9817), .A1(n9818) );
  inv01 U2746 ( .Y(n9811), .A(n9821) );
  nand02 U2747 ( .Y(n9822), .A0(n9819), .A1(n9820) );
  inv01 U2748 ( .Y(n9812), .A(n9822) );
  ao22 U2749 ( .Y(n9823), .A0(n13542), .A1(n14256), .B0(n13560), .B1(n14267)
         );
  inv01 U2750 ( .Y(n9824), .A(n9823) );
  ao22 U2751 ( .Y(n9825), .A0(n13564), .A1(n14196), .B0(n13569), .B1(n14330)
         );
  inv01 U2752 ( .Y(n9826), .A(n9825) );
  ao22 U2753 ( .Y(n9827), .A0(n13593), .A1(s_fract_48_i[1]), .B0(n13588), .B1(
        s_fract_48_i[4]) );
  inv01 U2754 ( .Y(n9828), .A(n9827) );
  ao22 U2755 ( .Y(n9829), .A0(n13561), .A1(n14277), .B0(n13556), .B1(n14278)
         );
  inv01 U2756 ( .Y(n9830), .A(n9829) );
  ao22 U2757 ( .Y(n9831), .A0(n13561), .A1(n14289), .B0(n13556), .B1(n14324)
         );
  inv01 U2758 ( .Y(n9832), .A(n9831) );
  nand02 U2759 ( .Y(n14295), .A0(n9833), .A1(n9834) );
  inv01 U2760 ( .Y(n9835), .A(n14248) );
  inv01 U2761 ( .Y(n9836), .A(n14247) );
  inv01 U2762 ( .Y(n9837), .A(n13561) );
  inv01 U2763 ( .Y(n9838), .A(n13556) );
  nand02 U2764 ( .Y(n9839), .A0(n9835), .A1(n9836) );
  nand02 U2765 ( .Y(n9840), .A0(n9835), .A1(n9837) );
  nand02 U2766 ( .Y(n9841), .A0(n9836), .A1(n9838) );
  nand02 U2767 ( .Y(n9842), .A0(n9837), .A1(n9838) );
  nand02 U2768 ( .Y(n9843), .A0(n9839), .A1(n9840) );
  inv01 U2769 ( .Y(n9833), .A(n9843) );
  nand02 U2770 ( .Y(n9844), .A0(n9841), .A1(n9842) );
  inv01 U2771 ( .Y(n9834), .A(n9844) );
  ao22 U2772 ( .Y(n9845), .A0(n13556), .A1(n14247), .B0(n13561), .B1(n14296)
         );
  inv01 U2773 ( .Y(n9846), .A(n9845) );
  nand02 U2774 ( .Y(n14368), .A0(n9847), .A1(n9848) );
  inv01 U2775 ( .Y(n9849), .A(n14265) );
  inv01 U2776 ( .Y(n9850), .A(n14264) );
  inv01 U2777 ( .Y(n9851), .A(n13576) );
  inv01 U2778 ( .Y(n9852), .A(n13557) );
  nand02 U2779 ( .Y(n9853), .A0(n9849), .A1(n9850) );
  nand02 U2780 ( .Y(n9854), .A0(n9849), .A1(n9851) );
  nand02 U2781 ( .Y(n9855), .A0(n9850), .A1(n9852) );
  nand02 U2782 ( .Y(n9856), .A0(n9851), .A1(n9852) );
  nand02 U2783 ( .Y(n9857), .A0(n9853), .A1(n9854) );
  inv01 U2784 ( .Y(n9847), .A(n9857) );
  nand02 U2785 ( .Y(n9858), .A0(n9855), .A1(n9856) );
  inv01 U2786 ( .Y(n9848), .A(n9858) );
  ao22 U2787 ( .Y(n9859), .A0(n13556), .A1(n14264), .B0(n13557), .B1(n14259)
         );
  inv01 U2788 ( .Y(n9860), .A(n9859) );
  ao22 U2789 ( .Y(n9861), .A0(n13566), .A1(n14250), .B0(n13560), .B1(n14240)
         );
  inv01 U2790 ( .Y(n9862), .A(n9861) );
  ao22 U2791 ( .Y(n9863), .A0(n13560), .A1(n14282), .B0(n13566), .B1(n14291)
         );
  inv01 U2792 ( .Y(n9864), .A(n9863) );
  ao22 U2793 ( .Y(n9865), .A0(n13556), .A1(n14284), .B0(n13557), .B1(n14288)
         );
  inv01 U2794 ( .Y(n9866), .A(n9865) );
  inv01 U2795 ( .Y(n14354), .A(n9867) );
  nor02 U2796 ( .Y(n9868), .A0(n13527), .A1(n14233) );
  nor02 U2797 ( .Y(n9869), .A0(n13563), .A1(n12917) );
  nor02 U2798 ( .Y(n9867), .A0(n9868), .A1(n9869) );
  ao22 U2799 ( .Y(n9870), .A0(n13542), .A1(n14282), .B0(n13560), .B1(n14291)
         );
  inv01 U2800 ( .Y(n9871), .A(n9870) );
  inv02 U2801 ( .Y(n13527), .A(n13565) );
  ao22 U2802 ( .Y(n9872), .A0(n13010), .A1(n13556), .B0(n13561), .B1(n14318)
         );
  inv01 U2803 ( .Y(n9873), .A(n9872) );
  ao22 U2804 ( .Y(n9874), .A0(n13566), .A1(n14280), .B0(n13560), .B1(n14269)
         );
  inv01 U2805 ( .Y(n9875), .A(n9874) );
  xor2 U2806 ( .Y(n9876), .A0(n____return6004_6_), .A1(n13963) );
  inv01 U2807 ( .Y(n9877), .A(n9876) );
  ao22 U2808 ( .Y(n9878), .A0(n14271), .A1(s_shr2_2_), .B0(n14273), .B1(n14353) );
  inv01 U2809 ( .Y(n9879), .A(n9878) );
  ao22 U2810 ( .Y(n9880), .A0(n12921), .A1(n14132), .B0(n13565), .B1(n14134)
         );
  inv01 U2811 ( .Y(n9881), .A(n9880) );
  ao22 U2812 ( .Y(n9882), .A0(n14255), .A1(s_shl2_2_), .B0(n14254), .B1(n14300) );
  inv01 U2813 ( .Y(n9883), .A(n9882) );
  ao22 U2814 ( .Y(n9884), .A0(n13593), .A1(s_fract_48_i[2]), .B0(n13588), .B1(
        n10376) );
  inv01 U2815 ( .Y(n9885), .A(n9884) );
  ao22 U2816 ( .Y(n9886), .A0(n13542), .A1(n14269), .B0(n13560), .B1(n14280)
         );
  inv01 U2817 ( .Y(n9887), .A(n9886) );
  buf02 U2818 ( .Y(n9888), .A(n14373) );
  ao22 U2819 ( .Y(n9889), .A0(n13569), .A1(n14309), .B0(n13564), .B1(n14191)
         );
  inv01 U2820 ( .Y(n9890), .A(n9889) );
  ao22 U2821 ( .Y(n9891), .A0(n13569), .A1(n14166), .B0(n13565), .B1(n14182)
         );
  inv01 U2822 ( .Y(n9892), .A(n9891) );
  ao22 U2823 ( .Y(n9893), .A0(n13569), .A1(n14220), .B0(n13564), .B1(n14185)
         );
  inv01 U2824 ( .Y(n9894), .A(n9893) );
  ao22 U2825 ( .Y(n9895), .A0(n13556), .A1(n14345), .B0(n13557), .B1(n14264)
         );
  inv01 U2826 ( .Y(n9896), .A(n9895) );
  ao22 U2827 ( .Y(n9897), .A0(n13593), .A1(s_fract_48_i[3]), .B0(n13588), .B1(
        s_fract_48_i[6]) );
  inv01 U2828 ( .Y(n9898), .A(n9897) );
  or02 U2829 ( .Y(n9899), .A0(n13511), .A1(n10846) );
  inv01 U2830 ( .Y(n9900), .A(n9899) );
  ao22 U2831 ( .Y(n9901), .A0(n13593), .A1(s_fract_48_i[4]), .B0(n13588), .B1(
        n10289) );
  inv01 U2832 ( .Y(n9902), .A(n9901) );
  ao22 U2833 ( .Y(n9903), .A0(s_fract_48_i[0]), .A1(n14108), .B0(n13586), .B1(
        s_fract_48_i[3]) );
  inv01 U2834 ( .Y(n9904), .A(n9903) );
  buf02 U2835 ( .Y(n9905), .A(n14374) );
  ao22 U2836 ( .Y(n9906), .A0(n13561), .A1(n14259), .B0(n13556), .B1(n14261)
         );
  inv01 U2837 ( .Y(n9907), .A(n9906) );
  nand02 U2838 ( .Y(n14188), .A0(n9908), .A1(n9909) );
  inv01 U2839 ( .Y(n9910), .A(s_fract_48_i[34]) );
  inv01 U2840 ( .Y(n9911), .A(s_fract_48_i[31]) );
  inv01 U2841 ( .Y(n9912), .A(n13593) );
  inv01 U2842 ( .Y(n9913), .A(n13588) );
  nand02 U2843 ( .Y(n9914), .A0(n9910), .A1(n9911) );
  nand02 U2844 ( .Y(n9915), .A0(n9910), .A1(n9912) );
  nand02 U2845 ( .Y(n9916), .A0(n9911), .A1(n9913) );
  nand02 U2846 ( .Y(n9917), .A0(n9912), .A1(n9913) );
  nand02 U2847 ( .Y(n9918), .A0(n9914), .A1(n9915) );
  inv01 U2848 ( .Y(n9908), .A(n9918) );
  nand02 U2849 ( .Y(n9919), .A0(n9916), .A1(n9917) );
  inv01 U2850 ( .Y(n9909), .A(n9919) );
  ao22 U2851 ( .Y(n9920), .A0(n13592), .A1(s_fract_48_i[31]), .B0(n13579), 
        .B1(n10884) );
  inv01 U2852 ( .Y(n9921), .A(n9920) );
  ao22 U2853 ( .Y(n9922), .A0(n13556), .A1(n14245), .B0(n13557), .B1(n14247)
         );
  inv01 U2854 ( .Y(n9923), .A(n9922) );
  ao22 U2855 ( .Y(n9924), .A0(n13556), .A1(n14276), .B0(n13557), .B1(n14277)
         );
  inv01 U2856 ( .Y(n9925), .A(n9924) );
  ao22 U2857 ( .Y(n9926), .A0(n13565), .A1(n14142), .B0(n13573), .B1(n14141)
         );
  inv01 U2858 ( .Y(n9927), .A(n9926) );
  ao22 U2859 ( .Y(n9928), .A0(n13565), .A1(n14148), .B0(n13573), .B1(n14147)
         );
  inv01 U2860 ( .Y(n9929), .A(n9928) );
  ao22 U2861 ( .Y(n9930), .A0(n14010), .A1(n13994), .B0(n10304), .B1(n13995)
         );
  inv01 U2862 ( .Y(n9931), .A(n9930) );
  nand02 U2863 ( .Y(n14149), .A0(n9932), .A1(n9933) );
  inv01 U2864 ( .Y(n9934), .A(n10395) );
  inv01 U2865 ( .Y(n9935), .A(s_fract_48_i[39]) );
  inv01 U2866 ( .Y(n9936), .A(n13593) );
  inv01 U2867 ( .Y(n9937), .A(n13586) );
  nand02 U2868 ( .Y(n9938), .A0(n9934), .A1(n9935) );
  nand02 U2869 ( .Y(n9939), .A0(n9934), .A1(n9936) );
  nand02 U2870 ( .Y(n9940), .A0(n9935), .A1(n9937) );
  nand02 U2871 ( .Y(n9941), .A0(n9936), .A1(n9937) );
  nand02 U2872 ( .Y(n9942), .A0(n9938), .A1(n9939) );
  inv01 U2873 ( .Y(n9932), .A(n9942) );
  nand02 U2874 ( .Y(n9943), .A0(n9940), .A1(n9941) );
  inv01 U2875 ( .Y(n9933), .A(n9943) );
  ao22 U2876 ( .Y(n9944), .A0(n13592), .A1(s_fract_48_i[39]), .B0(n13579), 
        .B1(s_fract_48_i[40]) );
  inv01 U2877 ( .Y(n9945), .A(n9944) );
  ao22 U2878 ( .Y(n9946), .A0(n13593), .A1(s_fract_48_i[30]), .B0(n13586), 
        .B1(s_fract_48_i[33]) );
  inv01 U2879 ( .Y(n9947), .A(n9946) );
  ao22 U2880 ( .Y(n9948), .A0(n13592), .A1(s_fract_48_i[30]), .B0(n13579), 
        .B1(s_fract_48_i[31]) );
  inv01 U2881 ( .Y(n9949), .A(n9948) );
  nand02 U2882 ( .Y(n14351), .A0(n9950), .A1(n9951) );
  inv01 U2883 ( .Y(n9952), .A(n10570) );
  inv01 U2884 ( .Y(n9953), .A(s_fract_48_i[15]) );
  inv01 U2885 ( .Y(n9954), .A(n13592) );
  inv01 U2886 ( .Y(n9955), .A(n13579) );
  nand02 U2887 ( .Y(n9956), .A0(n9952), .A1(n9953) );
  nand02 U2888 ( .Y(n9957), .A0(n9952), .A1(n9954) );
  nand02 U2889 ( .Y(n9958), .A0(n9953), .A1(n9955) );
  nand02 U2890 ( .Y(n9959), .A0(n9954), .A1(n9955) );
  nand02 U2891 ( .Y(n9960), .A0(n9956), .A1(n9957) );
  inv01 U2892 ( .Y(n9950), .A(n9960) );
  nand02 U2893 ( .Y(n9961), .A0(n9958), .A1(n9959) );
  inv01 U2894 ( .Y(n9951), .A(n9961) );
  ao22 U2895 ( .Y(n9962), .A0(n13593), .A1(s_fract_48_i[15]), .B0(n13586), 
        .B1(s_fract_48_i[18]) );
  inv01 U2896 ( .Y(n9963), .A(n9962) );
  ao22 U2897 ( .Y(n9964), .A0(n13556), .A1(n14116), .B0(n13561), .B1(n14284)
         );
  inv01 U2898 ( .Y(n9965), .A(n9964) );
  nand02 U2899 ( .Y(n14363), .A0(n9966), .A1(n9967) );
  inv01 U2900 ( .Y(n9968), .A(n10822) );
  inv01 U2901 ( .Y(n9969), .A(s_fract_48_i[34]) );
  inv01 U2902 ( .Y(n9970), .A(n13592) );
  inv01 U2903 ( .Y(n9971), .A(n13579) );
  nand02 U2904 ( .Y(n9972), .A0(n9968), .A1(n9969) );
  nand02 U2905 ( .Y(n9973), .A0(n9968), .A1(n9970) );
  nand02 U2906 ( .Y(n9974), .A0(n9969), .A1(n9971) );
  nand02 U2907 ( .Y(n9975), .A0(n9970), .A1(n9971) );
  nand02 U2908 ( .Y(n9976), .A0(n9972), .A1(n9973) );
  inv01 U2909 ( .Y(n9966), .A(n9976) );
  nand02 U2910 ( .Y(n9977), .A0(n9974), .A1(n9975) );
  inv01 U2911 ( .Y(n9967), .A(n9977) );
  ao22 U2912 ( .Y(n9978), .A0(n13593), .A1(s_fract_48_i[34]), .B0(n13588), 
        .B1(n10832) );
  inv01 U2913 ( .Y(n9979), .A(n9978) );
  ao22 U2914 ( .Y(n9980), .A0(n12921), .A1(n14124), .B0(n13565), .B1(n14126)
         );
  inv01 U2915 ( .Y(n9981), .A(n9980) );
  ao22 U2916 ( .Y(n9982), .A0(n13593), .A1(s_fract_48_i[23]), .B0(n13590), 
        .B1(n12348) );
  inv01 U2917 ( .Y(n9983), .A(n9982) );
  nand02 U2918 ( .Y(n14305), .A0(n9984), .A1(n9985) );
  inv01 U2919 ( .Y(n9986), .A(n12417) );
  inv01 U2920 ( .Y(n9987), .A(s_fract_48_i[17]) );
  inv01 U2921 ( .Y(n9988), .A(n13593) );
  inv01 U2922 ( .Y(n9989), .A(n13590) );
  nand02 U2923 ( .Y(n9990), .A0(n9986), .A1(n9987) );
  nand02 U2924 ( .Y(n9991), .A0(n9986), .A1(n9988) );
  nand02 U2925 ( .Y(n9992), .A0(n9987), .A1(n9989) );
  nand02 U2926 ( .Y(n9993), .A0(n9988), .A1(n9989) );
  nand02 U2927 ( .Y(n9994), .A0(n9990), .A1(n9991) );
  inv01 U2928 ( .Y(n9984), .A(n9994) );
  nand02 U2929 ( .Y(n9995), .A0(n9992), .A1(n9993) );
  inv01 U2930 ( .Y(n9985), .A(n9995) );
  ao22 U2931 ( .Y(n9996), .A0(n13592), .A1(s_fract_48_i[17]), .B0(n13579), 
        .B1(s_fract_48_i[18]) );
  inv01 U2932 ( .Y(n9997), .A(n9996) );
  ao22 U2933 ( .Y(n9998), .A0(n13592), .A1(s_fract_48_i[41]), .B0(n13579), 
        .B1(n10397) );
  inv01 U2934 ( .Y(n9999), .A(n9998) );
  ao22 U2935 ( .Y(n10000), .A0(n13592), .A1(s_fract_48_i[23]), .B0(n13579), 
        .B1(n12459) );
  inv01 U2936 ( .Y(n10001), .A(n10000) );
  ao22 U2937 ( .Y(n10002), .A0(n13593), .A1(s_fract_48_i[41]), .B0(n13590), 
        .B1(s_fract_48_i[44]) );
  inv01 U2938 ( .Y(n10003), .A(n10002) );
  nand02 U2939 ( .Y(n14251), .A0(n10004), .A1(n10005) );
  inv01 U2940 ( .Y(n10006), .A(n12408) );
  inv01 U2941 ( .Y(n10007), .A(s_fract_48_i[22]) );
  inv01 U2942 ( .Y(n10008), .A(n13593) );
  inv01 U2943 ( .Y(n10009), .A(n13588) );
  nand02 U2944 ( .Y(n10010), .A0(n10006), .A1(n10007) );
  nand02 U2945 ( .Y(n10011), .A0(n10006), .A1(n10008) );
  nand02 U2946 ( .Y(n10012), .A0(n10007), .A1(n10009) );
  nand02 U2947 ( .Y(n10013), .A0(n10008), .A1(n10009) );
  nand02 U2948 ( .Y(n10014), .A0(n10010), .A1(n10011) );
  inv01 U2949 ( .Y(n10004), .A(n10014) );
  nand02 U2950 ( .Y(n10015), .A0(n10012), .A1(n10013) );
  inv01 U2951 ( .Y(n10005), .A(n10015) );
  nand02 U2952 ( .Y(n14358), .A0(n10016), .A1(n10017) );
  inv01 U2953 ( .Y(n10018), .A(s_fract_48_i[15]) );
  inv01 U2954 ( .Y(n10019), .A(s_fract_48_i[14]) );
  inv01 U2955 ( .Y(n10020), .A(n13592) );
  inv01 U2956 ( .Y(n10021), .A(n13579) );
  nand02 U2957 ( .Y(n10022), .A0(n10018), .A1(n10019) );
  nand02 U2958 ( .Y(n10023), .A0(n10018), .A1(n10020) );
  nand02 U2959 ( .Y(n10024), .A0(n10019), .A1(n10021) );
  nand02 U2960 ( .Y(n10025), .A0(n10020), .A1(n10021) );
  nand02 U2961 ( .Y(n10026), .A0(n10022), .A1(n10023) );
  inv01 U2962 ( .Y(n10016), .A(n10026) );
  nand02 U2963 ( .Y(n10027), .A0(n10024), .A1(n10025) );
  inv01 U2964 ( .Y(n10017), .A(n10027) );
  ao22 U2965 ( .Y(n10028), .A0(n13592), .A1(s_fract_48_i[22]), .B0(n13579), 
        .B1(s_fract_48_i[23]) );
  inv01 U2966 ( .Y(n10029), .A(n10028) );
  ao22 U2967 ( .Y(n10030), .A0(n13593), .A1(s_fract_48_i[14]), .B0(n13590), 
        .B1(s_fract_48_i[17]) );
  inv01 U2968 ( .Y(n10031), .A(n10030) );
  ao22 U2969 ( .Y(n10032), .A0(n13592), .A1(s_fract_48_i[18]), .B0(n13579), 
        .B1(n10721) );
  inv01 U2970 ( .Y(n10033), .A(n10032) );
  nand02 U2971 ( .Y(n14179), .A0(n10034), .A1(n10035) );
  inv01 U2972 ( .Y(n10036), .A(n12257) );
  inv01 U2973 ( .Y(n10037), .A(s_fract_48_i[33]) );
  inv01 U2974 ( .Y(n10038), .A(n13593) );
  inv01 U2975 ( .Y(n10039), .A(n13586) );
  nand02 U2976 ( .Y(n10040), .A0(n10036), .A1(n10037) );
  nand02 U2977 ( .Y(n10041), .A0(n10036), .A1(n10038) );
  nand02 U2978 ( .Y(n10042), .A0(n10037), .A1(n10039) );
  nand02 U2979 ( .Y(n10043), .A0(n10038), .A1(n10039) );
  nand02 U2980 ( .Y(n10044), .A0(n10040), .A1(n10041) );
  inv01 U2981 ( .Y(n10034), .A(n10044) );
  nand02 U2982 ( .Y(n10045), .A0(n10042), .A1(n10043) );
  inv01 U2983 ( .Y(n10035), .A(n10045) );
  ao22 U2984 ( .Y(n10046), .A0(n13592), .A1(s_fract_48_i[33]), .B0(n13579), 
        .B1(s_fract_48_i[34]) );
  inv01 U2985 ( .Y(n10047), .A(n10046) );
  nand02 U2986 ( .Y(n14107), .A0(n10048), .A1(n10049) );
  inv01 U2987 ( .Y(n10050), .A(n13514) );
  inv01 U2988 ( .Y(n10051), .A(s_fract_48_i[44]) );
  inv01 U2989 ( .Y(n10052), .A(n13593) );
  inv01 U2990 ( .Y(n10053), .A(n13590) );
  nand02 U2991 ( .Y(n10054), .A0(n10050), .A1(n10051) );
  nand02 U2992 ( .Y(n10055), .A0(n10050), .A1(n10052) );
  nand02 U2993 ( .Y(n10056), .A0(n10051), .A1(n10053) );
  nand02 U2994 ( .Y(n10057), .A0(n10052), .A1(n10053) );
  nand02 U2995 ( .Y(n10058), .A0(n10054), .A1(n10055) );
  inv01 U2996 ( .Y(n10048), .A(n10058) );
  nand02 U2997 ( .Y(n10059), .A0(n10056), .A1(n10057) );
  inv01 U2998 ( .Y(n10049), .A(n10059) );
  ao22 U2999 ( .Y(n10060), .A0(n13592), .A1(s_fract_48_i[44]), .B0(n13579), 
        .B1(s_fract_48_i[45]) );
  inv01 U3000 ( .Y(n10061), .A(n10060) );
  ao22 U3001 ( .Y(n10062), .A0(n13592), .A1(s_fract_48_i[4]), .B0(n13579), 
        .B1(n10375) );
  inv01 U3002 ( .Y(n10063), .A(n10062) );
  ao22 U3003 ( .Y(n10064), .A0(n13593), .A1(s_fract_48_i[18]), .B0(n13586), 
        .B1(n10723) );
  inv01 U3004 ( .Y(n10065), .A(n10064) );
  ao22 U3005 ( .Y(n10066), .A0(n13593), .A1(s_fract_48_i[38]), .B0(n13590), 
        .B1(s_fract_48_i[41]) );
  inv01 U3006 ( .Y(n10067), .A(n10066) );
  inv02 U3007 ( .Y(n14300), .A(s_shl2_2_) );
  ao22 U3008 ( .Y(n10068), .A0(n13592), .A1(s_fract_48_i[38]), .B0(n13579), 
        .B1(s_fract_48_i[39]) );
  inv01 U3009 ( .Y(n10069), .A(n10068) );
  nand02 U3010 ( .Y(n14143), .A0(n10070), .A1(n10071) );
  inv01 U3011 ( .Y(n10072), .A(s_fract_48_i[43]) );
  inv01 U3012 ( .Y(n10073), .A(s_fract_48_i[40]) );
  inv01 U3013 ( .Y(n10074), .A(n13593) );
  inv01 U3014 ( .Y(n10075), .A(n13588) );
  nand02 U3015 ( .Y(n10076), .A0(n10072), .A1(n10073) );
  nand02 U3016 ( .Y(n10077), .A0(n10072), .A1(n10074) );
  nand02 U3017 ( .Y(n10078), .A0(n10073), .A1(n10075) );
  nand02 U3018 ( .Y(n10079), .A0(n10074), .A1(n10075) );
  nand02 U3019 ( .Y(n10080), .A0(n10076), .A1(n10077) );
  inv01 U3020 ( .Y(n10070), .A(n10080) );
  nand02 U3021 ( .Y(n10081), .A0(n10078), .A1(n10079) );
  inv01 U3022 ( .Y(n10071), .A(n10081) );
  ao22 U3023 ( .Y(n10082), .A0(n13592), .A1(s_fract_48_i[40]), .B0(n13579), 
        .B1(s_fract_48_i[41]) );
  inv01 U3024 ( .Y(n10083), .A(n10082) );
  nand02 U3025 ( .Y(n14355), .A0(n10084), .A1(n10085) );
  inv01 U3026 ( .Y(n10086), .A(n14272) );
  inv01 U3027 ( .Y(n10087), .A(n14338) );
  inv01 U3028 ( .Y(n10088), .A(n14317) );
  inv01 U3029 ( .Y(n10089), .A(n13562) );
  nand02 U3030 ( .Y(n10084), .A0(n10086), .A1(n10087) );
  nand02 U3031 ( .Y(n10085), .A0(n10088), .A1(n10089) );
  nand02 U3032 ( .Y(n14362), .A0(n10090), .A1(n10091) );
  inv01 U3033 ( .Y(n10092), .A(n14322) );
  inv01 U3034 ( .Y(n10093), .A(n14338) );
  inv01 U3035 ( .Y(n10094), .A(n14321) );
  inv01 U3036 ( .Y(n10095), .A(n13562) );
  nand02 U3037 ( .Y(n10090), .A0(n10092), .A1(n10093) );
  nand02 U3038 ( .Y(n10091), .A0(n10094), .A1(n10095) );
  inv01 U3039 ( .Y(n14337), .A(n10096) );
  nor02 U3040 ( .Y(n10097), .A0(n14338), .A1(n13418) );
  nor02 U3041 ( .Y(n10098), .A0(n13562), .A1(n14293) );
  nor02 U3042 ( .Y(n10096), .A0(n10097), .A1(n10098) );
  nand02 U3043 ( .Y(n10099), .A0(n____return5956_0_), .A1(n13511) );
  inv01 U3044 ( .Y(n14347), .A(n10100) );
  nor02 U3045 ( .Y(n10101), .A0(n14199), .A1(n14254) );
  nor02 U3046 ( .Y(n10102), .A0(n14204), .A1(n14255) );
  nor02 U3047 ( .Y(n10100), .A0(n10101), .A1(n10102) );
  inv01 U3048 ( .Y(n14341), .A(n10103) );
  nor02 U3049 ( .Y(n10104), .A0(n14204), .A1(n13394) );
  nor02 U3050 ( .Y(n10105), .A0(n14199), .A1(n13423) );
  nor02 U3051 ( .Y(n10103), .A0(n10104), .A1(n10105) );
  inv02 U3052 ( .Y(n14204), .A(n13542) );
  buf12 U3053 ( .Y(n13572), .A(n14221) );
  ao22 U3054 ( .Y(n10106), .A0(n10275), .A1(n13565), .B0(n13547), .B1(n14063)
         );
  inv01 U3055 ( .Y(n10107), .A(n10106) );
  ao22 U3056 ( .Y(n10108), .A0(n13565), .A1(n12753), .B0(n13541), .B1(n14091)
         );
  inv01 U3057 ( .Y(n10109), .A(n10108) );
  ao22 U3058 ( .Y(n10110), .A0(n13564), .A1(n14361), .B0(n13549), .B1(n14081)
         );
  inv01 U3059 ( .Y(n10111), .A(n10110) );
  ao22 U3060 ( .Y(n10112), .A0(n13553), .A1(n14129), .B0(n13544), .B1(n14130)
         );
  inv01 U3061 ( .Y(n10113), .A(n10112) );
  ao22 U3062 ( .Y(n10114), .A0(n13551), .A1(n14137), .B0(n10195), .B1(n14138)
         );
  inv01 U3063 ( .Y(n10115), .A(n10114) );
  ao22 U3064 ( .Y(n10116), .A0(n14056), .A1(n14085), .B0(n13565), .B1(n10859)
         );
  inv01 U3065 ( .Y(n10117), .A(n10116) );
  ao22 U3066 ( .Y(n10118), .A0(n14056), .A1(n14165), .B0(n13564), .B1(n14166)
         );
  inv01 U3067 ( .Y(n10119), .A(n10118) );
  ao22 U3068 ( .Y(n10120), .A0(n13544), .A1(n14203), .B0(n13545), .B1(n14156)
         );
  inv01 U3069 ( .Y(n10121), .A(n10120) );
  ao22 U3070 ( .Y(n10122), .A0(n13565), .A1(n14117), .B0(n13555), .B1(n14289)
         );
  inv01 U3071 ( .Y(n10123), .A(n10122) );
  ao22 U3072 ( .Y(n10124), .A0(n13565), .A1(n14114), .B0(n13555), .B1(n14277)
         );
  inv01 U3073 ( .Y(n10125), .A(n10124) );
  ao22 U3074 ( .Y(n10126), .A0(n13565), .A1(n14059), .B0(n13539), .B1(n14061)
         );
  inv01 U3075 ( .Y(n10127), .A(n10126) );
  ao22 U3076 ( .Y(n10128), .A0(n10195), .A1(n14194), .B0(n13545), .B1(n14153)
         );
  inv01 U3077 ( .Y(n10129), .A(n10128) );
  ao22 U3078 ( .Y(n10130), .A0(n10195), .A1(n14183), .B0(n13545), .B1(n14144)
         );
  inv01 U3079 ( .Y(n10131), .A(n10130) );
  ao22 U3080 ( .Y(n10132), .A0(n13544), .A1(n14189), .B0(n13545), .B1(n14150)
         );
  inv01 U3081 ( .Y(n10133), .A(n10132) );
  ao22 U3082 ( .Y(n10134), .A0(n14056), .A1(n14077), .B0(n13565), .B1(n14078)
         );
  inv01 U3083 ( .Y(n10135), .A(n10134) );
  ao22 U3084 ( .Y(n10136), .A0(n13565), .A1(n14069), .B0(n13549), .B1(n14070)
         );
  inv01 U3085 ( .Y(n10137), .A(n10136) );
  ao22 U3086 ( .Y(n10138), .A0(n13549), .A1(n14061), .B0(n13564), .B1(n14309)
         );
  inv01 U3087 ( .Y(n10139), .A(n10138) );
  ao22 U3088 ( .Y(n10140), .A0(n13541), .A1(n14073), .B0(n13555), .B1(n14316)
         );
  inv01 U3089 ( .Y(n10141), .A(n10140) );
  ao22 U3090 ( .Y(n10142), .A0(n13553), .A1(n14122), .B0(n10195), .B1(n14150)
         );
  inv01 U3091 ( .Y(n10143), .A(n10142) );
  ao22 U3092 ( .Y(n10144), .A0(n13544), .A1(n14176), .B0(n13535), .B1(n12753)
         );
  inv01 U3093 ( .Y(n10145), .A(n10144) );
  ao22 U3094 ( .Y(n10146), .A0(n13547), .A1(n14065), .B0(n13555), .B1(n14063)
         );
  inv01 U3095 ( .Y(n10147), .A(n10146) );
  ao22 U3096 ( .Y(n10148), .A0(n10195), .A1(n14180), .B0(n13536), .B1(n10275)
         );
  inv01 U3097 ( .Y(n10149), .A(n10148) );
  ao22 U3098 ( .Y(n10150), .A0(n13544), .A1(n14169), .B0(n13536), .B1(n10858)
         );
  inv01 U3099 ( .Y(n10151), .A(n10150) );
  ao22 U3100 ( .Y(n10152), .A0(n10195), .A1(n14173), .B0(n13535), .B1(n10859)
         );
  inv01 U3101 ( .Y(n10153), .A(n10152) );
  ao22 U3102 ( .Y(n10154), .A0(n13551), .A1(n14138), .B0(n10195), .B1(n14156)
         );
  inv01 U3103 ( .Y(n10155), .A(n10154) );
  ao22 U3104 ( .Y(n10156), .A0(n13551), .A1(n14130), .B0(n13544), .B1(n14153)
         );
  inv01 U3105 ( .Y(n10157), .A(n10156) );
  inv01 U3106 ( .Y(n10158), .A(n12438) );
  ao22 U3107 ( .Y(n10159), .A0(n13551), .A1(n14112), .B0(n13544), .B1(n14144)
         );
  inv01 U3108 ( .Y(n10160), .A(n10159) );
  nand02 U3109 ( .Y(n10161), .A0(n12416), .A1(n____return5956_2_) );
  buf04 U3110 ( .Y(n10162), .A(n13591) );
  ao22 U3111 ( .Y(n10163), .A0(n13564), .A1(n14220), .B0(n14056), .B1(n14185)
         );
  inv01 U3112 ( .Y(n10164), .A(n10163) );
  ao22 U3113 ( .Y(n10165), .A0(n12264), .A1(n12828), .B0(n13559), .B1(n14138)
         );
  inv01 U3114 ( .Y(n10166), .A(n10165) );
  ao22 U3115 ( .Y(n10167), .A0(n13564), .A1(n14066), .B0(n14056), .B1(n12809)
         );
  inv01 U3116 ( .Y(n10168), .A(n10167) );
  ao22 U3117 ( .Y(n10169), .A0(n13559), .A1(n14119), .B0(n13545), .B1(n14120)
         );
  inv01 U3118 ( .Y(n10170), .A(n10169) );
  ao22 U3119 ( .Y(n10171), .A0(n13559), .A1(n14127), .B0(n13545), .B1(n14128)
         );
  inv01 U3120 ( .Y(n10172), .A(n10171) );
  ao22 U3121 ( .Y(n10173), .A0(n13559), .A1(n14135), .B0(n13545), .B1(n14136)
         );
  inv01 U3122 ( .Y(n10174), .A(n10173) );
  ao22 U3123 ( .Y(n10175), .A0(n12266), .A1(n14218), .B0(n13554), .B1(n14083)
         );
  inv01 U3124 ( .Y(n10176), .A(n10175) );
  ao22 U3125 ( .Y(n10177), .A0(n13559), .A1(n14129), .B0(n13545), .B1(n14130)
         );
  inv01 U3126 ( .Y(n10178), .A(n10177) );
  ao22 U3127 ( .Y(n10179), .A0(n13559), .A1(n14137), .B0(n13545), .B1(n14138)
         );
  inv01 U3128 ( .Y(n10180), .A(n10179) );
  ao22 U3129 ( .Y(n10181), .A0(n12266), .A1(n14369), .B0(n13564), .B1(n14330)
         );
  inv01 U3130 ( .Y(n10182), .A(n10181) );
  ao22 U3131 ( .Y(n10183), .A0(n12266), .A1(n14159), .B0(n13554), .B1(n14075)
         );
  inv01 U3132 ( .Y(n10184), .A(n10183) );
  ao22 U3133 ( .Y(n10185), .A0(n13565), .A1(n14125), .B0(n13541), .B1(n14052)
         );
  inv01 U3134 ( .Y(n10186), .A(n10185) );
  ao22 U3135 ( .Y(n10187), .A0(n13565), .A1(n14147), .B0(n14056), .B1(n14146)
         );
  inv01 U3136 ( .Y(n10188), .A(n10187) );
  ao22 U3137 ( .Y(n10189), .A0(n12266), .A1(n14307), .B0(n13554), .B1(n14091)
         );
  inv01 U3138 ( .Y(n10190), .A(n10189) );
  ao22 U3139 ( .Y(n10191), .A0(n12927), .A1(n13010), .B0(n13564), .B1(n14205)
         );
  inv01 U3140 ( .Y(n10192), .A(n10191) );
  ao22 U3141 ( .Y(n10193), .A0(n13565), .A1(n14133), .B0(n13547), .B1(n14064)
         );
  inv01 U3142 ( .Y(n10194), .A(n10193) );
  buf08 U3143 ( .Y(n10195), .A(n13543) );
  ao22 U3144 ( .Y(n10196), .A0(n13559), .A1(n14099), .B0(n13545), .B1(n14112)
         );
  inv01 U3145 ( .Y(n10197), .A(n10196) );
  buf02 U3146 ( .Y(n10198), .A(v_count3287_0_) );
  ao21 U3147 ( .Y(n10199), .A0(n13901), .A1(n13902), .B0(n13601) );
  inv01 U3148 ( .Y(n10200), .A(n10199) );
  ao22 U3149 ( .Y(n10201), .A0(n13553), .A1(n14121), .B0(n13544), .B1(n14122)
         );
  inv01 U3150 ( .Y(n10202), .A(n10201) );
  nand02 U3151 ( .Y(n13617), .A0(n10203), .A1(n10204) );
  nand02 U3152 ( .Y(n10203), .A0(n14377), .A1(n14378) );
  inv01 U3153 ( .Y(n10204), .A(s_exp_10b[9]) );
  ao22 U3154 ( .Y(n10205), .A0(n12927), .A1(n14132), .B0(n13564), .B1(n14231)
         );
  inv01 U3155 ( .Y(n10206), .A(n10205) );
  buf02 U3156 ( .Y(n10207), .A(s_frac_rnd7043_12_) );
  buf02 U3157 ( .Y(n10208), .A(s_frac_rnd7043_10_) );
  buf02 U3158 ( .Y(n10209), .A(s_frac_rnd7043_9_) );
  buf02 U3159 ( .Y(n10210), .A(s_frac_rnd7043_19_) );
  buf02 U3160 ( .Y(n10211), .A(s_frac_rnd7043_20_) );
  buf02 U3161 ( .Y(n10212), .A(s_frac_rnd7043_11_) );
  buf02 U3162 ( .Y(n10213), .A(s_frac_rnd7043_3_) );
  buf02 U3163 ( .Y(n10214), .A(s_frac_rnd7043_16_) );
  buf02 U3164 ( .Y(n10215), .A(s_frac_rnd7043_7_) );
  buf02 U3165 ( .Y(n10216), .A(s_frac_rnd7043_21_) );
  buf02 U3166 ( .Y(n10217), .A(s_frac_rnd7043_15_) );
  buf02 U3167 ( .Y(n10218), .A(s_frac_rnd7043_5_) );
  buf02 U3168 ( .Y(n10219), .A(s_frac_rnd7043_17_) );
  buf02 U3169 ( .Y(n10220), .A(s_frac_rnd7043_6_) );
  buf02 U3170 ( .Y(n10221), .A(s_frac_rnd7043_4_) );
  buf02 U3171 ( .Y(n10222), .A(s_frac_rnd7043_13_) );
  buf02 U3172 ( .Y(n10223), .A(s_frac_rnd7043_2_) );
  buf02 U3173 ( .Y(n10224), .A(s_frac_rnd7043_8_) );
  buf02 U3174 ( .Y(n10225), .A(s_frac_rnd7043_14_) );
  buf02 U3175 ( .Y(n10226), .A(s_frac_rnd7043_24_) );
  buf02 U3176 ( .Y(n10227), .A(s_frac_rnd7043_22_) );
  buf02 U3177 ( .Y(n10228), .A(s_frac_rnd7043_18_) );
  buf02 U3178 ( .Y(n10229), .A(s_frac_rnd7043_1_) );
  ao22 U3179 ( .Y(n10230), .A0(n13564), .A1(n14055), .B0(n14056), .B1(n12797)
         );
  inv01 U3180 ( .Y(n10231), .A(n10230) );
  ao22 U3181 ( .Y(n10232), .A0(n13564), .A1(n14094), .B0(n14056), .B1(n14095)
         );
  inv01 U3182 ( .Y(n10233), .A(n10232) );
  ao22 U3183 ( .Y(n10234), .A0(n13564), .A1(n14088), .B0(n14056), .B1(n14089)
         );
  inv01 U3184 ( .Y(n10235), .A(n10234) );
  ao22 U3185 ( .Y(n10236), .A0(n13539), .A1(n14075), .B0(n13564), .B1(n14076)
         );
  inv01 U3186 ( .Y(n10237), .A(n10236) );
  ao22 U3187 ( .Y(n10238), .A0(n13559), .A1(n14120), .B0(n13545), .B1(n14121)
         );
  inv01 U3188 ( .Y(n10239), .A(n10238) );
  ao22 U3189 ( .Y(n10240), .A0(n12927), .A1(n14124), .B0(n13564), .B1(n14336)
         );
  inv01 U3190 ( .Y(n10241), .A(n10240) );
  ao22 U3191 ( .Y(n10242), .A0(n13559), .A1(n14136), .B0(n13545), .B1(n14137)
         );
  inv01 U3192 ( .Y(n10243), .A(n10242) );
  ao22 U3193 ( .Y(n10244), .A0(n13559), .A1(n14128), .B0(n13545), .B1(n14129)
         );
  inv01 U3194 ( .Y(n10245), .A(n10244) );
  ao22 U3195 ( .Y(n10246), .A0(n13539), .A1(n14083), .B0(n13564), .B1(n14084)
         );
  inv01 U3196 ( .Y(n10247), .A(n10246) );
  ao22 U3197 ( .Y(n10248), .A0(n12264), .A1(n14187), .B0(n13559), .B1(n14122)
         );
  inv01 U3198 ( .Y(n10249), .A(n10248) );
  ao22 U3199 ( .Y(n10250), .A0(n13559), .A1(n14103), .B0(n13545), .B1(n14099)
         );
  inv01 U3200 ( .Y(n10251), .A(n10250) );
  ao22 U3201 ( .Y(n10252), .A0(n12264), .A1(n14158), .B0(n13559), .B1(n14112)
         );
  inv01 U3202 ( .Y(n10253), .A(n10252) );
  ao22 U3203 ( .Y(n10254), .A0(n12927), .A1(n14116), .B0(n13564), .B1(n14212)
         );
  inv01 U3204 ( .Y(n10255), .A(n10254) );
  ao22 U3205 ( .Y(n10256), .A0(n12264), .A1(n14193), .B0(n13559), .B1(n14130)
         );
  inv01 U3206 ( .Y(n10257), .A(n10256) );
  or03 U3207 ( .Y(n10258), .A0(n10300), .A1(s_round), .A2(s_frac2a_23_) );
  inv01 U3208 ( .Y(n10259), .A(n10258) );
  nand02 U3209 ( .Y(n14170), .A0(n10260), .A1(n10261) );
  inv01 U3210 ( .Y(n10262), .A(n14122) );
  inv01 U3211 ( .Y(n10263), .A(n14121) );
  inv01 U3212 ( .Y(n10264), .A(n13559) );
  inv01 U3213 ( .Y(n10265), .A(n13545) );
  nand02 U3214 ( .Y(n10266), .A0(n10262), .A1(n10263) );
  nand02 U3215 ( .Y(n10267), .A0(n10262), .A1(n10264) );
  nand02 U3216 ( .Y(n10268), .A0(n10263), .A1(n10265) );
  nand02 U3217 ( .Y(n10269), .A0(n10264), .A1(n10265) );
  nand02 U3218 ( .Y(n10270), .A0(n10266), .A1(n10267) );
  inv01 U3219 ( .Y(n10260), .A(n10270) );
  nand02 U3220 ( .Y(n10271), .A0(n10268), .A1(n10269) );
  inv01 U3221 ( .Y(n10261), .A(n10271) );
  nand03 U3222 ( .Y(n10272), .A0(n13755), .A1(n13756), .A2(s_fract_48_i[14])
         );
  inv02 U3223 ( .Y(n10273), .A(n10272) );
  nand02 U3224 ( .Y(n10274), .A0(n9883), .A1(n14299) );
  inv04 U3225 ( .Y(n10275), .A(n10274) );
  or03 U3226 ( .Y(n10276), .A0(n10389), .A1(n13852), .A2(n13853) );
  inv01 U3227 ( .Y(n10277), .A(n10276) );
  nand03 U3228 ( .Y(n10278), .A0(n12411), .A1(n13927), .A2(n10833) );
  inv02 U3229 ( .Y(n10279), .A(n10278) );
  inv01 U3230 ( .Y(n10281), .A(n10280) );
  ao21 U3231 ( .Y(n10282), .A0(n10506), .A1(n13534), .B0(s_fract_48_i[45]) );
  inv01 U3232 ( .Y(n10283), .A(n10282) );
  or03 U3233 ( .Y(n10284), .A0(n14421), .A1(s_r_zeros_0_), .A2(n14422) );
  inv01 U3234 ( .Y(n10285), .A(n10284) );
  buf02 U3235 ( .Y(n10286), .A(s_fract_48_i[7]) );
  buf02 U3236 ( .Y(n10289), .A(s_fract_48_i[7]) );
  buf02 U3237 ( .Y(n10287), .A(s_fract_48_i[7]) );
  buf02 U3238 ( .Y(n10288), .A(s_fract_48_i[7]) );
  buf02 U3239 ( .Y(n10290), .A(s_fract_48_i[29]) );
  buf02 U3240 ( .Y(n10293), .A(s_fract_48_i[29]) );
  buf02 U3241 ( .Y(n10291), .A(s_fract_48_i[29]) );
  buf02 U3242 ( .Y(n10292), .A(s_fract_48_i[29]) );
  or02 U3243 ( .Y(n10294), .A0(n13582), .A1(n14398) );
  inv01 U3244 ( .Y(n10295), .A(n10294) );
  buf02 U3245 ( .Y(n10296), .A(U1086_U3_Z_0) );
  nor02 U3246 ( .Y(n13618), .A0(n13620), .A1(n10297) );
  nor02 U3247 ( .Y(n10298), .A0(n13621), .A1(n13619) );
  inv01 U3248 ( .Y(n10297), .A(n10298) );
  buf02 U3249 ( .Y(n10299), .A(n13911) );
  buf02 U3250 ( .Y(n10300), .A(n14042) );
  buf02 U3251 ( .Y(n10301), .A(n13845) );
  or03 U3252 ( .Y(n10302), .A0(s_r_zeros_1_), .A1(s_r_zeros_3_), .A2(
        s_r_zeros_2_) );
  inv01 U3253 ( .Y(n10303), .A(n10302) );
  buf02 U3254 ( .Y(n10304), .A(n14011) );
  nand02 U3255 ( .Y(n10305), .A0(n13951), .A1(n13796) );
  inv02 U3256 ( .Y(n10306), .A(n10305) );
  nand02 U3257 ( .Y(v_shl15711_5_), .A0(n10307), .A1(n10308) );
  inv01 U3258 ( .Y(n10309), .A(n13605) );
  inv01 U3259 ( .Y(n10310), .A(n13500) );
  inv01 U3260 ( .Y(n10311), .A(n13603) );
  inv01 U3261 ( .Y(n10312), .A(n13602) );
  nand02 U3262 ( .Y(n10307), .A0(n10309), .A1(n10310) );
  nand02 U3263 ( .Y(n10308), .A0(n10311), .A1(n10312) );
  inv01 U3264 ( .Y(v_shl15711_3_), .A(n10313) );
  nor02 U3265 ( .Y(n10314), .A0(n13500), .A1(n13609) );
  nor02 U3266 ( .Y(n10315), .A0(n13602), .A1(n13608) );
  nor02 U3267 ( .Y(n10313), .A0(n10314), .A1(n10315) );
  inv01 U3268 ( .Y(v_shl15711_2_), .A(n10316) );
  nor02 U3269 ( .Y(n10317), .A0(n13500), .A1(n13611) );
  nor02 U3270 ( .Y(n10318), .A0(n13602), .A1(n13610) );
  nor02 U3271 ( .Y(n10316), .A0(n10317), .A1(n10318) );
  inv02 U3272 ( .Y(n13602), .A(n13966) );
  inv01 U3273 ( .Y(v_shl15711_1_), .A(n10319) );
  nor02 U3274 ( .Y(n10320), .A0(n13500), .A1(n13613) );
  nor02 U3275 ( .Y(n10321), .A0(n13602), .A1(n13612) );
  nor02 U3276 ( .Y(n10319), .A0(n10320), .A1(n10321) );
  buf02 U3277 ( .Y(n13500), .A(n13604) );
  inv01 U3278 ( .Y(v_shl15711_4_), .A(n10322) );
  nor02 U3279 ( .Y(n10323), .A0(n13500), .A1(n13607) );
  nor02 U3280 ( .Y(n10324), .A0(n13602), .A1(n13606) );
  nor02 U3281 ( .Y(n10322), .A0(n10323), .A1(n10324) );
  inv01 U3282 ( .Y(v_shl15711_0_), .A(n10325) );
  nor02 U3283 ( .Y(n10326), .A0(n13500), .A1(n13615) );
  nor02 U3284 ( .Y(n10327), .A0(n13602), .A1(n13614) );
  nor02 U3285 ( .Y(n10325), .A0(n10326), .A1(n10327) );
  or02 U3286 ( .Y(n10328), .A0(n12220), .A1(n14389) );
  inv01 U3287 ( .Y(n10329), .A(n10328) );
  nand03 U3288 ( .Y(n10330), .A0(n13744), .A1(n13745), .A2(n10398) );
  inv02 U3289 ( .Y(n10331), .A(n10330) );
  inv01 U3290 ( .Y(n13675), .A(n10332) );
  inv01 U3291 ( .Y(n10333), .A(n13657) );
  inv01 U3292 ( .Y(n10334), .A(n13656) );
  inv01 U3293 ( .Y(n10335), .A(n13658) );
  nand02 U3294 ( .Y(n10332), .A0(n10335), .A1(n10336) );
  nand02 U3295 ( .Y(n10337), .A0(n10333), .A1(n10334) );
  inv01 U3296 ( .Y(n10336), .A(n10337) );
  buf02 U3297 ( .Y(n10338), .A(n13743) );
  buf02 U3298 ( .Y(n10339), .A(n13743) );
  inv01 U3299 ( .Y(s_output_o_0_), .A(n10340) );
  nor02 U3300 ( .Y(n10341), .A0(n13970), .A1(n14420) );
  nor02 U3301 ( .Y(n10342), .A0(n13972), .A1(n13992) );
  nor02 U3302 ( .Y(n10340), .A0(n10341), .A1(n10342) );
  ao21 U3303 ( .Y(n10343), .A0(n13425), .A1(n13761), .B0(n13716) );
  inv01 U3304 ( .Y(n10344), .A(n10343) );
  inv01 U3305 ( .Y(n13652), .A(n10345) );
  inv01 U3306 ( .Y(n10346), .A(n13660) );
  inv01 U3307 ( .Y(n10347), .A(n13659) );
  inv01 U3308 ( .Y(n10348), .A(n13661) );
  nand02 U3309 ( .Y(n10345), .A0(n10348), .A1(n10349) );
  nand02 U3310 ( .Y(n10350), .A0(n10346), .A1(n10347) );
  inv01 U3311 ( .Y(n10349), .A(n10350) );
  nand02 U3312 ( .Y(n10351), .A0(n13502), .A1(n9632) );
  inv02 U3313 ( .Y(n10352), .A(n10351) );
  or03 U3314 ( .Y(n10353), .A0(n13833), .A1(n13831), .A2(n13832) );
  inv01 U3315 ( .Y(n10354), .A(n10353) );
  or03 U3316 ( .Y(n10355), .A0(n13628), .A1(n13627), .A2(n12470) );
  inv01 U3317 ( .Y(n10356), .A(n10355) );
  nand02 U3318 ( .Y(n13713), .A0(n10357), .A1(n10358) );
  inv01 U3319 ( .Y(n10359), .A(n13716) );
  inv01 U3320 ( .Y(n10360), .A(n13714) );
  inv01 U3321 ( .Y(n10361), .A(n13600) );
  nand02 U3322 ( .Y(n10357), .A0(n10359), .A1(n10360) );
  nand02 U3323 ( .Y(n10358), .A0(n10359), .A1(n10361) );
  nand03 U3324 ( .Y(n10362), .A0(n13750), .A1(n13427), .A2(s_fract_48_i[22])
         );
  inv02 U3325 ( .Y(n10363), .A(n10362) );
  inv04 U3326 ( .Y(n10596), .A(n14074) );
  inv02 U3327 ( .Y(n14074), .A(n13401) );
  or03 U3328 ( .Y(n10364), .A0(n13655), .A1(n13653), .A2(n13654) );
  inv01 U3329 ( .Y(n10365), .A(n10364) );
  nand03 U3330 ( .Y(n10366), .A0(n13916), .A1(n13917), .A2(s_fract_48_i[4]) );
  inv02 U3331 ( .Y(n10367), .A(n10366) );
  buf02 U3332 ( .Y(n10368), .A(n14015) );
  buf02 U3333 ( .Y(n10369), .A(s_fract_48_i[10]) );
  buf02 U3334 ( .Y(n10370), .A(s_fract_48_i[6]) );
  buf02 U3335 ( .Y(n10371), .A(s_fract_48_i[12]) );
  or03 U3336 ( .Y(n10372), .A0(n13839), .A1(n13840), .A2(n10399) );
  inv01 U3337 ( .Y(n10373), .A(n10372) );
  buf02 U3338 ( .Y(n10374), .A(n13918) );
  buf02 U3339 ( .Y(n10375), .A(s_fract_48_i[5]) );
  buf02 U3340 ( .Y(n10378), .A(s_fract_48_i[5]) );
  buf02 U3341 ( .Y(n10376), .A(s_fract_48_i[5]) );
  buf02 U3342 ( .Y(n10377), .A(s_fract_48_i[5]) );
  inv01 U3343 ( .Y(n13694), .A(n10379) );
  inv01 U3344 ( .Y(n10380), .A(n13657) );
  inv01 U3345 ( .Y(n10381), .A(n13656) );
  inv01 U3346 ( .Y(n10382), .A(n13658) );
  nand02 U3347 ( .Y(n10379), .A0(n10382), .A1(n10383) );
  nand02 U3348 ( .Y(n10384), .A0(n10380), .A1(n10381) );
  inv01 U3349 ( .Y(n10383), .A(n10384) );
  or02 U3350 ( .Y(n10385), .A0(n13823), .A1(n13824) );
  inv01 U3351 ( .Y(n10386), .A(n10385) );
  ao21 U3352 ( .Y(n10387), .A0(n13998), .A1(n13997), .B0(n13988) );
  inv01 U3353 ( .Y(n10388), .A(n10387) );
  buf02 U3354 ( .Y(n10389), .A(n13854) );
  buf02 U3355 ( .Y(n10390), .A(n13854) );
  or03 U3356 ( .Y(n10391), .A0(s_opa_i_28_), .A1(s_opa_i_30_), .A2(s_opa_i_29_) );
  inv01 U3357 ( .Y(n10392), .A(n10391) );
  or03 U3358 ( .Y(n10393), .A0(s_opb_i_28_), .A1(s_opb_i_30_), .A2(s_opb_i_29_) );
  inv01 U3359 ( .Y(n10394), .A(n10393) );
  buf02 U3360 ( .Y(n10395), .A(s_fract_48_i[42]) );
  buf02 U3361 ( .Y(n10398), .A(s_fract_48_i[42]) );
  buf02 U3362 ( .Y(n10396), .A(s_fract_48_i[42]) );
  buf02 U3363 ( .Y(n10397), .A(s_fract_48_i[42]) );
  buf02 U3364 ( .Y(n10399), .A(n13856) );
  nand02 U3365 ( .Y(n10400), .A0(n12450), .A1(n____return5956_4_) );
  inv02 U3366 ( .Y(n10401), .A(n10400) );
  xor2 U3367 ( .Y(n10402), .A0(n14398), .A1(n10281) );
  inv01 U3368 ( .Y(n10403), .A(n10402) );
  nand03 U3369 ( .Y(n10404), .A0(n13421), .A1(n13792), .A2(n13771) );
  inv02 U3370 ( .Y(n10405), .A(n10404) );
  inv02 U3371 ( .Y(n10406), .A(s_exp_10a_9_) );
  inv08 U3372 ( .Y(n10407), .A(n10406) );
  or03 U3373 ( .Y(n10408), .A0(n12826), .A1(n10488), .A2(s_expo2b[8]) );
  inv01 U3374 ( .Y(n10409), .A(n10408) );
  inv01 U3375 ( .Y(n14040), .A(n10410) );
  inv01 U3376 ( .Y(n10411), .A(n10259) );
  inv01 U3377 ( .Y(n10412), .A(s_rmode_i_0_) );
  inv01 U3378 ( .Y(n10413), .A(n14043) );
  nand02 U3379 ( .Y(n10410), .A0(n10413), .A1(n10414) );
  nand02 U3380 ( .Y(n10415), .A0(n10411), .A1(n10412) );
  inv01 U3381 ( .Y(n10414), .A(n10415) );
  buf02 U3382 ( .Y(n10416), .A(s_fract_48_i[11]) );
  buf02 U3383 ( .Y(n10419), .A(s_fract_48_i[11]) );
  buf02 U3384 ( .Y(n10417), .A(s_fract_48_i[11]) );
  buf02 U3385 ( .Y(n10418), .A(s_fract_48_i[11]) );
  nand03 U3386 ( .Y(n10420), .A0(n13805), .A1(n13756), .A2(n10474) );
  inv02 U3387 ( .Y(n10421), .A(n10420) );
  nand03 U3388 ( .Y(n10422), .A0(n13752), .A1(n13806), .A2(n13751) );
  inv02 U3389 ( .Y(n10423), .A(n10422) );
  or03 U3390 ( .Y(n10424), .A0(n13982), .A1(n7170_8_), .A2(n13984) );
  inv01 U3391 ( .Y(n10425), .A(n10424) );
  or03 U3392 ( .Y(n10426), .A0(n13844), .A1(n13770), .A2(n13843) );
  inv01 U3393 ( .Y(n10427), .A(n10426) );
  inv01 U3394 ( .Y(n14369), .A(n10428) );
  nor02 U3395 ( .Y(n10429), .A0(n13931), .A1(n13582) );
  nor02 U3396 ( .Y(n10430), .A0(n13810), .A1(n13518) );
  nor02 U3397 ( .Y(n10431), .A0(n14308), .A1(n13598) );
  nor02 U3398 ( .Y(n10428), .A0(n10431), .A1(n10432) );
  nor02 U3399 ( .Y(n10433), .A0(n10429), .A1(n10430) );
  inv01 U3400 ( .Y(n10432), .A(n10433) );
  inv01 U3401 ( .Y(n14307), .A(n10434) );
  nor02 U3402 ( .Y(n10435), .A0(n13811), .A1(n13583) );
  nor02 U3403 ( .Y(n10436), .A0(n14308), .A1(n13518) );
  nor02 U3404 ( .Y(n10437), .A0(n13931), .A1(n13599) );
  nor02 U3405 ( .Y(n10434), .A0(n10437), .A1(n10438) );
  nor02 U3406 ( .Y(n10439), .A0(n10435), .A1(n10436) );
  inv01 U3407 ( .Y(n10438), .A(n10439) );
  inv02 U3408 ( .Y(n13931), .A(s_fract_48_i[3]) );
  buf02 U3409 ( .Y(n13518), .A(n14164) );
  inv01 U3410 ( .Y(n14218), .A(n10440) );
  nor02 U3411 ( .Y(n10441), .A0(n13917), .A1(n13582) );
  nor02 U3412 ( .Y(n10442), .A0(n13931), .A1(n13518) );
  nor02 U3413 ( .Y(n10443), .A0(n13811), .A1(n13598) );
  nor02 U3414 ( .Y(n10440), .A0(n10443), .A1(n10444) );
  nor02 U3415 ( .Y(n10445), .A0(n10441), .A1(n10442) );
  inv01 U3416 ( .Y(n10444), .A(n10445) );
  inv04 U3417 ( .Y(n13753), .A(n10417) );
  nand02 U3418 ( .Y(n14159), .A0(n10446), .A1(n10447) );
  inv01 U3419 ( .Y(n10448), .A(n13583) );
  inv01 U3420 ( .Y(n10449), .A(n13807) );
  inv01 U3421 ( .Y(n10450), .A(n13518) );
  inv01 U3422 ( .Y(n10451), .A(n13811) );
  inv01 U3423 ( .Y(n10452), .A(n13599) );
  inv01 U3424 ( .Y(n10453), .A(n13917) );
  nand02 U3425 ( .Y(n10454), .A0(n10448), .A1(n10449) );
  nand02 U3426 ( .Y(n10455), .A0(n10450), .A1(n10451) );
  nand02 U3427 ( .Y(n10446), .A0(n10452), .A1(n10453) );
  nand02 U3428 ( .Y(n10456), .A0(n10454), .A1(n10455) );
  inv01 U3429 ( .Y(n10447), .A(n10456) );
  inv02 U3430 ( .Y(n13811), .A(s_fract_48_i[4]) );
  nor02 U3431 ( .Y(n13703), .A0(n13641), .A1(n10457) );
  nor02 U3432 ( .Y(n10458), .A0(n13623), .A1(n13624) );
  inv01 U3433 ( .Y(n10457), .A(n10458) );
  or03 U3434 ( .Y(n10459), .A0(n13634), .A1(n13633), .A2(n13207) );
  inv01 U3435 ( .Y(n10460), .A(n10459) );
  inv02 U3436 ( .Y(n13641), .A(n13727) );
  inv01 U3437 ( .Y(n14343), .A(n10461) );
  nor02 U3438 ( .Y(n10462), .A0(n13931), .A1(n13580) );
  nor02 U3439 ( .Y(n10463), .A0(n13811), .A1(n13596) );
  inv01 U3440 ( .Y(n10464), .A(n9885) );
  nor02 U3441 ( .Y(n10461), .A0(n10464), .A1(n10465) );
  nor02 U3442 ( .Y(n10466), .A0(n10462), .A1(n10463) );
  inv01 U3443 ( .Y(n10465), .A(n10466) );
  inv01 U3444 ( .Y(n14339), .A(n10467) );
  nor02 U3445 ( .Y(n10468), .A0(n13746), .A1(n13582) );
  nor02 U3446 ( .Y(n10469), .A0(n13785), .A1(n13598) );
  inv01 U3447 ( .Y(n10470), .A(n9999) );
  nor02 U3448 ( .Y(n10467), .A0(n10470), .A1(n10471) );
  nor02 U3449 ( .Y(n10472), .A0(n10468), .A1(n10469) );
  inv01 U3450 ( .Y(n10471), .A(n10472) );
  buf02 U3451 ( .Y(n10473), .A(n14383) );
  buf02 U3452 ( .Y(n10474), .A(n13940) );
  buf02 U3453 ( .Y(n10475), .A(n13940) );
  nand02 U3454 ( .Y(n10476), .A0(n13780), .A1(n13803) );
  inv02 U3455 ( .Y(n10477), .A(n10476) );
  nand02 U3456 ( .Y(n10478), .A0(n13955), .A1(n13802) );
  inv02 U3457 ( .Y(n10479), .A(n10478) );
  nand02 U3458 ( .Y(n10480), .A0(n13788), .A1(n13797) );
  inv02 U3459 ( .Y(n10481), .A(n10480) );
  inv01 U3460 ( .Y(n14135), .A(n10482) );
  nor02 U3461 ( .Y(n10483), .A0(n13786), .A1(n13580) );
  nor02 U3462 ( .Y(n10484), .A0(n13785), .A1(n13595) );
  inv01 U3463 ( .Y(n10485), .A(n10003) );
  nor02 U3464 ( .Y(n10482), .A0(n10485), .A1(n10486) );
  nor02 U3465 ( .Y(n10487), .A0(n10483), .A1(n10484) );
  inv01 U3466 ( .Y(n10486), .A(n10487) );
  buf02 U3467 ( .Y(n10488), .A(n14012) );
  inv01 U3468 ( .Y(n14119), .A(n10489) );
  nor02 U3469 ( .Y(n10490), .A0(n13746), .A1(n13580) );
  nor02 U3470 ( .Y(n10491), .A0(n13747), .A1(n13595) );
  inv01 U3471 ( .Y(n10492), .A(n9644) );
  nor02 U3472 ( .Y(n10489), .A0(n10492), .A1(n10493) );
  nor02 U3473 ( .Y(n10494), .A0(n10490), .A1(n10491) );
  inv01 U3474 ( .Y(n10493), .A(n10494) );
  inv01 U3475 ( .Y(n14127), .A(n10495) );
  nor02 U3476 ( .Y(n10496), .A0(n13785), .A1(n13580) );
  nor02 U3477 ( .Y(n10497), .A0(n13746), .A1(n13596) );
  inv01 U3478 ( .Y(n10498), .A(n9744) );
  nor02 U3479 ( .Y(n10495), .A0(n10498), .A1(n10499) );
  nor02 U3480 ( .Y(n10500), .A0(n10496), .A1(n10497) );
  inv01 U3481 ( .Y(n10499), .A(n10500) );
  inv02 U3482 ( .Y(s_expo2b[2]), .A(n10488) );
  inv02 U3483 ( .Y(s_expo2b[8]), .A(n9888) );
  buf02 U3484 ( .Y(n10501), .A(s_fract_48_i[13]) );
  buf02 U3485 ( .Y(n10504), .A(s_fract_48_i[13]) );
  buf02 U3486 ( .Y(n10502), .A(s_fract_48_i[13]) );
  buf02 U3487 ( .Y(n10503), .A(s_fract_48_i[13]) );
  buf02 U3488 ( .Y(n13475), .A(s_exp_10a_4_) );
  inv02 U3489 ( .Y(n10505), .A(s_fract_48_i[43]) );
  inv04 U3490 ( .Y(n10506), .A(n10505) );
  buf02 U3491 ( .Y(n10507), .A(n14380) );
  inv01 U3492 ( .Y(n14356), .A(n10508) );
  nor02 U3493 ( .Y(n10509), .A0(n13786), .A1(n13582) );
  nor02 U3494 ( .Y(n10510), .A0(n13745), .A1(n13598) );
  inv01 U3495 ( .Y(n10511), .A(n9945) );
  nor02 U3496 ( .Y(n10508), .A0(n10511), .A1(n10512) );
  nor02 U3497 ( .Y(n10513), .A0(n10509), .A1(n10510) );
  inv01 U3498 ( .Y(n10512), .A(n10513) );
  inv01 U3499 ( .Y(n14348), .A(n10514) );
  nor02 U3500 ( .Y(n10515), .A0(n14308), .A1(n13580) );
  nor02 U3501 ( .Y(n10516), .A0(n13931), .A1(n13595) );
  inv01 U3502 ( .Y(n10517), .A(n9828) );
  nor02 U3503 ( .Y(n10514), .A0(n10517), .A1(n10518) );
  nor02 U3504 ( .Y(n10519), .A0(n10515), .A1(n10516) );
  inv01 U3505 ( .Y(n10518), .A(n10519) );
  inv01 U3506 ( .Y(n14101), .A(n10520) );
  nor02 U3507 ( .Y(n10521), .A0(n13747), .A1(n13580) );
  nor02 U3508 ( .Y(n10522), .A0(n14104), .A1(n13596) );
  inv01 U3509 ( .Y(n10523), .A(n14107) );
  nor02 U3510 ( .Y(n10520), .A0(n10523), .A1(n10524) );
  nor02 U3511 ( .Y(n10525), .A0(n10521), .A1(n10522) );
  inv01 U3512 ( .Y(n10524), .A(n10525) );
  nand02 U3513 ( .Y(n13987), .A0(n10526), .A1(n10527) );
  inv02 U3514 ( .Y(n10528), .A(n13474) );
  inv02 U3515 ( .Y(n10529), .A(n13471) );
  inv02 U3516 ( .Y(n10530), .A(n13989) );
  inv02 U3517 ( .Y(n10531), .A(n13988) );
  inv02 U3518 ( .Y(n10532), .A(s_frac_rnd_22_) );
  inv02 U3519 ( .Y(n10533), .A(s_frac_rnd_23_) );
  nand02 U3520 ( .Y(n10534), .A0(n10530), .A1(n10535) );
  nand02 U3521 ( .Y(n10536), .A0(n10531), .A1(n10537) );
  nand02 U3522 ( .Y(n10538), .A0(n10532), .A1(n10539) );
  nand02 U3523 ( .Y(n10540), .A0(n10532), .A1(n10541) );
  nand02 U3524 ( .Y(n10542), .A0(n10533), .A1(n10543) );
  nand02 U3525 ( .Y(n10544), .A0(n10533), .A1(n10545) );
  nand02 U3526 ( .Y(n10546), .A0(n10533), .A1(n10547) );
  nand02 U3527 ( .Y(n10548), .A0(n10533), .A1(n10549) );
  nand02 U3528 ( .Y(n10550), .A0(n10528), .A1(n10529) );
  inv01 U3529 ( .Y(n10535), .A(n10550) );
  nand02 U3530 ( .Y(n10551), .A0(n10528), .A1(n10529) );
  inv01 U3531 ( .Y(n10537), .A(n10551) );
  nand02 U3532 ( .Y(n10552), .A0(n10528), .A1(n10530) );
  inv01 U3533 ( .Y(n10539), .A(n10552) );
  nand02 U3534 ( .Y(n10553), .A0(n10528), .A1(n10531) );
  inv01 U3535 ( .Y(n10541), .A(n10553) );
  nand02 U3536 ( .Y(n10554), .A0(n10529), .A1(n10530) );
  inv01 U3537 ( .Y(n10543), .A(n10554) );
  nand02 U3538 ( .Y(n10555), .A0(n10529), .A1(n10531) );
  inv01 U3539 ( .Y(n10545), .A(n10555) );
  nand02 U3540 ( .Y(n10556), .A0(n10530), .A1(n10532) );
  inv01 U3541 ( .Y(n10547), .A(n10556) );
  nand02 U3542 ( .Y(n10557), .A0(n10531), .A1(n10532) );
  inv01 U3543 ( .Y(n10549), .A(n10557) );
  nand02 U3544 ( .Y(n10558), .A0(n10534), .A1(n10536) );
  inv01 U3545 ( .Y(n10559), .A(n10558) );
  nand02 U3546 ( .Y(n10560), .A0(n10538), .A1(n10540) );
  inv01 U3547 ( .Y(n10561), .A(n10560) );
  nand02 U3548 ( .Y(n10562), .A0(n10559), .A1(n10561) );
  inv01 U3549 ( .Y(n10526), .A(n10562) );
  nand02 U3550 ( .Y(n10563), .A0(n10542), .A1(n10544) );
  inv01 U3551 ( .Y(n10564), .A(n10563) );
  nand02 U3552 ( .Y(n10565), .A0(n10546), .A1(n10548) );
  inv01 U3553 ( .Y(n10566), .A(n10565) );
  nand02 U3554 ( .Y(n10567), .A0(n10564), .A1(n10566) );
  inv01 U3555 ( .Y(n10527), .A(n10567) );
  buf02 U3556 ( .Y(n10568), .A(s_fract_48_i[16]) );
  buf02 U3557 ( .Y(n10571), .A(s_fract_48_i[16]) );
  buf02 U3558 ( .Y(n10569), .A(s_fract_48_i[16]) );
  buf02 U3559 ( .Y(n10570), .A(s_fract_48_i[16]) );
  buf02 U3560 ( .Y(n10572), .A(s_fract_48_i[27]) );
  buf02 U3561 ( .Y(n10575), .A(s_fract_48_i[27]) );
  buf02 U3562 ( .Y(n10573), .A(s_fract_48_i[27]) );
  buf02 U3563 ( .Y(n10574), .A(s_fract_48_i[27]) );
  inv01 U3564 ( .Y(s_output_o_24_), .A(n10576) );
  nor02 U3565 ( .Y(n10577), .A0(n13982), .A1(n13972) );
  nor02 U3566 ( .Y(n10578), .A0(n13981), .A1(n13970) );
  inv01 U3567 ( .Y(n10579), .A(n13973) );
  nor02 U3568 ( .Y(n10576), .A0(n10579), .A1(n10580) );
  nor02 U3569 ( .Y(n10581), .A0(n10577), .A1(n10578) );
  inv01 U3570 ( .Y(n10580), .A(n10581) );
  inv01 U3571 ( .Y(s_output_o_27_), .A(n10582) );
  nor02 U3572 ( .Y(n10583), .A0(n13979), .A1(n13972) );
  nor02 U3573 ( .Y(n10584), .A0(n13978), .A1(n13970) );
  inv01 U3574 ( .Y(n10585), .A(n13973) );
  nor02 U3575 ( .Y(n10582), .A0(n10585), .A1(n10586) );
  nor02 U3576 ( .Y(n10587), .A0(n10583), .A1(n10584) );
  inv01 U3577 ( .Y(n10586), .A(n10587) );
  inv01 U3578 ( .Y(s_output_o_29_), .A(n10588) );
  nor02 U3579 ( .Y(n10589), .A0(n13975), .A1(n13972) );
  nor02 U3580 ( .Y(n10590), .A0(n13974), .A1(n13970) );
  inv01 U3581 ( .Y(n10591), .A(n13973) );
  nor02 U3582 ( .Y(n10588), .A0(n10591), .A1(n10592) );
  nor02 U3583 ( .Y(n10593), .A0(n10589), .A1(n10590) );
  inv01 U3584 ( .Y(n10592), .A(n10593) );
  inv04 U3585 ( .Y(n13970), .A(n13470) );
  inv04 U3586 ( .Y(n13972), .A(n13473) );
  nand02 U3587 ( .Y(n14350), .A0(n10594), .A1(n10595) );
  inv02 U3588 ( .Y(n10597), .A(n14056) );
  inv02 U3589 ( .Y(n10598), .A(n14072) );
  inv02 U3590 ( .Y(n10599), .A(n13547) );
  inv02 U3591 ( .Y(n10600), .A(n14140) );
  inv02 U3592 ( .Y(n10601), .A(n13554) );
  nand02 U3593 ( .Y(n10602), .A0(n10598), .A1(n10603) );
  nand02 U3594 ( .Y(n10604), .A0(n10599), .A1(n10605) );
  nand02 U3595 ( .Y(n10606), .A0(n10600), .A1(n10607) );
  nand02 U3596 ( .Y(n10608), .A0(n10600), .A1(n10609) );
  nand02 U3597 ( .Y(n10610), .A0(n10601), .A1(n10611) );
  nand02 U3598 ( .Y(n10612), .A0(n10601), .A1(n10613) );
  nand02 U3599 ( .Y(n10614), .A0(n10601), .A1(n10615) );
  nand02 U3600 ( .Y(n10616), .A0(n10601), .A1(n10617) );
  nand02 U3601 ( .Y(n10618), .A0(n10596), .A1(n10597) );
  inv01 U3602 ( .Y(n10603), .A(n10618) );
  nand02 U3603 ( .Y(n10619), .A0(n10596), .A1(n10597) );
  inv01 U3604 ( .Y(n10605), .A(n10619) );
  nand02 U3605 ( .Y(n10620), .A0(n10596), .A1(n10598) );
  inv01 U3606 ( .Y(n10607), .A(n10620) );
  nand02 U3607 ( .Y(n10621), .A0(n10596), .A1(n10599) );
  inv01 U3608 ( .Y(n10609), .A(n10621) );
  nand02 U3609 ( .Y(n10622), .A0(n10597), .A1(n10598) );
  inv01 U3610 ( .Y(n10611), .A(n10622) );
  nand02 U3611 ( .Y(n10623), .A0(n10597), .A1(n10599) );
  inv01 U3612 ( .Y(n10613), .A(n10623) );
  nand02 U3613 ( .Y(n10624), .A0(n10598), .A1(n10600) );
  inv01 U3614 ( .Y(n10615), .A(n10624) );
  nand02 U3615 ( .Y(n10625), .A0(n10599), .A1(n10600) );
  inv01 U3616 ( .Y(n10617), .A(n10625) );
  nand02 U3617 ( .Y(n10626), .A0(n10602), .A1(n10604) );
  inv01 U3618 ( .Y(n10627), .A(n10626) );
  nand02 U3619 ( .Y(n10628), .A0(n10606), .A1(n10608) );
  inv01 U3620 ( .Y(n10629), .A(n10628) );
  nand02 U3621 ( .Y(n10630), .A0(n10627), .A1(n10629) );
  inv01 U3622 ( .Y(n10594), .A(n10630) );
  nand02 U3623 ( .Y(n10631), .A0(n10610), .A1(n10612) );
  inv01 U3624 ( .Y(n10632), .A(n10631) );
  nand02 U3625 ( .Y(n10633), .A0(n10614), .A1(n10616) );
  inv01 U3626 ( .Y(n10634), .A(n10633) );
  nand02 U3627 ( .Y(n10635), .A0(n10632), .A1(n10634) );
  inv01 U3628 ( .Y(n10595), .A(n10635) );
  inv04 U3629 ( .Y(n13547), .A(n13546) );
  inv02 U3630 ( .Y(n14140), .A(n14232) );
  inv04 U3631 ( .Y(n14056), .A(n14346) );
  inv01 U3632 ( .Y(n13695), .A(n10636) );
  inv01 U3633 ( .Y(n10637), .A(n13699) );
  inv01 U3634 ( .Y(n10638), .A(n13698) );
  inv01 U3635 ( .Y(n10639), .A(n13697) );
  inv01 U3636 ( .Y(n10640), .A(n13696) );
  nand02 U3637 ( .Y(n10636), .A0(n10641), .A1(n10642) );
  nand02 U3638 ( .Y(n10643), .A0(n10637), .A1(n10638) );
  inv01 U3639 ( .Y(n10641), .A(n10643) );
  nand02 U3640 ( .Y(n10644), .A0(n10639), .A1(n10640) );
  inv01 U3641 ( .Y(n10642), .A(n10644) );
  or04 U3642 ( .Y(n10645), .A0(n13663), .A1(n13664), .A2(n13665), .A3(n13666)
         );
  inv01 U3643 ( .Y(n10646), .A(n10645) );
  nand02 U3644 ( .Y(n14096), .A0(n10647), .A1(n10648) );
  inv02 U3645 ( .Y(n10649), .A(n14114) );
  inv02 U3646 ( .Y(n10650), .A(n14112) );
  inv02 U3647 ( .Y(n10651), .A(n14110) );
  inv02 U3648 ( .Y(n10652), .A(n13573) );
  inv02 U3649 ( .Y(n10653), .A(n10195) );
  inv02 U3650 ( .Y(n10654), .A(n13536) );
  nand02 U3651 ( .Y(n10655), .A0(n10651), .A1(n10656) );
  nand02 U3652 ( .Y(n10657), .A0(n10652), .A1(n10658) );
  nand02 U3653 ( .Y(n10659), .A0(n10653), .A1(n10660) );
  nand02 U3654 ( .Y(n10661), .A0(n10653), .A1(n10662) );
  nand02 U3655 ( .Y(n10663), .A0(n10654), .A1(n10664) );
  nand02 U3656 ( .Y(n10665), .A0(n10654), .A1(n10666) );
  nand02 U3657 ( .Y(n10667), .A0(n10654), .A1(n10668) );
  nand02 U3658 ( .Y(n10669), .A0(n10654), .A1(n10670) );
  nand02 U3659 ( .Y(n10671), .A0(n10649), .A1(n10650) );
  inv01 U3660 ( .Y(n10656), .A(n10671) );
  nand02 U3661 ( .Y(n10672), .A0(n10649), .A1(n10650) );
  inv01 U3662 ( .Y(n10658), .A(n10672) );
  nand02 U3663 ( .Y(n10673), .A0(n10649), .A1(n10651) );
  inv01 U3664 ( .Y(n10660), .A(n10673) );
  nand02 U3665 ( .Y(n10674), .A0(n10649), .A1(n10652) );
  inv01 U3666 ( .Y(n10662), .A(n10674) );
  nand02 U3667 ( .Y(n10675), .A0(n10650), .A1(n10651) );
  inv01 U3668 ( .Y(n10664), .A(n10675) );
  nand02 U3669 ( .Y(n10676), .A0(n10650), .A1(n10652) );
  inv01 U3670 ( .Y(n10666), .A(n10676) );
  nand02 U3671 ( .Y(n10677), .A0(n10651), .A1(n10653) );
  inv01 U3672 ( .Y(n10668), .A(n10677) );
  nand02 U3673 ( .Y(n10678), .A0(n10652), .A1(n10653) );
  inv01 U3674 ( .Y(n10670), .A(n10678) );
  nand02 U3675 ( .Y(n10679), .A0(n10655), .A1(n10657) );
  inv01 U3676 ( .Y(n10680), .A(n10679) );
  nand02 U3677 ( .Y(n10681), .A0(n10659), .A1(n10661) );
  inv01 U3678 ( .Y(n10682), .A(n10681) );
  nand02 U3679 ( .Y(n10683), .A0(n10680), .A1(n10682) );
  inv01 U3680 ( .Y(n10647), .A(n10683) );
  nand02 U3681 ( .Y(n10684), .A0(n10663), .A1(n10665) );
  inv01 U3682 ( .Y(n10685), .A(n10684) );
  nand02 U3683 ( .Y(n10686), .A0(n10667), .A1(n10669) );
  inv01 U3684 ( .Y(n10687), .A(n10686) );
  nand02 U3685 ( .Y(n10688), .A0(n10685), .A1(n10687) );
  inv01 U3686 ( .Y(n10648), .A(n10688) );
  or04 U3687 ( .Y(n10689), .A0(n14457), .A1(n14458), .A2(n14459), .A3(n14460)
         );
  inv01 U3688 ( .Y(n10690), .A(n10689) );
  or04 U3689 ( .Y(n10691), .A0(n14449), .A1(n14450), .A2(n14451), .A3(n14452)
         );
  inv01 U3690 ( .Y(n10692), .A(n10691) );
  inv02 U3691 ( .Y(n13615), .A(n____return5956_0_) );
  nor02 U3692 ( .Y(n13717), .A0(n10693), .A1(n10694) );
  nor02 U3693 ( .Y(n10695), .A0(n13718), .A1(n13719) );
  inv01 U3694 ( .Y(n10693), .A(n10695) );
  nor02 U3695 ( .Y(n10696), .A0(n13720), .A1(n13721) );
  inv01 U3696 ( .Y(n10694), .A(n10696) );
  nor02 U3697 ( .Y(n13676), .A0(n10697), .A1(n10698) );
  nor02 U3698 ( .Y(n10699), .A0(n13677), .A1(n13678) );
  inv01 U3699 ( .Y(n10697), .A(n10699) );
  nor02 U3700 ( .Y(n10700), .A0(n13679), .A1(n13680) );
  inv01 U3701 ( .Y(n10698), .A(n10700) );
  inv01 U3702 ( .Y(s_output_o_30_), .A(n10701) );
  nor02 U3703 ( .Y(n10702), .A0(n13971), .A1(n13972) );
  nor02 U3704 ( .Y(n10703), .A0(n13969), .A1(n13970) );
  inv01 U3705 ( .Y(n10704), .A(n13973) );
  nor02 U3706 ( .Y(n10701), .A0(n10704), .A1(n10705) );
  nor02 U3707 ( .Y(n10706), .A0(n10702), .A1(n10703) );
  inv01 U3708 ( .Y(n10705), .A(n10706) );
  inv01 U3709 ( .Y(s_output_o_23_), .A(n10707) );
  nor02 U3710 ( .Y(n10708), .A0(n13984), .A1(n13972) );
  nor02 U3711 ( .Y(n10709), .A0(n12826), .A1(n13970) );
  inv01 U3712 ( .Y(n10710), .A(n13973) );
  nor02 U3713 ( .Y(n10707), .A0(n10710), .A1(n10711) );
  nor02 U3714 ( .Y(n10712), .A0(n10708), .A1(n10709) );
  inv01 U3715 ( .Y(n10711), .A(n10712) );
  inv01 U3716 ( .Y(s_output_o_28_), .A(n10713) );
  nor02 U3717 ( .Y(n10714), .A0(n13977), .A1(n13972) );
  nor02 U3718 ( .Y(n10715), .A0(n13976), .A1(n13970) );
  inv01 U3719 ( .Y(n10716), .A(n13973) );
  nor02 U3720 ( .Y(n10713), .A0(n10716), .A1(n10717) );
  nor02 U3721 ( .Y(n10718), .A0(n10714), .A1(n10715) );
  inv01 U3722 ( .Y(n10717), .A(n10718) );
  buf02 U3723 ( .Y(n10719), .A(s_fract_48_i[19]) );
  buf02 U3724 ( .Y(n10722), .A(s_fract_48_i[19]) );
  buf02 U3725 ( .Y(n10720), .A(s_fract_48_i[19]) );
  buf02 U3726 ( .Y(n10721), .A(s_fract_48_i[19]) );
  buf02 U3727 ( .Y(n10723), .A(s_fract_48_i[21]) );
  buf02 U3728 ( .Y(n10726), .A(s_fract_48_i[21]) );
  buf02 U3729 ( .Y(n10724), .A(s_fract_48_i[21]) );
  buf02 U3730 ( .Y(n10725), .A(s_fract_48_i[21]) );
  inv01 U3731 ( .Y(s_frac2a6207_28_), .A(n10727) );
  nor02 U3732 ( .Y(n10728), .A0(n14226), .A1(n13568) );
  nor02 U3733 ( .Y(n10729), .A0(n12833), .A1(n14221) );
  inv01 U3734 ( .Y(n10730), .A(n9881) );
  nor02 U3735 ( .Y(n10727), .A0(n10730), .A1(n10731) );
  nor02 U3736 ( .Y(n10732), .A0(n10728), .A1(n10729) );
  inv01 U3737 ( .Y(n10731), .A(n10732) );
  buf04 U3738 ( .Y(n13568), .A(n14222) );
  inv01 U3739 ( .Y(s_frac2a6207_26_), .A(n10733) );
  nor02 U3740 ( .Y(n10734), .A0(n12914), .A1(n13568) );
  nor02 U3741 ( .Y(n10735), .A0(n12262), .A1(n13563) );
  inv01 U3742 ( .Y(n10736), .A(n9929) );
  nor02 U3743 ( .Y(n10733), .A0(n10736), .A1(n10737) );
  nor02 U3744 ( .Y(n10738), .A0(n10734), .A1(n10735) );
  inv01 U3745 ( .Y(n10737), .A(n10738) );
  inv01 U3746 ( .Y(s_frac2a6207_27_), .A(n10739) );
  nor02 U3747 ( .Y(n10740), .A0(n13563), .A1(n14232) );
  nor02 U3748 ( .Y(n10741), .A0(n12917), .A1(n13568) );
  inv01 U3749 ( .Y(n10742), .A(n9927) );
  nor02 U3750 ( .Y(n10739), .A0(n10742), .A1(n10743) );
  nor02 U3751 ( .Y(n10744), .A0(n10740), .A1(n10741) );
  inv01 U3752 ( .Y(n10743), .A(n10744) );
  nand02 U3753 ( .Y(s_frac2a6207_29_), .A0(n9981), .A1(n10745) );
  inv01 U3754 ( .Y(n10746), .A(n13568) );
  inv01 U3755 ( .Y(n10747), .A(n12891) );
  inv01 U3756 ( .Y(n10748), .A(n14221) );
  inv01 U3757 ( .Y(n10749), .A(n12835) );
  nand02 U3758 ( .Y(n10750), .A0(n10746), .A1(n10747) );
  nand02 U3759 ( .Y(n10751), .A0(n10748), .A1(n10749) );
  nand02 U3760 ( .Y(n10752), .A0(n10750), .A1(n10751) );
  inv01 U3761 ( .Y(n10745), .A(n10752) );
  inv01 U3762 ( .Y(s_frac2a6207_16_), .A(n10753) );
  nor02 U3763 ( .Y(n10754), .A0(n14329), .A1(n13527) );
  nor02 U3764 ( .Y(n10755), .A0(n14255), .A1(n13210) );
  inv01 U3765 ( .Y(n10756), .A(n9826) );
  nor02 U3766 ( .Y(n10753), .A0(n10756), .A1(n10757) );
  nor02 U3767 ( .Y(n10758), .A0(n10754), .A1(n10755) );
  inv01 U3768 ( .Y(n10757), .A(n10758) );
  inv01 U3769 ( .Y(s_frac2a6207_24_), .A(n10759) );
  nor02 U3770 ( .Y(n10760), .A0(n14068), .A1(n13568) );
  nor02 U3771 ( .Y(n10761), .A0(n14252), .A1(n13527) );
  inv01 U3772 ( .Y(n10762), .A(n9773) );
  nor02 U3773 ( .Y(n10759), .A0(n10762), .A1(n10763) );
  nor02 U3774 ( .Y(n10764), .A0(n10760), .A1(n10761) );
  inv01 U3775 ( .Y(n10763), .A(n10764) );
  nand02 U3776 ( .Y(n14097), .A0(n10765), .A1(n10766) );
  inv02 U3777 ( .Y(n10767), .A(n14103) );
  inv02 U3778 ( .Y(n10768), .A(n14101) );
  inv02 U3779 ( .Y(n10769), .A(n14099) );
  inv02 U3780 ( .Y(n10770), .A(n13553) );
  inv02 U3781 ( .Y(n10771), .A(n13559) );
  inv02 U3782 ( .Y(n10772), .A(n13545) );
  nand02 U3783 ( .Y(n10773), .A0(n10769), .A1(n10774) );
  nand02 U3784 ( .Y(n10775), .A0(n10770), .A1(n10776) );
  nand02 U3785 ( .Y(n10777), .A0(n10771), .A1(n10778) );
  nand02 U3786 ( .Y(n10779), .A0(n10771), .A1(n10780) );
  nand02 U3787 ( .Y(n10781), .A0(n10772), .A1(n10782) );
  nand02 U3788 ( .Y(n10783), .A0(n10772), .A1(n10784) );
  nand02 U3789 ( .Y(n10785), .A0(n10772), .A1(n10786) );
  nand02 U3790 ( .Y(n10787), .A0(n10772), .A1(n10788) );
  nand02 U3791 ( .Y(n10789), .A0(n10767), .A1(n10768) );
  inv01 U3792 ( .Y(n10774), .A(n10789) );
  nand02 U3793 ( .Y(n10790), .A0(n10767), .A1(n10768) );
  inv01 U3794 ( .Y(n10776), .A(n10790) );
  nand02 U3795 ( .Y(n10791), .A0(n10767), .A1(n10769) );
  inv01 U3796 ( .Y(n10778), .A(n10791) );
  nand02 U3797 ( .Y(n10792), .A0(n10767), .A1(n10770) );
  inv01 U3798 ( .Y(n10780), .A(n10792) );
  nand02 U3799 ( .Y(n10793), .A0(n10768), .A1(n10769) );
  inv01 U3800 ( .Y(n10782), .A(n10793) );
  nand02 U3801 ( .Y(n10794), .A0(n10768), .A1(n10770) );
  inv01 U3802 ( .Y(n10784), .A(n10794) );
  nand02 U3803 ( .Y(n10795), .A0(n10769), .A1(n10771) );
  inv01 U3804 ( .Y(n10786), .A(n10795) );
  nand02 U3805 ( .Y(n10796), .A0(n10770), .A1(n10771) );
  inv01 U3806 ( .Y(n10788), .A(n10796) );
  nand02 U3807 ( .Y(n10797), .A0(n10773), .A1(n10775) );
  inv01 U3808 ( .Y(n10798), .A(n10797) );
  nand02 U3809 ( .Y(n10799), .A0(n10777), .A1(n10779) );
  inv01 U3810 ( .Y(n10800), .A(n10799) );
  nand02 U3811 ( .Y(n10801), .A0(n10798), .A1(n10800) );
  inv01 U3812 ( .Y(n10765), .A(n10801) );
  nand02 U3813 ( .Y(n10802), .A0(n10781), .A1(n10783) );
  inv01 U3814 ( .Y(n10803), .A(n10802) );
  nand02 U3815 ( .Y(n10804), .A0(n10785), .A1(n10787) );
  inv01 U3816 ( .Y(n10805), .A(n10804) );
  nand02 U3817 ( .Y(n10806), .A0(n10803), .A1(n10805) );
  inv01 U3818 ( .Y(n10766), .A(n10806) );
  buf04 U3819 ( .Y(n13545), .A(n14102) );
  inv01 U3820 ( .Y(s_frac2a6207_19_), .A(n10807) );
  nor02 U3821 ( .Y(n10808), .A0(n14312), .A1(n13563) );
  nor02 U3822 ( .Y(n10809), .A0(n14310), .A1(n13210) );
  inv01 U3823 ( .Y(n10810), .A(n9892) );
  nor02 U3824 ( .Y(n10807), .A0(n10810), .A1(n10811) );
  nor02 U3825 ( .Y(n10812), .A0(n10808), .A1(n10809) );
  inv01 U3826 ( .Y(n10811), .A(n10812) );
  inv01 U3827 ( .Y(s_frac2a6207_17_), .A(n10813) );
  nor02 U3828 ( .Y(n10814), .A0(n14327), .A1(n13527) );
  nor02 U3829 ( .Y(n10815), .A0(n13393), .A1(n13210) );
  inv01 U3830 ( .Y(n10816), .A(n9890) );
  nor02 U3831 ( .Y(n10813), .A0(n10816), .A1(n10817) );
  nor02 U3832 ( .Y(n10818), .A0(n10814), .A1(n10815) );
  inv01 U3833 ( .Y(n10817), .A(n10818) );
  buf04 U3834 ( .Y(n13563), .A(n14230) );
  buf02 U3835 ( .Y(n10819), .A(s_fract_48_i[35]) );
  buf02 U3836 ( .Y(n10822), .A(s_fract_48_i[35]) );
  buf02 U3837 ( .Y(n10820), .A(s_fract_48_i[35]) );
  buf02 U3838 ( .Y(n10821), .A(s_fract_48_i[35]) );
  inv01 U3839 ( .Y(s_frac2a6207_18_), .A(n10823) );
  nor02 U3840 ( .Y(n10824), .A0(n14320), .A1(n14198) );
  nor02 U3841 ( .Y(n10825), .A0(n14319), .A1(n13210) );
  inv01 U3842 ( .Y(n10826), .A(n9894) );
  nor02 U3843 ( .Y(n10823), .A0(n10826), .A1(n10827) );
  nor02 U3844 ( .Y(n10828), .A0(n10824), .A1(n10825) );
  inv01 U3845 ( .Y(n10827), .A(n10828) );
  buf02 U3846 ( .Y(n10829), .A(s_fract_48_i[37]) );
  buf02 U3847 ( .Y(n10832), .A(s_fract_48_i[37]) );
  buf02 U3848 ( .Y(n10830), .A(s_fract_48_i[37]) );
  buf02 U3849 ( .Y(n10831), .A(s_fract_48_i[37]) );
  buf02 U3850 ( .Y(n10833), .A(n13926) );
  or04 U3851 ( .Y(n10834), .A0(n13458), .A1(n13455), .A2(n13461), .A3(n13447)
         );
  inv01 U3852 ( .Y(n10835), .A(n10834) );
  inv01 U3853 ( .Y(n14377), .A(n10836) );
  inv01 U3854 ( .Y(n10837), .A(s_exp_10b[0]) );
  inv01 U3855 ( .Y(n10838), .A(s_exp_10b[1]) );
  inv01 U3856 ( .Y(n10839), .A(s_exp_10b[2]) );
  inv01 U3857 ( .Y(n10840), .A(s_exp_10b[3]) );
  nand02 U3858 ( .Y(n10836), .A0(n10841), .A1(n10842) );
  nand02 U3859 ( .Y(n10843), .A0(n10837), .A1(n10838) );
  inv01 U3860 ( .Y(n10841), .A(n10843) );
  nand02 U3861 ( .Y(n10844), .A0(n10839), .A1(n10840) );
  inv01 U3862 ( .Y(n10842), .A(n10844) );
  or04 U3863 ( .Y(n10845), .A0(n13857), .A1(n13858), .A2(n13859), .A3(n13860)
         );
  inv02 U3864 ( .Y(n10846), .A(n10845) );
  or04 U3865 ( .Y(n10847), .A0(n13812), .A1(n13813), .A2(n13814), .A3(n13815)
         );
  inv02 U3866 ( .Y(n10848), .A(n10847) );
  inv02 U3867 ( .Y(n13885), .A(n10849) );
  inv01 U3868 ( .Y(n10850), .A(n13889) );
  inv01 U3869 ( .Y(n10851), .A(n13888) );
  inv01 U3870 ( .Y(n10852), .A(n13887) );
  inv02 U3871 ( .Y(n10853), .A(n13886) );
  nand02 U3872 ( .Y(n10849), .A0(n10854), .A1(n10855) );
  nand02 U3873 ( .Y(n10856), .A0(n10850), .A1(n10851) );
  inv01 U3874 ( .Y(n10854), .A(n10856) );
  nand02 U3875 ( .Y(n10857), .A0(n10852), .A1(n10853) );
  inv01 U3876 ( .Y(n10855), .A(n10857) );
  ao22 U3877 ( .Y(n10858), .A0(n14269), .A1(n13574), .B0(n14158), .B1(n13566)
         );
  buf02 U3878 ( .Y(n10859), .A(n14086) );
  buf12 U3879 ( .Y(n13574), .A(n14201) );
  or04 U3880 ( .Y(n10860), .A0(n14461), .A1(n14462), .A2(n14463), .A3(n14464)
         );
  inv01 U3881 ( .Y(n10861), .A(n10860) );
  or04 U3882 ( .Y(n10862), .A0(n14453), .A1(n14454), .A2(n14455), .A3(n14456)
         );
  inv01 U3883 ( .Y(n10863), .A(n10862) );
  inv02 U3884 ( .Y(n13903), .A(n10864) );
  inv01 U3885 ( .Y(n10865), .A(n13907) );
  inv01 U3886 ( .Y(n10866), .A(n13906) );
  inv01 U3887 ( .Y(n10867), .A(n13905) );
  inv02 U3888 ( .Y(n10868), .A(n13904) );
  nand02 U3889 ( .Y(n10864), .A0(n10869), .A1(n10870) );
  nand02 U3890 ( .Y(n10871), .A0(n10865), .A1(n10866) );
  inv01 U3891 ( .Y(n10869), .A(n10871) );
  nand02 U3892 ( .Y(n10872), .A0(n10867), .A1(n10868) );
  inv01 U3893 ( .Y(n10870), .A(n10872) );
  inv02 U3894 ( .Y(n13869), .A(n10873) );
  inv01 U3895 ( .Y(n10874), .A(n13873) );
  inv01 U3896 ( .Y(n10875), .A(n13872) );
  inv01 U3897 ( .Y(n10876), .A(n13871) );
  inv02 U3898 ( .Y(n10877), .A(n13870) );
  nand02 U3899 ( .Y(n10873), .A0(n10878), .A1(n10879) );
  nand02 U3900 ( .Y(n10880), .A0(n10874), .A1(n10875) );
  inv01 U3901 ( .Y(n10878), .A(n10880) );
  nand02 U3902 ( .Y(n10881), .A0(n10876), .A1(n10877) );
  inv01 U3903 ( .Y(n10879), .A(n10881) );
  inv02 U3904 ( .Y(n13605), .A(n____return5956_5_) );
  buf02 U3905 ( .Y(n10882), .A(s_fract_48_i[32]) );
  buf02 U3906 ( .Y(n10885), .A(s_fract_48_i[32]) );
  buf02 U3907 ( .Y(n10883), .A(s_fract_48_i[32]) );
  buf02 U3908 ( .Y(n10884), .A(s_fract_48_i[32]) );
  nand02 U3909 ( .Y(n14306), .A0(n10886), .A1(n10887) );
  inv02 U3910 ( .Y(n10888), .A(n14193) );
  inv02 U3911 ( .Y(n10889), .A(n14191) );
  inv02 U3912 ( .Y(n10890), .A(n14052) );
  inv02 U3913 ( .Y(n10891), .A(n13555) );
  inv02 U3914 ( .Y(n10892), .A(n14056) );
  inv02 U3915 ( .Y(n10893), .A(n13559) );
  nand02 U3916 ( .Y(n10894), .A0(n10890), .A1(n10895) );
  nand02 U3917 ( .Y(n10896), .A0(n10891), .A1(n10897) );
  nand02 U3918 ( .Y(n10898), .A0(n10892), .A1(n10899) );
  nand02 U3919 ( .Y(n10900), .A0(n10892), .A1(n10901) );
  nand02 U3920 ( .Y(n10902), .A0(n10893), .A1(n10903) );
  nand02 U3921 ( .Y(n10904), .A0(n10893), .A1(n10905) );
  nand02 U3922 ( .Y(n10906), .A0(n10893), .A1(n10907) );
  nand02 U3923 ( .Y(n10908), .A0(n10893), .A1(n10909) );
  nand02 U3924 ( .Y(n10910), .A0(n10888), .A1(n10889) );
  inv01 U3925 ( .Y(n10895), .A(n10910) );
  nand02 U3926 ( .Y(n10911), .A0(n10888), .A1(n10889) );
  inv01 U3927 ( .Y(n10897), .A(n10911) );
  nand02 U3928 ( .Y(n10912), .A0(n10888), .A1(n10890) );
  inv01 U3929 ( .Y(n10899), .A(n10912) );
  nand02 U3930 ( .Y(n10913), .A0(n10888), .A1(n10891) );
  inv01 U3931 ( .Y(n10901), .A(n10913) );
  nand02 U3932 ( .Y(n10914), .A0(n10889), .A1(n10890) );
  inv01 U3933 ( .Y(n10903), .A(n10914) );
  nand02 U3934 ( .Y(n10915), .A0(n10889), .A1(n10891) );
  inv01 U3935 ( .Y(n10905), .A(n10915) );
  nand02 U3936 ( .Y(n10916), .A0(n10890), .A1(n10892) );
  inv01 U3937 ( .Y(n10907), .A(n10916) );
  nand02 U3938 ( .Y(n10917), .A0(n10891), .A1(n10892) );
  inv01 U3939 ( .Y(n10909), .A(n10917) );
  nand02 U3940 ( .Y(n10918), .A0(n10894), .A1(n10896) );
  inv01 U3941 ( .Y(n10919), .A(n10918) );
  nand02 U3942 ( .Y(n10920), .A0(n10898), .A1(n10900) );
  inv01 U3943 ( .Y(n10921), .A(n10920) );
  nand02 U3944 ( .Y(n10922), .A0(n10919), .A1(n10921) );
  inv01 U3945 ( .Y(n10886), .A(n10922) );
  nand02 U3946 ( .Y(n10923), .A0(n10902), .A1(n10904) );
  inv01 U3947 ( .Y(n10924), .A(n10923) );
  nand02 U3948 ( .Y(n10925), .A0(n10906), .A1(n10908) );
  inv01 U3949 ( .Y(n10926), .A(n10925) );
  nand02 U3950 ( .Y(n10927), .A0(n10924), .A1(n10926) );
  inv01 U3951 ( .Y(n10887), .A(n10927) );
  nand02 U3952 ( .Y(n14071), .A0(n10928), .A1(n10929) );
  inv02 U3953 ( .Y(n10930), .A(n14073) );
  inv02 U3954 ( .Y(n10931), .A(n14072) );
  inv02 U3955 ( .Y(n10932), .A(n13555) );
  inv02 U3956 ( .Y(n10933), .A(n13554) );
  inv02 U3957 ( .Y(n10934), .A(n13548) );
  nand02 U3958 ( .Y(n10935), .A0(n10931), .A1(n10936) );
  nand02 U3959 ( .Y(n10937), .A0(n10932), .A1(n10938) );
  nand02 U3960 ( .Y(n10939), .A0(n10933), .A1(n10940) );
  nand02 U3961 ( .Y(n10941), .A0(n10933), .A1(n10942) );
  nand02 U3962 ( .Y(n10943), .A0(n10934), .A1(n10944) );
  nand02 U3963 ( .Y(n10945), .A0(n10934), .A1(n10946) );
  nand02 U3964 ( .Y(n10947), .A0(n10934), .A1(n10948) );
  nand02 U3965 ( .Y(n10949), .A0(n10934), .A1(n10950) );
  nand02 U3966 ( .Y(n10951), .A0(n10596), .A1(n10930) );
  inv01 U3967 ( .Y(n10936), .A(n10951) );
  nand02 U3968 ( .Y(n10952), .A0(n10596), .A1(n10930) );
  inv01 U3969 ( .Y(n10938), .A(n10952) );
  nand02 U3970 ( .Y(n10953), .A0(n10596), .A1(n10931) );
  inv01 U3971 ( .Y(n10940), .A(n10953) );
  nand02 U3972 ( .Y(n10954), .A0(n10596), .A1(n10932) );
  inv01 U3973 ( .Y(n10942), .A(n10954) );
  nand02 U3974 ( .Y(n10955), .A0(n10930), .A1(n10931) );
  inv01 U3975 ( .Y(n10944), .A(n10955) );
  nand02 U3976 ( .Y(n10956), .A0(n10930), .A1(n10932) );
  inv01 U3977 ( .Y(n10946), .A(n10956) );
  nand02 U3978 ( .Y(n10957), .A0(n10931), .A1(n10933) );
  inv01 U3979 ( .Y(n10948), .A(n10957) );
  nand02 U3980 ( .Y(n10958), .A0(n10932), .A1(n10933) );
  inv01 U3981 ( .Y(n10950), .A(n10958) );
  nand02 U3982 ( .Y(n10959), .A0(n10935), .A1(n10937) );
  inv01 U3983 ( .Y(n10960), .A(n10959) );
  nand02 U3984 ( .Y(n10961), .A0(n10939), .A1(n10941) );
  inv01 U3985 ( .Y(n10962), .A(n10961) );
  nand02 U3986 ( .Y(n10963), .A0(n10960), .A1(n10962) );
  inv01 U3987 ( .Y(n10928), .A(n10963) );
  nand02 U3988 ( .Y(n10964), .A0(n10943), .A1(n10945) );
  inv01 U3989 ( .Y(n10965), .A(n10964) );
  nand02 U3990 ( .Y(n10966), .A0(n10947), .A1(n10949) );
  inv01 U3991 ( .Y(n10967), .A(n10966) );
  nand02 U3992 ( .Y(n10968), .A0(n10965), .A1(n10967) );
  inv01 U3993 ( .Y(n10929), .A(n10968) );
  nand02 U3994 ( .Y(n14334), .A0(n10969), .A1(n10970) );
  inv02 U3995 ( .Y(n10971), .A(n14325) );
  inv02 U3996 ( .Y(n10972), .A(n14081) );
  inv02 U3997 ( .Y(n10973), .A(n14082) );
  inv02 U3998 ( .Y(n10974), .A(n13541) );
  inv02 U3999 ( .Y(n10975), .A(n13554) );
  inv02 U4000 ( .Y(n10976), .A(n13548) );
  nand02 U4001 ( .Y(n10977), .A0(n10973), .A1(n10978) );
  nand02 U4002 ( .Y(n10979), .A0(n10974), .A1(n10980) );
  nand02 U4003 ( .Y(n10981), .A0(n10975), .A1(n10982) );
  nand02 U4004 ( .Y(n10983), .A0(n10975), .A1(n10984) );
  nand02 U4005 ( .Y(n10985), .A0(n10976), .A1(n10986) );
  nand02 U4006 ( .Y(n10987), .A0(n10976), .A1(n10988) );
  nand02 U4007 ( .Y(n10989), .A0(n10976), .A1(n10990) );
  nand02 U4008 ( .Y(n10991), .A0(n10976), .A1(n10992) );
  nand02 U4009 ( .Y(n10993), .A0(n10971), .A1(n10972) );
  inv01 U4010 ( .Y(n10978), .A(n10993) );
  nand02 U4011 ( .Y(n10994), .A0(n10971), .A1(n10972) );
  inv01 U4012 ( .Y(n10980), .A(n10994) );
  nand02 U4013 ( .Y(n10995), .A0(n10971), .A1(n10973) );
  inv01 U4014 ( .Y(n10982), .A(n10995) );
  nand02 U4015 ( .Y(n10996), .A0(n10971), .A1(n10974) );
  inv01 U4016 ( .Y(n10984), .A(n10996) );
  nand02 U4017 ( .Y(n10997), .A0(n10972), .A1(n10973) );
  inv01 U4018 ( .Y(n10986), .A(n10997) );
  nand02 U4019 ( .Y(n10998), .A0(n10972), .A1(n10974) );
  inv01 U4020 ( .Y(n10988), .A(n10998) );
  nand02 U4021 ( .Y(n10999), .A0(n10973), .A1(n10975) );
  inv01 U4022 ( .Y(n10990), .A(n10999) );
  nand02 U4023 ( .Y(n11000), .A0(n10974), .A1(n10975) );
  inv01 U4024 ( .Y(n10992), .A(n11000) );
  nand02 U4025 ( .Y(n11001), .A0(n10977), .A1(n10979) );
  inv01 U4026 ( .Y(n11002), .A(n11001) );
  nand02 U4027 ( .Y(n11003), .A0(n10981), .A1(n10983) );
  inv01 U4028 ( .Y(n11004), .A(n11003) );
  nand02 U4029 ( .Y(n11005), .A0(n11002), .A1(n11004) );
  inv01 U4030 ( .Y(n10969), .A(n11005) );
  nand02 U4031 ( .Y(n11006), .A0(n10985), .A1(n10987) );
  inv01 U4032 ( .Y(n11007), .A(n11006) );
  nand02 U4033 ( .Y(n11008), .A0(n10989), .A1(n10991) );
  inv01 U4034 ( .Y(n11009), .A(n11008) );
  nand02 U4035 ( .Y(n11010), .A0(n11007), .A1(n11009) );
  inv01 U4036 ( .Y(n10970), .A(n11010) );
  nand02 U4037 ( .Y(n14131), .A0(n11011), .A1(n11012) );
  inv02 U4038 ( .Y(n11013), .A(n14134) );
  inv02 U4039 ( .Y(n11014), .A(n14133) );
  inv02 U4040 ( .Y(n11015), .A(n14132) );
  inv02 U4041 ( .Y(n11016), .A(n13541) );
  inv02 U4042 ( .Y(n11017), .A(n13535) );
  inv02 U4043 ( .Y(n11018), .A(n13573) );
  nand02 U4044 ( .Y(n11019), .A0(n11015), .A1(n11020) );
  nand02 U4045 ( .Y(n11021), .A0(n11016), .A1(n11022) );
  nand02 U4046 ( .Y(n11023), .A0(n11017), .A1(n11024) );
  nand02 U4047 ( .Y(n11025), .A0(n11017), .A1(n11026) );
  nand02 U4048 ( .Y(n11027), .A0(n11018), .A1(n11028) );
  nand02 U4049 ( .Y(n11029), .A0(n11018), .A1(n11030) );
  nand02 U4050 ( .Y(n11031), .A0(n11018), .A1(n11032) );
  nand02 U4051 ( .Y(n11033), .A0(n11018), .A1(n11034) );
  nand02 U4052 ( .Y(n11035), .A0(n11013), .A1(n11014) );
  inv01 U4053 ( .Y(n11020), .A(n11035) );
  nand02 U4054 ( .Y(n11036), .A0(n11013), .A1(n11014) );
  inv01 U4055 ( .Y(n11022), .A(n11036) );
  nand02 U4056 ( .Y(n11037), .A0(n11013), .A1(n11015) );
  inv01 U4057 ( .Y(n11024), .A(n11037) );
  nand02 U4058 ( .Y(n11038), .A0(n11013), .A1(n11016) );
  inv01 U4059 ( .Y(n11026), .A(n11038) );
  nand02 U4060 ( .Y(n11039), .A0(n11014), .A1(n11015) );
  inv01 U4061 ( .Y(n11028), .A(n11039) );
  nand02 U4062 ( .Y(n11040), .A0(n11014), .A1(n11016) );
  inv01 U4063 ( .Y(n11030), .A(n11040) );
  nand02 U4064 ( .Y(n11041), .A0(n11015), .A1(n11017) );
  inv01 U4065 ( .Y(n11032), .A(n11041) );
  nand02 U4066 ( .Y(n11042), .A0(n11016), .A1(n11017) );
  inv01 U4067 ( .Y(n11034), .A(n11042) );
  nand02 U4068 ( .Y(n11043), .A0(n11019), .A1(n11021) );
  inv01 U4069 ( .Y(n11044), .A(n11043) );
  nand02 U4070 ( .Y(n11045), .A0(n11023), .A1(n11025) );
  inv01 U4071 ( .Y(n11046), .A(n11045) );
  nand02 U4072 ( .Y(n11047), .A0(n11044), .A1(n11046) );
  inv01 U4073 ( .Y(n11011), .A(n11047) );
  nand02 U4074 ( .Y(n11048), .A0(n11027), .A1(n11029) );
  inv01 U4075 ( .Y(n11049), .A(n11048) );
  nand02 U4076 ( .Y(n11050), .A0(n11031), .A1(n11033) );
  inv01 U4077 ( .Y(n11051), .A(n11050) );
  nand02 U4078 ( .Y(n11052), .A0(n11049), .A1(n11051) );
  inv01 U4079 ( .Y(n11012), .A(n11052) );
  inv02 U4080 ( .Y(n13541), .A(n13538) );
  buf02 U4081 ( .Y(n11053), .A(n14350) );
  nand02 U4082 ( .Y(n14087), .A0(n11054), .A1(n11055) );
  inv02 U4083 ( .Y(n11056), .A(n14052) );
  inv02 U4084 ( .Y(n11057), .A(n14061) );
  inv02 U4085 ( .Y(n11058), .A(n13555) );
  inv02 U4086 ( .Y(n11059), .A(n13554) );
  inv02 U4087 ( .Y(n11060), .A(n13548) );
  nand02 U4088 ( .Y(n11061), .A0(n11180), .A1(n11062) );
  nand02 U4089 ( .Y(n11063), .A0(n11058), .A1(n11064) );
  nand02 U4090 ( .Y(n11065), .A0(n11059), .A1(n11066) );
  nand02 U4091 ( .Y(n11067), .A0(n11059), .A1(n11068) );
  nand02 U4092 ( .Y(n11069), .A0(n11060), .A1(n11070) );
  nand02 U4093 ( .Y(n11071), .A0(n11060), .A1(n11072) );
  nand02 U4094 ( .Y(n11073), .A0(n11060), .A1(n11074) );
  nand02 U4095 ( .Y(n11075), .A0(n11060), .A1(n11076) );
  nand02 U4096 ( .Y(n11077), .A0(n11056), .A1(n11057) );
  inv01 U4097 ( .Y(n11062), .A(n11077) );
  nand02 U4098 ( .Y(n11078), .A0(n11056), .A1(n11057) );
  inv01 U4099 ( .Y(n11064), .A(n11078) );
  nand02 U4100 ( .Y(n11079), .A0(n11056), .A1(n11180) );
  inv01 U4101 ( .Y(n11066), .A(n11079) );
  nand02 U4102 ( .Y(n11080), .A0(n11056), .A1(n11058) );
  inv01 U4103 ( .Y(n11068), .A(n11080) );
  nand02 U4104 ( .Y(n11081), .A0(n11057), .A1(n14328) );
  inv01 U4105 ( .Y(n11070), .A(n11081) );
  nand02 U4106 ( .Y(n11082), .A0(n11057), .A1(n11058) );
  inv01 U4107 ( .Y(n11072), .A(n11082) );
  nand02 U4108 ( .Y(n11083), .A0(n11180), .A1(n11059) );
  inv01 U4109 ( .Y(n11074), .A(n11083) );
  nand02 U4110 ( .Y(n11084), .A0(n11058), .A1(n11059) );
  inv01 U4111 ( .Y(n11076), .A(n11084) );
  nand02 U4112 ( .Y(n11085), .A0(n11061), .A1(n11063) );
  inv01 U4113 ( .Y(n11086), .A(n11085) );
  nand02 U4114 ( .Y(n11087), .A0(n11065), .A1(n11067) );
  inv01 U4115 ( .Y(n11088), .A(n11087) );
  nand02 U4116 ( .Y(n11089), .A0(n11086), .A1(n11088) );
  inv01 U4117 ( .Y(n11054), .A(n11089) );
  nand02 U4118 ( .Y(n11090), .A0(n11069), .A1(n11071) );
  inv01 U4119 ( .Y(n11091), .A(n11090) );
  nand02 U4120 ( .Y(n11092), .A0(n11073), .A1(n11075) );
  inv01 U4121 ( .Y(n11093), .A(n11092) );
  nand02 U4122 ( .Y(n11094), .A0(n11091), .A1(n11093) );
  inv01 U4123 ( .Y(n11055), .A(n11094) );
  nand02 U4124 ( .Y(n14217), .A0(n11095), .A1(n11096) );
  inv02 U4125 ( .Y(n11097), .A(n14080) );
  inv02 U4126 ( .Y(n11098), .A(n14187) );
  inv02 U4127 ( .Y(n11099), .A(n14082) );
  inv02 U4128 ( .Y(n11100), .A(n13555) );
  inv02 U4129 ( .Y(n11101), .A(n13559) );
  inv02 U4130 ( .Y(n11102), .A(n13548) );
  nand02 U4131 ( .Y(n11103), .A0(n11099), .A1(n11104) );
  nand02 U4132 ( .Y(n11105), .A0(n11100), .A1(n11106) );
  nand02 U4133 ( .Y(n11107), .A0(n11101), .A1(n11108) );
  nand02 U4134 ( .Y(n11109), .A0(n11101), .A1(n11110) );
  nand02 U4135 ( .Y(n11111), .A0(n11102), .A1(n11112) );
  nand02 U4136 ( .Y(n11113), .A0(n11102), .A1(n11114) );
  nand02 U4137 ( .Y(n11115), .A0(n11102), .A1(n11116) );
  nand02 U4138 ( .Y(n11117), .A0(n11102), .A1(n11118) );
  nand02 U4139 ( .Y(n11119), .A0(n11097), .A1(n11098) );
  inv01 U4140 ( .Y(n11104), .A(n11119) );
  nand02 U4141 ( .Y(n11120), .A0(n11097), .A1(n11098) );
  inv01 U4142 ( .Y(n11106), .A(n11120) );
  nand02 U4143 ( .Y(n11121), .A0(n11097), .A1(n11099) );
  inv01 U4144 ( .Y(n11108), .A(n11121) );
  nand02 U4145 ( .Y(n11122), .A0(n11097), .A1(n11100) );
  inv01 U4146 ( .Y(n11110), .A(n11122) );
  nand02 U4147 ( .Y(n11123), .A0(n11098), .A1(n11099) );
  inv01 U4148 ( .Y(n11112), .A(n11123) );
  nand02 U4149 ( .Y(n11124), .A0(n11098), .A1(n11100) );
  inv01 U4150 ( .Y(n11114), .A(n11124) );
  nand02 U4151 ( .Y(n11125), .A0(n11099), .A1(n11101) );
  inv01 U4152 ( .Y(n11116), .A(n11125) );
  nand02 U4153 ( .Y(n11126), .A0(n11100), .A1(n11101) );
  inv01 U4154 ( .Y(n11118), .A(n11126) );
  nand02 U4155 ( .Y(n11127), .A0(n11103), .A1(n11105) );
  inv01 U4156 ( .Y(n11128), .A(n11127) );
  nand02 U4157 ( .Y(n11129), .A0(n11107), .A1(n11109) );
  inv01 U4158 ( .Y(n11130), .A(n11129) );
  nand02 U4159 ( .Y(n11131), .A0(n11128), .A1(n11130) );
  inv01 U4160 ( .Y(n11095), .A(n11131) );
  nand02 U4161 ( .Y(n11132), .A0(n11111), .A1(n11113) );
  inv01 U4162 ( .Y(n11133), .A(n11132) );
  nand02 U4163 ( .Y(n11134), .A0(n11115), .A1(n11117) );
  inv01 U4164 ( .Y(n11135), .A(n11134) );
  nand02 U4165 ( .Y(n11136), .A0(n11133), .A1(n11135) );
  inv01 U4166 ( .Y(n11096), .A(n11136) );
  nand02 U4167 ( .Y(n14157), .A0(n11137), .A1(n11138) );
  inv02 U4168 ( .Y(n11139), .A(n14073) );
  inv02 U4169 ( .Y(n11140), .A(n14158) );
  inv02 U4170 ( .Y(n11141), .A(n13555) );
  inv02 U4171 ( .Y(n11142), .A(n13559) );
  inv02 U4172 ( .Y(n11143), .A(n13549) );
  nand02 U4173 ( .Y(n11144), .A0(n10596), .A1(n11145) );
  nand02 U4174 ( .Y(n11146), .A0(n11141), .A1(n11147) );
  nand02 U4175 ( .Y(n11148), .A0(n11142), .A1(n11149) );
  nand02 U4176 ( .Y(n11150), .A0(n11142), .A1(n11151) );
  nand02 U4177 ( .Y(n11152), .A0(n11143), .A1(n11153) );
  nand02 U4178 ( .Y(n11154), .A0(n11143), .A1(n11155) );
  nand02 U4179 ( .Y(n11156), .A0(n11143), .A1(n11157) );
  nand02 U4180 ( .Y(n11158), .A0(n11143), .A1(n11159) );
  nand02 U4181 ( .Y(n11160), .A0(n11139), .A1(n11140) );
  inv01 U4182 ( .Y(n11145), .A(n11160) );
  nand02 U4183 ( .Y(n11161), .A0(n11139), .A1(n11140) );
  inv01 U4184 ( .Y(n11147), .A(n11161) );
  nand02 U4185 ( .Y(n11162), .A0(n11139), .A1(n10596) );
  inv01 U4186 ( .Y(n11149), .A(n11162) );
  nand02 U4187 ( .Y(n11163), .A0(n11139), .A1(n11141) );
  inv01 U4188 ( .Y(n11151), .A(n11163) );
  nand02 U4189 ( .Y(n11164), .A0(n11140), .A1(n10596) );
  inv01 U4190 ( .Y(n11153), .A(n11164) );
  nand02 U4191 ( .Y(n11165), .A0(n11140), .A1(n11141) );
  inv01 U4192 ( .Y(n11155), .A(n11165) );
  nand02 U4193 ( .Y(n11166), .A0(n10596), .A1(n11142) );
  inv01 U4194 ( .Y(n11157), .A(n11166) );
  nand02 U4195 ( .Y(n11167), .A0(n11141), .A1(n11142) );
  inv01 U4196 ( .Y(n11159), .A(n11167) );
  nand02 U4197 ( .Y(n11168), .A0(n11144), .A1(n11146) );
  inv01 U4198 ( .Y(n11169), .A(n11168) );
  nand02 U4199 ( .Y(n11170), .A0(n11148), .A1(n11150) );
  inv01 U4200 ( .Y(n11171), .A(n11170) );
  nand02 U4201 ( .Y(n11172), .A0(n11169), .A1(n11171) );
  inv01 U4202 ( .Y(n11137), .A(n11172) );
  nand02 U4203 ( .Y(n11173), .A0(n11152), .A1(n11154) );
  inv01 U4204 ( .Y(n11174), .A(n11173) );
  nand02 U4205 ( .Y(n11175), .A0(n11156), .A1(n11158) );
  inv01 U4206 ( .Y(n11176), .A(n11175) );
  nand02 U4207 ( .Y(n11177), .A0(n11174), .A1(n11176) );
  inv01 U4208 ( .Y(n11138), .A(n11177) );
  nand02 U4209 ( .Y(n14335), .A0(n11178), .A1(n11179) );
  inv02 U4210 ( .Y(n11180), .A(n14054) );
  inv02 U4211 ( .Y(n11181), .A(n14296) );
  inv02 U4212 ( .Y(n11182), .A(n14050) );
  inv02 U4213 ( .Y(n11183), .A(n13549) );
  inv02 U4214 ( .Y(n11184), .A(n13555) );
  inv02 U4215 ( .Y(n11185), .A(n13554) );
  nand02 U4216 ( .Y(n11186), .A0(n11182), .A1(n11187) );
  nand02 U4217 ( .Y(n11188), .A0(n11183), .A1(n11189) );
  nand02 U4218 ( .Y(n11190), .A0(n11184), .A1(n11191) );
  nand02 U4219 ( .Y(n11192), .A0(n11184), .A1(n11193) );
  nand02 U4220 ( .Y(n11194), .A0(n11185), .A1(n11195) );
  nand02 U4221 ( .Y(n11196), .A0(n11185), .A1(n11197) );
  nand02 U4222 ( .Y(n11198), .A0(n11185), .A1(n11199) );
  nand02 U4223 ( .Y(n11200), .A0(n11185), .A1(n11201) );
  nand02 U4224 ( .Y(n11202), .A0(n11180), .A1(n11181) );
  inv01 U4225 ( .Y(n11187), .A(n11202) );
  nand02 U4226 ( .Y(n11203), .A0(n11180), .A1(n11181) );
  inv01 U4227 ( .Y(n11189), .A(n11203) );
  nand02 U4228 ( .Y(n11204), .A0(n11180), .A1(n11182) );
  inv01 U4229 ( .Y(n11191), .A(n11204) );
  nand02 U4230 ( .Y(n11205), .A0(n11180), .A1(n11183) );
  inv01 U4231 ( .Y(n11193), .A(n11205) );
  nand02 U4232 ( .Y(n11206), .A0(n11181), .A1(n11182) );
  inv01 U4233 ( .Y(n11195), .A(n11206) );
  nand02 U4234 ( .Y(n11207), .A0(n11181), .A1(n11183) );
  inv01 U4235 ( .Y(n11197), .A(n11207) );
  nand02 U4236 ( .Y(n11208), .A0(n11182), .A1(n11184) );
  inv01 U4237 ( .Y(n11199), .A(n11208) );
  nand02 U4238 ( .Y(n11209), .A0(n11183), .A1(n11184) );
  inv01 U4239 ( .Y(n11201), .A(n11209) );
  nand02 U4240 ( .Y(n11210), .A0(n11186), .A1(n11188) );
  inv01 U4241 ( .Y(n11211), .A(n11210) );
  nand02 U4242 ( .Y(n11212), .A0(n11190), .A1(n11192) );
  inv01 U4243 ( .Y(n11213), .A(n11212) );
  nand02 U4244 ( .Y(n11214), .A0(n11211), .A1(n11213) );
  inv01 U4245 ( .Y(n11178), .A(n11214) );
  nand02 U4246 ( .Y(n11215), .A0(n11194), .A1(n11196) );
  inv01 U4247 ( .Y(n11216), .A(n11215) );
  nand02 U4248 ( .Y(n11217), .A0(n11198), .A1(n11200) );
  inv01 U4249 ( .Y(n11218), .A(n11217) );
  nand02 U4250 ( .Y(n11219), .A0(n11216), .A1(n11218) );
  inv01 U4251 ( .Y(n11179), .A(n11219) );
  nand02 U4252 ( .Y(n14062), .A0(n11220), .A1(n11221) );
  inv02 U4253 ( .Y(n11222), .A(n14065) );
  inv02 U4254 ( .Y(n11223), .A(n14064) );
  inv02 U4255 ( .Y(n11224), .A(n14063) );
  inv02 U4256 ( .Y(n11225), .A(n13554) );
  inv02 U4257 ( .Y(n11226), .A(n13555) );
  inv02 U4258 ( .Y(n11227), .A(n13540) );
  nand02 U4259 ( .Y(n11228), .A0(n11224), .A1(n11229) );
  nand02 U4260 ( .Y(n11230), .A0(n11225), .A1(n11231) );
  nand02 U4261 ( .Y(n11232), .A0(n11226), .A1(n11233) );
  nand02 U4262 ( .Y(n11234), .A0(n11226), .A1(n11235) );
  nand02 U4263 ( .Y(n11236), .A0(n11227), .A1(n11237) );
  nand02 U4264 ( .Y(n11238), .A0(n11227), .A1(n11239) );
  nand02 U4265 ( .Y(n11240), .A0(n11227), .A1(n11241) );
  nand02 U4266 ( .Y(n11242), .A0(n11227), .A1(n11243) );
  nand02 U4267 ( .Y(n11244), .A0(n11222), .A1(n11223) );
  inv01 U4268 ( .Y(n11229), .A(n11244) );
  nand02 U4269 ( .Y(n11245), .A0(n11222), .A1(n11223) );
  inv01 U4270 ( .Y(n11231), .A(n11245) );
  nand02 U4271 ( .Y(n11246), .A0(n11222), .A1(n11224) );
  inv01 U4272 ( .Y(n11233), .A(n11246) );
  nand02 U4273 ( .Y(n11247), .A0(n11222), .A1(n11225) );
  inv01 U4274 ( .Y(n11235), .A(n11247) );
  nand02 U4275 ( .Y(n11248), .A0(n11223), .A1(n11224) );
  inv01 U4276 ( .Y(n11237), .A(n11248) );
  nand02 U4277 ( .Y(n11249), .A0(n11223), .A1(n11225) );
  inv01 U4278 ( .Y(n11239), .A(n11249) );
  nand02 U4279 ( .Y(n11250), .A0(n11224), .A1(n11226) );
  inv01 U4280 ( .Y(n11241), .A(n11250) );
  nand02 U4281 ( .Y(n11251), .A0(n11225), .A1(n11226) );
  inv01 U4282 ( .Y(n11243), .A(n11251) );
  nand02 U4283 ( .Y(n11252), .A0(n11228), .A1(n11230) );
  inv01 U4284 ( .Y(n11253), .A(n11252) );
  nand02 U4285 ( .Y(n11254), .A0(n11232), .A1(n11234) );
  inv01 U4286 ( .Y(n11255), .A(n11254) );
  nand02 U4287 ( .Y(n11256), .A0(n11253), .A1(n11255) );
  inv01 U4288 ( .Y(n11220), .A(n11256) );
  nand02 U4289 ( .Y(n11257), .A0(n11236), .A1(n11238) );
  inv01 U4290 ( .Y(n11258), .A(n11257) );
  nand02 U4291 ( .Y(n11259), .A0(n11240), .A1(n11242) );
  inv01 U4292 ( .Y(n11260), .A(n11259) );
  nand02 U4293 ( .Y(n11261), .A0(n11258), .A1(n11260) );
  inv01 U4294 ( .Y(n11221), .A(n11261) );
  inv01 U4295 ( .Y(n14333), .A(n11262) );
  nor02 U4296 ( .Y(n11263), .A0(n14074), .A1(n11264) );
  nor02 U4297 ( .Y(n11265), .A0(n14074), .A1(n11266) );
  nor02 U4298 ( .Y(n11267), .A0(n14074), .A1(n11268) );
  nor02 U4299 ( .Y(n11269), .A0(n14074), .A1(n11270) );
  nor02 U4300 ( .Y(n11271), .A0(n13540), .A1(n11272) );
  nor02 U4301 ( .Y(n11273), .A0(n13540), .A1(n11274) );
  nor02 U4302 ( .Y(n11275), .A0(n13540), .A1(n11276) );
  nor02 U4303 ( .Y(n11277), .A0(n13540), .A1(n11278) );
  nor02 U4304 ( .Y(n11262), .A0(n11279), .A1(n11280) );
  inv01 U4305 ( .Y(n11264), .A(n11284) );
  nor02 U4306 ( .Y(n11281), .A0(n13554), .A1(n14316) );
  inv01 U4307 ( .Y(n11266), .A(n11281) );
  nor02 U4308 ( .Y(n11282), .A0(n14072), .A1(n13548) );
  inv01 U4309 ( .Y(n11268), .A(n11282) );
  nor02 U4310 ( .Y(n11283), .A0(n13554), .A1(n13548) );
  inv01 U4311 ( .Y(n11270), .A(n11283) );
  nor02 U4312 ( .Y(n11284), .A0(n14072), .A1(n14316) );
  inv01 U4313 ( .Y(n11272), .A(n11284) );
  nor02 U4314 ( .Y(n11285), .A0(n13554), .A1(n14316) );
  inv01 U4315 ( .Y(n11274), .A(n11285) );
  nor02 U4316 ( .Y(n11286), .A0(n14072), .A1(n13548) );
  inv01 U4317 ( .Y(n11276), .A(n11286) );
  nor02 U4318 ( .Y(n11287), .A0(n13554), .A1(n13548) );
  inv01 U4319 ( .Y(n11278), .A(n11287) );
  nor02 U4320 ( .Y(n11288), .A0(n11263), .A1(n11265) );
  inv01 U4321 ( .Y(n11289), .A(n11288) );
  nor02 U4322 ( .Y(n11290), .A0(n11267), .A1(n11269) );
  inv01 U4323 ( .Y(n11291), .A(n11290) );
  nor02 U4324 ( .Y(n11292), .A0(n11289), .A1(n11291) );
  inv01 U4325 ( .Y(n11279), .A(n11292) );
  nor02 U4326 ( .Y(n11293), .A0(n11271), .A1(n11273) );
  inv01 U4327 ( .Y(n11294), .A(n11293) );
  nor02 U4328 ( .Y(n11295), .A0(n11275), .A1(n11277) );
  inv01 U4329 ( .Y(n11296), .A(n11295) );
  nor02 U4330 ( .Y(n11297), .A0(n11294), .A1(n11296) );
  inv01 U4331 ( .Y(n11280), .A(n11297) );
  inv01 U4332 ( .Y(n14048), .A(n11298) );
  nor02 U4333 ( .Y(n11299), .A0(n14054), .A1(n11300) );
  nor02 U4334 ( .Y(n11301), .A0(n14054), .A1(n11302) );
  nor02 U4335 ( .Y(n11303), .A0(n14054), .A1(n11304) );
  nor02 U4336 ( .Y(n11305), .A0(n14054), .A1(n11306) );
  nor02 U4337 ( .Y(n11307), .A0(n13547), .A1(n11308) );
  nor02 U4338 ( .Y(n11309), .A0(n13547), .A1(n11310) );
  nor02 U4339 ( .Y(n11311), .A0(n13547), .A1(n11312) );
  nor02 U4340 ( .Y(n11313), .A0(n13547), .A1(n11314) );
  nor02 U4341 ( .Y(n11298), .A0(n11315), .A1(n11316) );
  inv01 U4342 ( .Y(n11300), .A(n11320) );
  nor02 U4343 ( .Y(n11317), .A0(n13555), .A1(n14052) );
  inv01 U4344 ( .Y(n11302), .A(n11317) );
  nor02 U4345 ( .Y(n11318), .A0(n14050), .A1(n13554) );
  inv01 U4346 ( .Y(n11304), .A(n11318) );
  nor02 U4347 ( .Y(n11319), .A0(n13555), .A1(n13554) );
  inv01 U4348 ( .Y(n11306), .A(n11319) );
  nor02 U4349 ( .Y(n11320), .A0(n14050), .A1(n14052) );
  inv01 U4350 ( .Y(n11308), .A(n11320) );
  nor02 U4351 ( .Y(n11321), .A0(n13555), .A1(n14052) );
  inv01 U4352 ( .Y(n11310), .A(n11321) );
  nor02 U4353 ( .Y(n11322), .A0(n14050), .A1(n13554) );
  inv01 U4354 ( .Y(n11312), .A(n11322) );
  nor02 U4355 ( .Y(n11323), .A0(n13555), .A1(n13554) );
  inv01 U4356 ( .Y(n11314), .A(n11323) );
  nor02 U4357 ( .Y(n11324), .A0(n11299), .A1(n11301) );
  inv01 U4358 ( .Y(n11325), .A(n11324) );
  nor02 U4359 ( .Y(n11326), .A0(n11303), .A1(n11305) );
  inv01 U4360 ( .Y(n11327), .A(n11326) );
  nor02 U4361 ( .Y(n11328), .A0(n11325), .A1(n11327) );
  inv01 U4362 ( .Y(n11315), .A(n11328) );
  nor02 U4363 ( .Y(n11329), .A0(n11307), .A1(n11309) );
  inv01 U4364 ( .Y(n11330), .A(n11329) );
  nor02 U4365 ( .Y(n11331), .A0(n11311), .A1(n11313) );
  inv01 U4366 ( .Y(n11332), .A(n11331) );
  nor02 U4367 ( .Y(n11333), .A0(n11330), .A1(n11332) );
  inv01 U4368 ( .Y(n11316), .A(n11333) );
  inv04 U4369 ( .Y(n13548), .A(n13546) );
  nand02 U4370 ( .Y(n14357), .A0(n11334), .A1(n11335) );
  inv02 U4371 ( .Y(n11336), .A(n14080) );
  inv02 U4372 ( .Y(n11337), .A(n14325) );
  inv02 U4373 ( .Y(n11338), .A(n14082) );
  inv02 U4374 ( .Y(n11339), .A(n13554) );
  inv02 U4375 ( .Y(n11340), .A(n13555) );
  inv02 U4376 ( .Y(n11341), .A(n13540) );
  nand02 U4377 ( .Y(n11342), .A0(n11338), .A1(n11343) );
  nand02 U4378 ( .Y(n11344), .A0(n11339), .A1(n11345) );
  nand02 U4379 ( .Y(n11346), .A0(n11340), .A1(n11347) );
  nand02 U4380 ( .Y(n11348), .A0(n11340), .A1(n11349) );
  nand02 U4381 ( .Y(n11350), .A0(n11341), .A1(n11351) );
  nand02 U4382 ( .Y(n11352), .A0(n11341), .A1(n11353) );
  nand02 U4383 ( .Y(n11354), .A0(n11341), .A1(n11355) );
  nand02 U4384 ( .Y(n11356), .A0(n11341), .A1(n11357) );
  nand02 U4385 ( .Y(n11358), .A0(n11336), .A1(n11337) );
  inv01 U4386 ( .Y(n11343), .A(n11358) );
  nand02 U4387 ( .Y(n11359), .A0(n11336), .A1(n11337) );
  inv01 U4388 ( .Y(n11345), .A(n11359) );
  nand02 U4389 ( .Y(n11360), .A0(n11336), .A1(n11338) );
  inv01 U4390 ( .Y(n11347), .A(n11360) );
  nand02 U4391 ( .Y(n11361), .A0(n11336), .A1(n11339) );
  inv01 U4392 ( .Y(n11349), .A(n11361) );
  nand02 U4393 ( .Y(n11362), .A0(n11337), .A1(n11338) );
  inv01 U4394 ( .Y(n11351), .A(n11362) );
  nand02 U4395 ( .Y(n11363), .A0(n11337), .A1(n11339) );
  inv01 U4396 ( .Y(n11353), .A(n11363) );
  nand02 U4397 ( .Y(n11364), .A0(n11338), .A1(n11340) );
  inv01 U4398 ( .Y(n11355), .A(n11364) );
  nand02 U4399 ( .Y(n11365), .A0(n11339), .A1(n11340) );
  inv01 U4400 ( .Y(n11357), .A(n11365) );
  nand02 U4401 ( .Y(n11366), .A0(n11342), .A1(n11344) );
  inv01 U4402 ( .Y(n11367), .A(n11366) );
  nand02 U4403 ( .Y(n11368), .A0(n11346), .A1(n11348) );
  inv01 U4404 ( .Y(n11369), .A(n11368) );
  nand02 U4405 ( .Y(n11370), .A0(n11367), .A1(n11369) );
  inv01 U4406 ( .Y(n11334), .A(n11370) );
  nand02 U4407 ( .Y(n11371), .A0(n11350), .A1(n11352) );
  inv01 U4408 ( .Y(n11372), .A(n11371) );
  nand02 U4409 ( .Y(n11373), .A0(n11354), .A1(n11356) );
  inv01 U4410 ( .Y(n11374), .A(n11373) );
  nand02 U4411 ( .Y(n11375), .A0(n11372), .A1(n11374) );
  inv01 U4412 ( .Y(n11335), .A(n11375) );
  nand02 U4413 ( .Y(n14092), .A0(n11376), .A1(n11377) );
  inv02 U4414 ( .Y(n11378), .A(n14093) );
  inv02 U4415 ( .Y(n11379), .A(n14070) );
  inv02 U4416 ( .Y(n11380), .A(n14065) );
  inv02 U4417 ( .Y(n11381), .A(n13554) );
  inv02 U4418 ( .Y(n11382), .A(n13555) );
  inv02 U4419 ( .Y(n11383), .A(n13540) );
  nand02 U4420 ( .Y(n11384), .A0(n11380), .A1(n11385) );
  nand02 U4421 ( .Y(n11386), .A0(n11381), .A1(n11387) );
  nand02 U4422 ( .Y(n11388), .A0(n11382), .A1(n11389) );
  nand02 U4423 ( .Y(n11390), .A0(n11382), .A1(n11391) );
  nand02 U4424 ( .Y(n11392), .A0(n11383), .A1(n11393) );
  nand02 U4425 ( .Y(n11394), .A0(n11383), .A1(n11395) );
  nand02 U4426 ( .Y(n11396), .A0(n11383), .A1(n11397) );
  nand02 U4427 ( .Y(n11398), .A0(n11383), .A1(n11399) );
  nand02 U4428 ( .Y(n11400), .A0(n11378), .A1(n11379) );
  inv01 U4429 ( .Y(n11385), .A(n11400) );
  nand02 U4430 ( .Y(n11401), .A0(n11378), .A1(n11379) );
  inv01 U4431 ( .Y(n11387), .A(n11401) );
  nand02 U4432 ( .Y(n11402), .A0(n11378), .A1(n11380) );
  inv01 U4433 ( .Y(n11389), .A(n11402) );
  nand02 U4434 ( .Y(n11403), .A0(n11378), .A1(n11381) );
  inv01 U4435 ( .Y(n11391), .A(n11403) );
  nand02 U4436 ( .Y(n11404), .A0(n11379), .A1(n11380) );
  inv01 U4437 ( .Y(n11393), .A(n11404) );
  nand02 U4438 ( .Y(n11405), .A0(n11379), .A1(n11381) );
  inv01 U4439 ( .Y(n11395), .A(n11405) );
  nand02 U4440 ( .Y(n11406), .A0(n11380), .A1(n11382) );
  inv01 U4441 ( .Y(n11397), .A(n11406) );
  nand02 U4442 ( .Y(n11407), .A0(n11381), .A1(n11382) );
  inv01 U4443 ( .Y(n11399), .A(n11407) );
  nand02 U4444 ( .Y(n11408), .A0(n11384), .A1(n11386) );
  inv01 U4445 ( .Y(n11409), .A(n11408) );
  nand02 U4446 ( .Y(n11410), .A0(n11388), .A1(n11390) );
  inv01 U4447 ( .Y(n11411), .A(n11410) );
  nand02 U4448 ( .Y(n11412), .A0(n11409), .A1(n11411) );
  inv01 U4449 ( .Y(n11376), .A(n11412) );
  nand02 U4450 ( .Y(n11413), .A0(n11392), .A1(n11394) );
  inv01 U4451 ( .Y(n11414), .A(n11413) );
  nand02 U4452 ( .Y(n11415), .A0(n11396), .A1(n11398) );
  inv01 U4453 ( .Y(n11416), .A(n11415) );
  nand02 U4454 ( .Y(n11417), .A0(n11414), .A1(n11416) );
  inv01 U4455 ( .Y(n11377), .A(n11417) );
  nand02 U4456 ( .Y(n14079), .A0(n11418), .A1(n11419) );
  inv02 U4457 ( .Y(n11420), .A(n14082) );
  inv02 U4458 ( .Y(n11421), .A(n14081) );
  inv02 U4459 ( .Y(n11422), .A(n14080) );
  inv02 U4460 ( .Y(n11423), .A(n13554) );
  inv02 U4461 ( .Y(n11424), .A(n13555) );
  inv02 U4462 ( .Y(n11425), .A(n13549) );
  nand02 U4463 ( .Y(n11426), .A0(n11422), .A1(n11427) );
  nand02 U4464 ( .Y(n11428), .A0(n11423), .A1(n11429) );
  nand02 U4465 ( .Y(n11430), .A0(n11424), .A1(n11431) );
  nand02 U4466 ( .Y(n11432), .A0(n11424), .A1(n11433) );
  nand02 U4467 ( .Y(n11434), .A0(n11425), .A1(n11435) );
  nand02 U4468 ( .Y(n11436), .A0(n11425), .A1(n11437) );
  nand02 U4469 ( .Y(n11438), .A0(n11425), .A1(n11439) );
  nand02 U4470 ( .Y(n11440), .A0(n11425), .A1(n11441) );
  nand02 U4471 ( .Y(n11442), .A0(n11420), .A1(n11421) );
  inv01 U4472 ( .Y(n11427), .A(n11442) );
  nand02 U4473 ( .Y(n11443), .A0(n11420), .A1(n11421) );
  inv01 U4474 ( .Y(n11429), .A(n11443) );
  nand02 U4475 ( .Y(n11444), .A0(n11420), .A1(n11422) );
  inv01 U4476 ( .Y(n11431), .A(n11444) );
  nand02 U4477 ( .Y(n11445), .A0(n11420), .A1(n11423) );
  inv01 U4478 ( .Y(n11433), .A(n11445) );
  nand02 U4479 ( .Y(n11446), .A0(n11421), .A1(n11422) );
  inv01 U4480 ( .Y(n11435), .A(n11446) );
  nand02 U4481 ( .Y(n11447), .A0(n11421), .A1(n11423) );
  inv01 U4482 ( .Y(n11437), .A(n11447) );
  nand02 U4483 ( .Y(n11448), .A0(n11422), .A1(n11424) );
  inv01 U4484 ( .Y(n11439), .A(n11448) );
  nand02 U4485 ( .Y(n11449), .A0(n11423), .A1(n11424) );
  inv01 U4486 ( .Y(n11441), .A(n11449) );
  nand02 U4487 ( .Y(n11450), .A0(n11426), .A1(n11428) );
  inv01 U4488 ( .Y(n11451), .A(n11450) );
  nand02 U4489 ( .Y(n11452), .A0(n11430), .A1(n11432) );
  inv01 U4490 ( .Y(n11453), .A(n11452) );
  nand02 U4491 ( .Y(n11454), .A0(n11451), .A1(n11453) );
  inv01 U4492 ( .Y(n11418), .A(n11454) );
  nand02 U4493 ( .Y(n11455), .A0(n11434), .A1(n11436) );
  inv01 U4494 ( .Y(n11456), .A(n11455) );
  nand02 U4495 ( .Y(n11457), .A0(n11438), .A1(n11440) );
  inv01 U4496 ( .Y(n11458), .A(n11457) );
  nand02 U4497 ( .Y(n11459), .A0(n11456), .A1(n11458) );
  inv01 U4498 ( .Y(n11419), .A(n11459) );
  inv01 U4499 ( .Y(n14344), .A(n11460) );
  nor02 U4500 ( .Y(n11461), .A0(n14063), .A1(n11462) );
  nor02 U4501 ( .Y(n11463), .A0(n14063), .A1(n11464) );
  nor02 U4502 ( .Y(n11465), .A0(n14063), .A1(n11466) );
  nor02 U4503 ( .Y(n11467), .A0(n14063), .A1(n11468) );
  nor02 U4504 ( .Y(n11469), .A0(n13540), .A1(n11470) );
  nor02 U4505 ( .Y(n11471), .A0(n13540), .A1(n11472) );
  nor02 U4506 ( .Y(n11473), .A0(n13540), .A1(n11474) );
  nor02 U4507 ( .Y(n11475), .A0(n13540), .A1(n11476) );
  nor02 U4508 ( .Y(n11460), .A0(n11477), .A1(n11478) );
  nor02 U4509 ( .Y(n11479), .A0(n14070), .A1(n14259) );
  inv01 U4510 ( .Y(n11462), .A(n11479) );
  nor02 U4511 ( .Y(n11480), .A0(n13554), .A1(n14259) );
  inv01 U4512 ( .Y(n11464), .A(n11480) );
  nor02 U4513 ( .Y(n11481), .A0(n14070), .A1(n13555) );
  inv01 U4514 ( .Y(n11466), .A(n11481) );
  nor02 U4515 ( .Y(n11482), .A0(n13554), .A1(n13555) );
  inv01 U4516 ( .Y(n11468), .A(n11482) );
  nor02 U4517 ( .Y(n11483), .A0(n14070), .A1(n14259) );
  inv01 U4518 ( .Y(n11470), .A(n11483) );
  nor02 U4519 ( .Y(n11484), .A0(n13554), .A1(n14259) );
  inv01 U4520 ( .Y(n11472), .A(n11484) );
  nor02 U4521 ( .Y(n11485), .A0(n14070), .A1(n13555) );
  inv01 U4522 ( .Y(n11474), .A(n11485) );
  nor02 U4523 ( .Y(n11486), .A0(n13554), .A1(n13555) );
  inv01 U4524 ( .Y(n11476), .A(n11486) );
  nor02 U4525 ( .Y(n11487), .A0(n11461), .A1(n11463) );
  inv01 U4526 ( .Y(n11488), .A(n11487) );
  nor02 U4527 ( .Y(n11489), .A0(n11465), .A1(n11467) );
  inv01 U4528 ( .Y(n11490), .A(n11489) );
  nor02 U4529 ( .Y(n11491), .A0(n11488), .A1(n11490) );
  inv01 U4530 ( .Y(n11477), .A(n11491) );
  nor02 U4531 ( .Y(n11492), .A0(n11469), .A1(n11471) );
  inv01 U4532 ( .Y(n11493), .A(n11492) );
  nor02 U4533 ( .Y(n11494), .A0(n11473), .A1(n11475) );
  inv01 U4534 ( .Y(n11495), .A(n11494) );
  nor02 U4535 ( .Y(n11496), .A0(n11493), .A1(n11495) );
  inv01 U4536 ( .Y(n11478), .A(n11496) );
  buf08 U4537 ( .Y(n13555), .A(n14049) );
  inv02 U4538 ( .Y(n13549), .A(n13546) );
  inv04 U4539 ( .Y(n13540), .A(n13538) );
  inv01 U4540 ( .Y(n11497), .A(n14366) );
  nand02 U4541 ( .Y(n14123), .A0(n11498), .A1(n11499) );
  inv02 U4542 ( .Y(n11500), .A(n14126) );
  inv02 U4543 ( .Y(n11501), .A(n14125) );
  inv02 U4544 ( .Y(n11502), .A(n14124) );
  inv02 U4545 ( .Y(n11503), .A(n13539) );
  inv02 U4546 ( .Y(n11504), .A(n13536) );
  inv02 U4547 ( .Y(n11505), .A(n13573) );
  nand02 U4548 ( .Y(n11506), .A0(n11502), .A1(n11507) );
  nand02 U4549 ( .Y(n11508), .A0(n11503), .A1(n11509) );
  nand02 U4550 ( .Y(n11510), .A0(n11504), .A1(n11511) );
  nand02 U4551 ( .Y(n11512), .A0(n11504), .A1(n11513) );
  nand02 U4552 ( .Y(n11514), .A0(n11505), .A1(n11515) );
  nand02 U4553 ( .Y(n11516), .A0(n11505), .A1(n11517) );
  nand02 U4554 ( .Y(n11518), .A0(n11505), .A1(n11519) );
  nand02 U4555 ( .Y(n11520), .A0(n11505), .A1(n11521) );
  nand02 U4556 ( .Y(n11522), .A0(n11500), .A1(n11501) );
  inv01 U4557 ( .Y(n11507), .A(n11522) );
  nand02 U4558 ( .Y(n11523), .A0(n11500), .A1(n11501) );
  inv01 U4559 ( .Y(n11509), .A(n11523) );
  nand02 U4560 ( .Y(n11524), .A0(n11500), .A1(n11502) );
  inv01 U4561 ( .Y(n11511), .A(n11524) );
  nand02 U4562 ( .Y(n11525), .A0(n11500), .A1(n11503) );
  inv01 U4563 ( .Y(n11513), .A(n11525) );
  nand02 U4564 ( .Y(n11526), .A0(n11501), .A1(n11502) );
  inv01 U4565 ( .Y(n11515), .A(n11526) );
  nand02 U4566 ( .Y(n11527), .A0(n11501), .A1(n11503) );
  inv01 U4567 ( .Y(n11517), .A(n11527) );
  nand02 U4568 ( .Y(n11528), .A0(n11502), .A1(n11504) );
  inv01 U4569 ( .Y(n11519), .A(n11528) );
  nand02 U4570 ( .Y(n11529), .A0(n11503), .A1(n11504) );
  inv01 U4571 ( .Y(n11521), .A(n11529) );
  nand02 U4572 ( .Y(n11530), .A0(n11506), .A1(n11508) );
  inv01 U4573 ( .Y(n11531), .A(n11530) );
  nand02 U4574 ( .Y(n11532), .A0(n11510), .A1(n11512) );
  inv01 U4575 ( .Y(n11533), .A(n11532) );
  nand02 U4576 ( .Y(n11534), .A0(n11531), .A1(n11533) );
  inv01 U4577 ( .Y(n11498), .A(n11534) );
  nand02 U4578 ( .Y(n11535), .A0(n11514), .A1(n11516) );
  inv01 U4579 ( .Y(n11536), .A(n11535) );
  nand02 U4580 ( .Y(n11537), .A0(n11518), .A1(n11520) );
  inv01 U4581 ( .Y(n11538), .A(n11537) );
  nand02 U4582 ( .Y(n11539), .A0(n11536), .A1(n11538) );
  inv01 U4583 ( .Y(n11499), .A(n11539) );
  nand02 U4584 ( .Y(n14139), .A0(n11540), .A1(n11541) );
  inv02 U4585 ( .Y(n11542), .A(n14142) );
  inv02 U4586 ( .Y(n11543), .A(n14141) );
  inv02 U4587 ( .Y(n11544), .A(n13569) );
  inv02 U4588 ( .Y(n11545), .A(n14140) );
  inv02 U4589 ( .Y(n11546), .A(n13535) );
  inv02 U4590 ( .Y(n11547), .A(n13573) );
  nand02 U4591 ( .Y(n11548), .A0(n11544), .A1(n11549) );
  nand02 U4592 ( .Y(n11550), .A0(n11545), .A1(n11551) );
  nand02 U4593 ( .Y(n11552), .A0(n11546), .A1(n11553) );
  nand02 U4594 ( .Y(n11554), .A0(n11546), .A1(n11555) );
  nand02 U4595 ( .Y(n11556), .A0(n11547), .A1(n11557) );
  nand02 U4596 ( .Y(n11558), .A0(n11547), .A1(n11559) );
  nand02 U4597 ( .Y(n11560), .A0(n11547), .A1(n11561) );
  nand02 U4598 ( .Y(n11562), .A0(n11547), .A1(n11563) );
  nand02 U4599 ( .Y(n11564), .A0(n11542), .A1(n11543) );
  inv01 U4600 ( .Y(n11549), .A(n11564) );
  nand02 U4601 ( .Y(n11565), .A0(n11542), .A1(n11543) );
  inv01 U4602 ( .Y(n11551), .A(n11565) );
  nand02 U4603 ( .Y(n11566), .A0(n11542), .A1(n11544) );
  inv01 U4604 ( .Y(n11553), .A(n11566) );
  nand02 U4605 ( .Y(n11567), .A0(n11542), .A1(n11545) );
  inv01 U4606 ( .Y(n11555), .A(n11567) );
  nand02 U4607 ( .Y(n11568), .A0(n11543), .A1(n11544) );
  inv01 U4608 ( .Y(n11557), .A(n11568) );
  nand02 U4609 ( .Y(n11569), .A0(n11543), .A1(n11545) );
  inv01 U4610 ( .Y(n11559), .A(n11569) );
  nand02 U4611 ( .Y(n11570), .A0(n11544), .A1(n11546) );
  inv01 U4612 ( .Y(n11561), .A(n11570) );
  nand02 U4613 ( .Y(n11571), .A0(n11545), .A1(n11546) );
  inv01 U4614 ( .Y(n11563), .A(n11571) );
  nand02 U4615 ( .Y(n11572), .A0(n11548), .A1(n11550) );
  inv01 U4616 ( .Y(n11573), .A(n11572) );
  nand02 U4617 ( .Y(n11574), .A0(n11552), .A1(n11554) );
  inv01 U4618 ( .Y(n11575), .A(n11574) );
  nand02 U4619 ( .Y(n11576), .A0(n11573), .A1(n11575) );
  inv01 U4620 ( .Y(n11540), .A(n11576) );
  nand02 U4621 ( .Y(n11577), .A0(n11556), .A1(n11558) );
  inv01 U4622 ( .Y(n11578), .A(n11577) );
  nand02 U4623 ( .Y(n11579), .A0(n11560), .A1(n11562) );
  inv01 U4624 ( .Y(n11580), .A(n11579) );
  nand02 U4625 ( .Y(n11581), .A0(n11578), .A1(n11580) );
  inv01 U4626 ( .Y(n11541), .A(n11581) );
  nand02 U4627 ( .Y(n14115), .A0(n11582), .A1(n11583) );
  inv02 U4628 ( .Y(n11584), .A(n14118) );
  inv02 U4629 ( .Y(n11585), .A(n14117) );
  inv02 U4630 ( .Y(n11586), .A(n14116) );
  inv02 U4631 ( .Y(n11587), .A(n13539) );
  inv02 U4632 ( .Y(n11588), .A(n13573) );
  nand02 U4633 ( .Y(n11589), .A0(n11586), .A1(n11590) );
  nand02 U4634 ( .Y(n11591), .A0(n11587), .A1(n11592) );
  nand02 U4635 ( .Y(n11593), .A0(n11839), .A1(n11594) );
  nand02 U4636 ( .Y(n11595), .A0(n11546), .A1(n11596) );
  nand02 U4637 ( .Y(n11597), .A0(n11588), .A1(n11598) );
  nand02 U4638 ( .Y(n11599), .A0(n11588), .A1(n11600) );
  nand02 U4639 ( .Y(n11601), .A0(n11588), .A1(n11602) );
  nand02 U4640 ( .Y(n11603), .A0(n11588), .A1(n11604) );
  nand02 U4641 ( .Y(n11605), .A0(n11584), .A1(n11585) );
  inv01 U4642 ( .Y(n11590), .A(n11605) );
  nand02 U4643 ( .Y(n11606), .A0(n11584), .A1(n11585) );
  inv01 U4644 ( .Y(n11592), .A(n11606) );
  nand02 U4645 ( .Y(n11607), .A0(n11584), .A1(n11586) );
  inv01 U4646 ( .Y(n11594), .A(n11607) );
  nand02 U4647 ( .Y(n11608), .A0(n11584), .A1(n11587) );
  inv01 U4648 ( .Y(n11596), .A(n11608) );
  nand02 U4649 ( .Y(n11609), .A0(n11585), .A1(n11586) );
  inv01 U4650 ( .Y(n11598), .A(n11609) );
  nand02 U4651 ( .Y(n11610), .A0(n11585), .A1(n11587) );
  inv01 U4652 ( .Y(n11600), .A(n11610) );
  nand02 U4653 ( .Y(n11611), .A0(n11586), .A1(n10654) );
  inv01 U4654 ( .Y(n11602), .A(n11611) );
  nand02 U4655 ( .Y(n11612), .A0(n11587), .A1(n12049) );
  inv01 U4656 ( .Y(n11604), .A(n11612) );
  nand02 U4657 ( .Y(n11613), .A0(n11589), .A1(n11591) );
  inv01 U4658 ( .Y(n11614), .A(n11613) );
  nand02 U4659 ( .Y(n11615), .A0(n11593), .A1(n11595) );
  inv01 U4660 ( .Y(n11616), .A(n11615) );
  nand02 U4661 ( .Y(n11617), .A0(n11614), .A1(n11616) );
  inv01 U4662 ( .Y(n11582), .A(n11617) );
  nand02 U4663 ( .Y(n11618), .A0(n11597), .A1(n11599) );
  inv01 U4664 ( .Y(n11619), .A(n11618) );
  nand02 U4665 ( .Y(n11620), .A0(n11601), .A1(n11603) );
  inv01 U4666 ( .Y(n11621), .A(n11620) );
  nand02 U4667 ( .Y(n11622), .A0(n11619), .A1(n11621) );
  inv01 U4668 ( .Y(n11583), .A(n11622) );
  inv02 U4669 ( .Y(n13611), .A(n____return5956_2_) );
  nand02 U4670 ( .Y(n14364), .A0(n11623), .A1(n11624) );
  inv02 U4671 ( .Y(n11625), .A(n12828) );
  inv02 U4672 ( .Y(n11626), .A(n14093) );
  inv02 U4673 ( .Y(n11627), .A(n14196) );
  inv02 U4674 ( .Y(n11628), .A(n14056) );
  inv02 U4675 ( .Y(n11629), .A(n13554) );
  inv02 U4676 ( .Y(n11630), .A(n13559) );
  nand02 U4677 ( .Y(n11631), .A0(n11627), .A1(n11632) );
  nand02 U4678 ( .Y(n11633), .A0(n11628), .A1(n11634) );
  nand02 U4679 ( .Y(n11635), .A0(n11629), .A1(n11636) );
  nand02 U4680 ( .Y(n11637), .A0(n11629), .A1(n11638) );
  nand02 U4681 ( .Y(n11639), .A0(n11630), .A1(n11640) );
  nand02 U4682 ( .Y(n11641), .A0(n11630), .A1(n11642) );
  nand02 U4683 ( .Y(n11643), .A0(n11630), .A1(n11644) );
  nand02 U4684 ( .Y(n11645), .A0(n11630), .A1(n11646) );
  nand02 U4685 ( .Y(n11647), .A0(n11625), .A1(n11626) );
  inv01 U4686 ( .Y(n11632), .A(n11647) );
  nand02 U4687 ( .Y(n11648), .A0(n11625), .A1(n11626) );
  inv01 U4688 ( .Y(n11634), .A(n11648) );
  nand02 U4689 ( .Y(n11649), .A0(n11625), .A1(n11627) );
  inv01 U4690 ( .Y(n11636), .A(n11649) );
  nand02 U4691 ( .Y(n11650), .A0(n11625), .A1(n11628) );
  inv01 U4692 ( .Y(n11638), .A(n11650) );
  nand02 U4693 ( .Y(n11651), .A0(n11626), .A1(n11627) );
  inv01 U4694 ( .Y(n11640), .A(n11651) );
  nand02 U4695 ( .Y(n11652), .A0(n11626), .A1(n11628) );
  inv01 U4696 ( .Y(n11642), .A(n11652) );
  nand02 U4697 ( .Y(n11653), .A0(n11627), .A1(n11629) );
  inv01 U4698 ( .Y(n11644), .A(n11653) );
  nand02 U4699 ( .Y(n11654), .A0(n11628), .A1(n11629) );
  inv01 U4700 ( .Y(n11646), .A(n11654) );
  nand02 U4701 ( .Y(n11655), .A0(n11631), .A1(n11633) );
  inv01 U4702 ( .Y(n11656), .A(n11655) );
  nand02 U4703 ( .Y(n11657), .A0(n11635), .A1(n11637) );
  inv01 U4704 ( .Y(n11658), .A(n11657) );
  nand02 U4705 ( .Y(n11659), .A0(n11656), .A1(n11658) );
  inv01 U4706 ( .Y(n11623), .A(n11659) );
  nand02 U4707 ( .Y(n11660), .A0(n11639), .A1(n11641) );
  inv01 U4708 ( .Y(n11661), .A(n11660) );
  nand02 U4709 ( .Y(n11662), .A0(n11643), .A1(n11645) );
  inv01 U4710 ( .Y(n11663), .A(n11662) );
  nand02 U4711 ( .Y(n11664), .A0(n11661), .A1(n11663) );
  inv01 U4712 ( .Y(n11624), .A(n11664) );
  buf08 U4713 ( .Y(n13554), .A(n14051) );
  buf08 U4714 ( .Y(n13559), .A(n14100) );
  inv12 U4715 ( .Y(n13573), .A(n13572) );
  nand02 U4716 ( .Y(n14190), .A0(n11665), .A1(n11666) );
  inv02 U4717 ( .Y(n11667), .A(n14192) );
  inv02 U4718 ( .Y(n11668), .A(n14176) );
  inv02 U4719 ( .Y(n11669), .A(n14191) );
  inv02 U4720 ( .Y(n11670), .A(n13569) );
  inv02 U4721 ( .Y(n11671), .A(n13551) );
  inv02 U4722 ( .Y(n11672), .A(n13573) );
  nand02 U4723 ( .Y(n11673), .A0(n11669), .A1(n11674) );
  nand02 U4724 ( .Y(n11675), .A0(n11670), .A1(n11676) );
  nand02 U4725 ( .Y(n11677), .A0(n11671), .A1(n11678) );
  nand02 U4726 ( .Y(n11679), .A0(n11671), .A1(n11680) );
  nand02 U4727 ( .Y(n11681), .A0(n11672), .A1(n11682) );
  nand02 U4728 ( .Y(n11683), .A0(n11672), .A1(n11684) );
  nand02 U4729 ( .Y(n11685), .A0(n11672), .A1(n11686) );
  nand02 U4730 ( .Y(n11687), .A0(n11672), .A1(n11688) );
  nand02 U4731 ( .Y(n11689), .A0(n11667), .A1(n11668) );
  inv01 U4732 ( .Y(n11674), .A(n11689) );
  nand02 U4733 ( .Y(n11690), .A0(n11667), .A1(n11668) );
  inv01 U4734 ( .Y(n11676), .A(n11690) );
  nand02 U4735 ( .Y(n11691), .A0(n11667), .A1(n11669) );
  inv01 U4736 ( .Y(n11678), .A(n11691) );
  nand02 U4737 ( .Y(n11692), .A0(n11667), .A1(n11670) );
  inv01 U4738 ( .Y(n11680), .A(n11692) );
  nand02 U4739 ( .Y(n11693), .A0(n11668), .A1(n11669) );
  inv01 U4740 ( .Y(n11682), .A(n11693) );
  nand02 U4741 ( .Y(n11694), .A0(n11668), .A1(n11670) );
  inv01 U4742 ( .Y(n11684), .A(n11694) );
  nand02 U4743 ( .Y(n11695), .A0(n11669), .A1(n11671) );
  inv01 U4744 ( .Y(n11686), .A(n11695) );
  nand02 U4745 ( .Y(n11696), .A0(n11670), .A1(n11671) );
  inv01 U4746 ( .Y(n11688), .A(n11696) );
  nand02 U4747 ( .Y(n11697), .A0(n11673), .A1(n11675) );
  inv01 U4748 ( .Y(n11698), .A(n11697) );
  nand02 U4749 ( .Y(n11699), .A0(n11677), .A1(n11679) );
  inv01 U4750 ( .Y(n11700), .A(n11699) );
  nand02 U4751 ( .Y(n11701), .A0(n11698), .A1(n11700) );
  inv01 U4752 ( .Y(n11665), .A(n11701) );
  nand02 U4753 ( .Y(n11702), .A0(n11681), .A1(n11683) );
  inv01 U4754 ( .Y(n11703), .A(n11702) );
  nand02 U4755 ( .Y(n11704), .A0(n11685), .A1(n11687) );
  inv01 U4756 ( .Y(n11705), .A(n11704) );
  nand02 U4757 ( .Y(n11706), .A0(n11703), .A1(n11705) );
  inv01 U4758 ( .Y(n11666), .A(n11706) );
  nand02 U4759 ( .Y(n14154), .A0(n11707), .A1(n11708) );
  inv02 U4760 ( .Y(n11709), .A(n14155) );
  inv02 U4761 ( .Y(n11710), .A(n14069) );
  inv02 U4762 ( .Y(n11711), .A(n12809) );
  inv02 U4763 ( .Y(n11712), .A(n13569) );
  inv02 U4764 ( .Y(n11713), .A(n13535) );
  inv02 U4765 ( .Y(n11714), .A(n13573) );
  nand02 U4766 ( .Y(n11715), .A0(n11711), .A1(n11716) );
  nand02 U4767 ( .Y(n11717), .A0(n11712), .A1(n11718) );
  nand02 U4768 ( .Y(n11719), .A0(n11713), .A1(n11720) );
  nand02 U4769 ( .Y(n11721), .A0(n11713), .A1(n11722) );
  nand02 U4770 ( .Y(n11723), .A0(n11714), .A1(n11724) );
  nand02 U4771 ( .Y(n11725), .A0(n11714), .A1(n11726) );
  nand02 U4772 ( .Y(n11727), .A0(n11714), .A1(n11728) );
  nand02 U4773 ( .Y(n11729), .A0(n11714), .A1(n11730) );
  nand02 U4774 ( .Y(n11731), .A0(n11709), .A1(n11710) );
  inv01 U4775 ( .Y(n11716), .A(n11731) );
  nand02 U4776 ( .Y(n11732), .A0(n11709), .A1(n11710) );
  inv01 U4777 ( .Y(n11718), .A(n11732) );
  nand02 U4778 ( .Y(n11733), .A0(n11709), .A1(n11711) );
  inv01 U4779 ( .Y(n11720), .A(n11733) );
  nand02 U4780 ( .Y(n11734), .A0(n11709), .A1(n11712) );
  inv01 U4781 ( .Y(n11722), .A(n11734) );
  nand02 U4782 ( .Y(n11735), .A0(n11710), .A1(n11711) );
  inv01 U4783 ( .Y(n11724), .A(n11735) );
  nand02 U4784 ( .Y(n11736), .A0(n11710), .A1(n11712) );
  inv01 U4785 ( .Y(n11726), .A(n11736) );
  nand02 U4786 ( .Y(n11737), .A0(n11711), .A1(n11713) );
  inv01 U4787 ( .Y(n11728), .A(n11737) );
  nand02 U4788 ( .Y(n11738), .A0(n11712), .A1(n11713) );
  inv01 U4789 ( .Y(n11730), .A(n11738) );
  nand02 U4790 ( .Y(n11739), .A0(n11715), .A1(n11717) );
  inv01 U4791 ( .Y(n11740), .A(n11739) );
  nand02 U4792 ( .Y(n11741), .A0(n11719), .A1(n11721) );
  inv01 U4793 ( .Y(n11742), .A(n11741) );
  nand02 U4794 ( .Y(n11743), .A0(n11740), .A1(n11742) );
  inv01 U4795 ( .Y(n11707), .A(n11743) );
  nand02 U4796 ( .Y(n11744), .A0(n11723), .A1(n11725) );
  inv01 U4797 ( .Y(n11745), .A(n11744) );
  nand02 U4798 ( .Y(n11746), .A0(n11727), .A1(n11729) );
  inv01 U4799 ( .Y(n11747), .A(n11746) );
  nand02 U4800 ( .Y(n11748), .A0(n11745), .A1(n11747) );
  inv01 U4801 ( .Y(n11708), .A(n11748) );
  inv04 U4802 ( .Y(n13551), .A(n13550) );
  buf04 U4803 ( .Y(n13535), .A(n14113) );
  nand02 U4804 ( .Y(n14171), .A0(n11749), .A1(n11750) );
  inv02 U4805 ( .Y(n11751), .A(n14172) );
  inv02 U4806 ( .Y(n11752), .A(n14150) );
  inv02 U4807 ( .Y(n11753), .A(n14085) );
  inv02 U4808 ( .Y(n11754), .A(n13569) );
  inv02 U4809 ( .Y(n11755), .A(n13552) );
  inv02 U4810 ( .Y(n11756), .A(n13573) );
  nand02 U4811 ( .Y(n11757), .A0(n11753), .A1(n11758) );
  nand02 U4812 ( .Y(n11759), .A0(n11754), .A1(n11760) );
  nand02 U4813 ( .Y(n11761), .A0(n11755), .A1(n11762) );
  nand02 U4814 ( .Y(n11763), .A0(n11755), .A1(n11764) );
  nand02 U4815 ( .Y(n11765), .A0(n11756), .A1(n11766) );
  nand02 U4816 ( .Y(n11767), .A0(n11756), .A1(n11768) );
  nand02 U4817 ( .Y(n11769), .A0(n11756), .A1(n11770) );
  nand02 U4818 ( .Y(n11771), .A0(n11756), .A1(n11772) );
  nand02 U4819 ( .Y(n11773), .A0(n11751), .A1(n11752) );
  inv01 U4820 ( .Y(n11758), .A(n11773) );
  nand02 U4821 ( .Y(n11774), .A0(n11751), .A1(n11752) );
  inv01 U4822 ( .Y(n11760), .A(n11774) );
  nand02 U4823 ( .Y(n11775), .A0(n11751), .A1(n11753) );
  inv01 U4824 ( .Y(n11762), .A(n11775) );
  nand02 U4825 ( .Y(n11776), .A0(n11751), .A1(n11754) );
  inv01 U4826 ( .Y(n11764), .A(n11776) );
  nand02 U4827 ( .Y(n11777), .A0(n11752), .A1(n11753) );
  inv01 U4828 ( .Y(n11766), .A(n11777) );
  nand02 U4829 ( .Y(n11778), .A0(n11752), .A1(n11754) );
  inv01 U4830 ( .Y(n11768), .A(n11778) );
  nand02 U4831 ( .Y(n11779), .A0(n11753), .A1(n11755) );
  inv01 U4832 ( .Y(n11770), .A(n11779) );
  nand02 U4833 ( .Y(n11780), .A0(n11754), .A1(n11755) );
  inv01 U4834 ( .Y(n11772), .A(n11780) );
  nand02 U4835 ( .Y(n11781), .A0(n11757), .A1(n11759) );
  inv01 U4836 ( .Y(n11782), .A(n11781) );
  nand02 U4837 ( .Y(n11783), .A0(n11761), .A1(n11763) );
  inv01 U4838 ( .Y(n11784), .A(n11783) );
  nand02 U4839 ( .Y(n11785), .A0(n11782), .A1(n11784) );
  inv01 U4840 ( .Y(n11749), .A(n11785) );
  nand02 U4841 ( .Y(n11786), .A0(n11765), .A1(n11767) );
  inv01 U4842 ( .Y(n11787), .A(n11786) );
  nand02 U4843 ( .Y(n11788), .A0(n11769), .A1(n11771) );
  inv01 U4844 ( .Y(n11789), .A(n11788) );
  nand02 U4845 ( .Y(n11790), .A0(n11787), .A1(n11789) );
  inv01 U4846 ( .Y(n11750), .A(n11790) );
  nand02 U4847 ( .Y(n14174), .A0(n11791), .A1(n11792) );
  inv02 U4848 ( .Y(n11793), .A(n14175) );
  inv02 U4849 ( .Y(n11794), .A(n14153) );
  inv02 U4850 ( .Y(n11795), .A(n14089) );
  inv02 U4851 ( .Y(n11796), .A(n13569) );
  inv02 U4852 ( .Y(n11797), .A(n13552) );
  inv02 U4853 ( .Y(n11798), .A(n13573) );
  nand02 U4854 ( .Y(n11799), .A0(n11795), .A1(n11800) );
  nand02 U4855 ( .Y(n11801), .A0(n11796), .A1(n11802) );
  nand02 U4856 ( .Y(n11803), .A0(n11797), .A1(n11804) );
  nand02 U4857 ( .Y(n11805), .A0(n11797), .A1(n11806) );
  nand02 U4858 ( .Y(n11807), .A0(n11798), .A1(n11808) );
  nand02 U4859 ( .Y(n11809), .A0(n11798), .A1(n11810) );
  nand02 U4860 ( .Y(n11811), .A0(n11798), .A1(n11812) );
  nand02 U4861 ( .Y(n11813), .A0(n11798), .A1(n11814) );
  nand02 U4862 ( .Y(n11815), .A0(n11793), .A1(n11794) );
  inv01 U4863 ( .Y(n11800), .A(n11815) );
  nand02 U4864 ( .Y(n11816), .A0(n11793), .A1(n11794) );
  inv01 U4865 ( .Y(n11802), .A(n11816) );
  nand02 U4866 ( .Y(n11817), .A0(n11793), .A1(n11795) );
  inv01 U4867 ( .Y(n11804), .A(n11817) );
  nand02 U4868 ( .Y(n11818), .A0(n11793), .A1(n11796) );
  inv01 U4869 ( .Y(n11806), .A(n11818) );
  nand02 U4870 ( .Y(n11819), .A0(n11794), .A1(n11795) );
  inv01 U4871 ( .Y(n11808), .A(n11819) );
  nand02 U4872 ( .Y(n11820), .A0(n11794), .A1(n11796) );
  inv01 U4873 ( .Y(n11810), .A(n11820) );
  nand02 U4874 ( .Y(n11821), .A0(n11795), .A1(n11797) );
  inv01 U4875 ( .Y(n11812), .A(n11821) );
  nand02 U4876 ( .Y(n11822), .A0(n11796), .A1(n11797) );
  inv01 U4877 ( .Y(n11814), .A(n11822) );
  nand02 U4878 ( .Y(n11823), .A0(n11799), .A1(n11801) );
  inv01 U4879 ( .Y(n11824), .A(n11823) );
  nand02 U4880 ( .Y(n11825), .A0(n11803), .A1(n11805) );
  inv01 U4881 ( .Y(n11826), .A(n11825) );
  nand02 U4882 ( .Y(n11827), .A0(n11824), .A1(n11826) );
  inv01 U4883 ( .Y(n11791), .A(n11827) );
  nand02 U4884 ( .Y(n11828), .A0(n11807), .A1(n11809) );
  inv01 U4885 ( .Y(n11829), .A(n11828) );
  nand02 U4886 ( .Y(n11830), .A0(n11811), .A1(n11813) );
  inv01 U4887 ( .Y(n11831), .A(n11830) );
  nand02 U4888 ( .Y(n11832), .A0(n11829), .A1(n11831) );
  inv01 U4889 ( .Y(n11792), .A(n11832) );
  inv04 U4890 ( .Y(n13552), .A(n13550) );
  nand02 U4891 ( .Y(n14151), .A0(n11833), .A1(n11834) );
  inv02 U4892 ( .Y(n11835), .A(n14152) );
  inv02 U4893 ( .Y(n11836), .A(n14059) );
  inv02 U4894 ( .Y(n11837), .A(n12797) );
  inv02 U4895 ( .Y(n11838), .A(n13569) );
  inv02 U4896 ( .Y(n11839), .A(n13536) );
  inv02 U4897 ( .Y(n11840), .A(n13573) );
  nand02 U4898 ( .Y(n11841), .A0(n11837), .A1(n11842) );
  nand02 U4899 ( .Y(n11843), .A0(n11838), .A1(n11844) );
  nand02 U4900 ( .Y(n11845), .A0(n11839), .A1(n11846) );
  nand02 U4901 ( .Y(n11847), .A0(n11839), .A1(n11848) );
  nand02 U4902 ( .Y(n11849), .A0(n11840), .A1(n11850) );
  nand02 U4903 ( .Y(n11851), .A0(n11840), .A1(n11852) );
  nand02 U4904 ( .Y(n11853), .A0(n11840), .A1(n11854) );
  nand02 U4905 ( .Y(n11855), .A0(n11840), .A1(n11856) );
  nand02 U4906 ( .Y(n11857), .A0(n11835), .A1(n11836) );
  inv01 U4907 ( .Y(n11842), .A(n11857) );
  nand02 U4908 ( .Y(n11858), .A0(n11835), .A1(n11836) );
  inv01 U4909 ( .Y(n11844), .A(n11858) );
  nand02 U4910 ( .Y(n11859), .A0(n11835), .A1(n11837) );
  inv01 U4911 ( .Y(n11846), .A(n11859) );
  nand02 U4912 ( .Y(n11860), .A0(n11835), .A1(n11838) );
  inv01 U4913 ( .Y(n11848), .A(n11860) );
  nand02 U4914 ( .Y(n11861), .A0(n11836), .A1(n11837) );
  inv01 U4915 ( .Y(n11850), .A(n11861) );
  nand02 U4916 ( .Y(n11862), .A0(n11836), .A1(n11838) );
  inv01 U4917 ( .Y(n11852), .A(n11862) );
  nand02 U4918 ( .Y(n11863), .A0(n11837), .A1(n11839) );
  inv01 U4919 ( .Y(n11854), .A(n11863) );
  nand02 U4920 ( .Y(n11864), .A0(n11838), .A1(n11839) );
  inv01 U4921 ( .Y(n11856), .A(n11864) );
  nand02 U4922 ( .Y(n11865), .A0(n11841), .A1(n11843) );
  inv01 U4923 ( .Y(n11866), .A(n11865) );
  nand02 U4924 ( .Y(n11867), .A0(n11845), .A1(n11847) );
  inv01 U4925 ( .Y(n11868), .A(n11867) );
  nand02 U4926 ( .Y(n11869), .A0(n11866), .A1(n11868) );
  inv01 U4927 ( .Y(n11833), .A(n11869) );
  nand02 U4928 ( .Y(n11870), .A0(n11849), .A1(n11851) );
  inv01 U4929 ( .Y(n11871), .A(n11870) );
  nand02 U4930 ( .Y(n11872), .A0(n11853), .A1(n11855) );
  inv01 U4931 ( .Y(n11873), .A(n11872) );
  nand02 U4932 ( .Y(n11874), .A0(n11871), .A1(n11873) );
  inv01 U4933 ( .Y(n11834), .A(n11874) );
  nand02 U4934 ( .Y(n14184), .A0(n11875), .A1(n11876) );
  inv02 U4935 ( .Y(n11877), .A(n14186) );
  inv02 U4936 ( .Y(n11878), .A(n14173) );
  inv02 U4937 ( .Y(n11879), .A(n14185) );
  inv02 U4938 ( .Y(n11880), .A(n13569) );
  inv02 U4939 ( .Y(n11881), .A(n13552) );
  inv02 U4940 ( .Y(n11882), .A(n13573) );
  nand02 U4941 ( .Y(n11883), .A0(n11879), .A1(n11884) );
  nand02 U4942 ( .Y(n11885), .A0(n11880), .A1(n11886) );
  nand02 U4943 ( .Y(n11887), .A0(n11881), .A1(n11888) );
  nand02 U4944 ( .Y(n11889), .A0(n11881), .A1(n11890) );
  nand02 U4945 ( .Y(n11891), .A0(n11882), .A1(n11892) );
  nand02 U4946 ( .Y(n11893), .A0(n11882), .A1(n11894) );
  nand02 U4947 ( .Y(n11895), .A0(n11882), .A1(n11896) );
  nand02 U4948 ( .Y(n11897), .A0(n11882), .A1(n11898) );
  nand02 U4949 ( .Y(n11899), .A0(n11877), .A1(n11878) );
  inv01 U4950 ( .Y(n11884), .A(n11899) );
  nand02 U4951 ( .Y(n11900), .A0(n11877), .A1(n11878) );
  inv01 U4952 ( .Y(n11886), .A(n11900) );
  nand02 U4953 ( .Y(n11901), .A0(n11877), .A1(n11879) );
  inv01 U4954 ( .Y(n11888), .A(n11901) );
  nand02 U4955 ( .Y(n11902), .A0(n11877), .A1(n11880) );
  inv01 U4956 ( .Y(n11890), .A(n11902) );
  nand02 U4957 ( .Y(n11903), .A0(n11878), .A1(n11879) );
  inv01 U4958 ( .Y(n11892), .A(n11903) );
  nand02 U4959 ( .Y(n11904), .A0(n11878), .A1(n11880) );
  inv01 U4960 ( .Y(n11894), .A(n11904) );
  nand02 U4961 ( .Y(n11905), .A0(n11879), .A1(n11881) );
  inv01 U4962 ( .Y(n11896), .A(n11905) );
  nand02 U4963 ( .Y(n11906), .A0(n11880), .A1(n11881) );
  inv01 U4964 ( .Y(n11898), .A(n11906) );
  nand02 U4965 ( .Y(n11907), .A0(n11883), .A1(n11885) );
  inv01 U4966 ( .Y(n11908), .A(n11907) );
  nand02 U4967 ( .Y(n11909), .A0(n11887), .A1(n11889) );
  inv01 U4968 ( .Y(n11910), .A(n11909) );
  nand02 U4969 ( .Y(n11911), .A0(n11908), .A1(n11910) );
  inv01 U4970 ( .Y(n11875), .A(n11911) );
  nand02 U4971 ( .Y(n11912), .A0(n11891), .A1(n11893) );
  inv01 U4972 ( .Y(n11913), .A(n11912) );
  nand02 U4973 ( .Y(n11914), .A0(n11895), .A1(n11897) );
  inv01 U4974 ( .Y(n11915), .A(n11914) );
  nand02 U4975 ( .Y(n11916), .A0(n11913), .A1(n11915) );
  inv01 U4976 ( .Y(n11876), .A(n11916) );
  nand02 U4977 ( .Y(n14195), .A0(n11917), .A1(n11918) );
  inv02 U4978 ( .Y(n11919), .A(n14197) );
  inv02 U4979 ( .Y(n11920), .A(n14180) );
  inv02 U4980 ( .Y(n11921), .A(n14196) );
  inv02 U4981 ( .Y(n11922), .A(n13569) );
  inv02 U4982 ( .Y(n11923), .A(n13553) );
  inv02 U4983 ( .Y(n11924), .A(n13573) );
  nand02 U4984 ( .Y(n11925), .A0(n11921), .A1(n11926) );
  nand02 U4985 ( .Y(n11927), .A0(n11922), .A1(n11928) );
  nand02 U4986 ( .Y(n11929), .A0(n11923), .A1(n11930) );
  nand02 U4987 ( .Y(n11931), .A0(n11923), .A1(n11932) );
  nand02 U4988 ( .Y(n11933), .A0(n11924), .A1(n11934) );
  nand02 U4989 ( .Y(n11935), .A0(n11924), .A1(n11936) );
  nand02 U4990 ( .Y(n11937), .A0(n11924), .A1(n11938) );
  nand02 U4991 ( .Y(n11939), .A0(n11924), .A1(n11940) );
  nand02 U4992 ( .Y(n11941), .A0(n11919), .A1(n11920) );
  inv01 U4993 ( .Y(n11926), .A(n11941) );
  nand02 U4994 ( .Y(n11942), .A0(n11919), .A1(n11920) );
  inv01 U4995 ( .Y(n11928), .A(n11942) );
  nand02 U4996 ( .Y(n11943), .A0(n11919), .A1(n11921) );
  inv01 U4997 ( .Y(n11930), .A(n11943) );
  nand02 U4998 ( .Y(n11944), .A0(n11919), .A1(n11922) );
  inv01 U4999 ( .Y(n11932), .A(n11944) );
  nand02 U5000 ( .Y(n11945), .A0(n11920), .A1(n11921) );
  inv01 U5001 ( .Y(n11934), .A(n11945) );
  nand02 U5002 ( .Y(n11946), .A0(n11920), .A1(n11922) );
  inv01 U5003 ( .Y(n11936), .A(n11946) );
  nand02 U5004 ( .Y(n11947), .A0(n11921), .A1(n11923) );
  inv01 U5005 ( .Y(n11938), .A(n11947) );
  nand02 U5006 ( .Y(n11948), .A0(n11922), .A1(n11923) );
  inv01 U5007 ( .Y(n11940), .A(n11948) );
  nand02 U5008 ( .Y(n11949), .A0(n11925), .A1(n11927) );
  inv01 U5009 ( .Y(n11950), .A(n11949) );
  nand02 U5010 ( .Y(n11951), .A0(n11929), .A1(n11931) );
  inv01 U5011 ( .Y(n11952), .A(n11951) );
  nand02 U5012 ( .Y(n11953), .A0(n11950), .A1(n11952) );
  inv01 U5013 ( .Y(n11917), .A(n11953) );
  nand02 U5014 ( .Y(n11954), .A0(n11933), .A1(n11935) );
  inv01 U5015 ( .Y(n11955), .A(n11954) );
  nand02 U5016 ( .Y(n11956), .A0(n11937), .A1(n11939) );
  inv01 U5017 ( .Y(n11957), .A(n11956) );
  nand02 U5018 ( .Y(n11958), .A0(n11955), .A1(n11957) );
  inv01 U5019 ( .Y(n11918), .A(n11958) );
  nand02 U5020 ( .Y(n14167), .A0(n11959), .A1(n11960) );
  inv02 U5021 ( .Y(n11961), .A(n14168) );
  inv02 U5022 ( .Y(n11962), .A(n14144) );
  inv02 U5023 ( .Y(n11963), .A(n14077) );
  inv02 U5024 ( .Y(n11964), .A(n13569) );
  inv02 U5025 ( .Y(n11965), .A(n13552) );
  inv02 U5026 ( .Y(n11966), .A(n13573) );
  nand02 U5027 ( .Y(n11967), .A0(n11963), .A1(n11968) );
  nand02 U5028 ( .Y(n11969), .A0(n11964), .A1(n11970) );
  nand02 U5029 ( .Y(n11971), .A0(n11965), .A1(n11972) );
  nand02 U5030 ( .Y(n11973), .A0(n11965), .A1(n11974) );
  nand02 U5031 ( .Y(n11975), .A0(n11966), .A1(n11976) );
  nand02 U5032 ( .Y(n11977), .A0(n11966), .A1(n11978) );
  nand02 U5033 ( .Y(n11979), .A0(n11966), .A1(n11980) );
  nand02 U5034 ( .Y(n11981), .A0(n11966), .A1(n11982) );
  nand02 U5035 ( .Y(n11983), .A0(n11961), .A1(n11962) );
  inv01 U5036 ( .Y(n11968), .A(n11983) );
  nand02 U5037 ( .Y(n11984), .A0(n11961), .A1(n11962) );
  inv01 U5038 ( .Y(n11970), .A(n11984) );
  nand02 U5039 ( .Y(n11985), .A0(n11961), .A1(n11963) );
  inv01 U5040 ( .Y(n11972), .A(n11985) );
  nand02 U5041 ( .Y(n11986), .A0(n11961), .A1(n11964) );
  inv01 U5042 ( .Y(n11974), .A(n11986) );
  nand02 U5043 ( .Y(n11987), .A0(n11962), .A1(n11963) );
  inv01 U5044 ( .Y(n11976), .A(n11987) );
  nand02 U5045 ( .Y(n11988), .A0(n11962), .A1(n11964) );
  inv01 U5046 ( .Y(n11978), .A(n11988) );
  nand02 U5047 ( .Y(n11989), .A0(n11963), .A1(n11965) );
  inv01 U5048 ( .Y(n11980), .A(n11989) );
  nand02 U5049 ( .Y(n11990), .A0(n11964), .A1(n11965) );
  inv01 U5050 ( .Y(n11982), .A(n11990) );
  nand02 U5051 ( .Y(n11991), .A0(n11967), .A1(n11969) );
  inv01 U5052 ( .Y(n11992), .A(n11991) );
  nand02 U5053 ( .Y(n11993), .A0(n11971), .A1(n11973) );
  inv01 U5054 ( .Y(n11994), .A(n11993) );
  nand02 U5055 ( .Y(n11995), .A0(n11992), .A1(n11994) );
  inv01 U5056 ( .Y(n11959), .A(n11995) );
  nand02 U5057 ( .Y(n11996), .A0(n11975), .A1(n11977) );
  inv01 U5058 ( .Y(n11997), .A(n11996) );
  nand02 U5059 ( .Y(n11998), .A0(n11979), .A1(n11981) );
  inv01 U5060 ( .Y(n11999), .A(n11998) );
  nand02 U5061 ( .Y(n12000), .A0(n11997), .A1(n11999) );
  inv01 U5062 ( .Y(n11960), .A(n12000) );
  inv02 U5063 ( .Y(n13553), .A(n13550) );
  nand02 U5064 ( .Y(n14177), .A0(n12001), .A1(n12002) );
  inv02 U5065 ( .Y(n12003), .A(n14178) );
  inv02 U5066 ( .Y(n12004), .A(n14156) );
  inv02 U5067 ( .Y(n12005), .A(n14095) );
  inv02 U5068 ( .Y(n12006), .A(n13569) );
  inv02 U5069 ( .Y(n12007), .A(n13551) );
  inv02 U5070 ( .Y(n12008), .A(n13573) );
  nand02 U5071 ( .Y(n12009), .A0(n12005), .A1(n12010) );
  nand02 U5072 ( .Y(n12011), .A0(n12006), .A1(n12012) );
  nand02 U5073 ( .Y(n12013), .A0(n12007), .A1(n12014) );
  nand02 U5074 ( .Y(n12015), .A0(n12007), .A1(n12016) );
  nand02 U5075 ( .Y(n12017), .A0(n12008), .A1(n12018) );
  nand02 U5076 ( .Y(n12019), .A0(n12008), .A1(n12020) );
  nand02 U5077 ( .Y(n12021), .A0(n12008), .A1(n12022) );
  nand02 U5078 ( .Y(n12023), .A0(n12008), .A1(n12024) );
  nand02 U5079 ( .Y(n12025), .A0(n12003), .A1(n12004) );
  inv01 U5080 ( .Y(n12010), .A(n12025) );
  nand02 U5081 ( .Y(n12026), .A0(n12003), .A1(n12004) );
  inv01 U5082 ( .Y(n12012), .A(n12026) );
  nand02 U5083 ( .Y(n12027), .A0(n12003), .A1(n12005) );
  inv01 U5084 ( .Y(n12014), .A(n12027) );
  nand02 U5085 ( .Y(n12028), .A0(n12003), .A1(n12006) );
  inv01 U5086 ( .Y(n12016), .A(n12028) );
  nand02 U5087 ( .Y(n12029), .A0(n12004), .A1(n12005) );
  inv01 U5088 ( .Y(n12018), .A(n12029) );
  nand02 U5089 ( .Y(n12030), .A0(n12004), .A1(n12006) );
  inv01 U5090 ( .Y(n12020), .A(n12030) );
  nand02 U5091 ( .Y(n12031), .A0(n12005), .A1(n12007) );
  inv01 U5092 ( .Y(n12022), .A(n12031) );
  nand02 U5093 ( .Y(n12032), .A0(n12006), .A1(n12007) );
  inv01 U5094 ( .Y(n12024), .A(n12032) );
  nand02 U5095 ( .Y(n12033), .A0(n12009), .A1(n12011) );
  inv01 U5096 ( .Y(n12034), .A(n12033) );
  nand02 U5097 ( .Y(n12035), .A0(n12013), .A1(n12015) );
  inv01 U5098 ( .Y(n12036), .A(n12035) );
  nand02 U5099 ( .Y(n12037), .A0(n12034), .A1(n12036) );
  inv01 U5100 ( .Y(n12001), .A(n12037) );
  nand02 U5101 ( .Y(n12038), .A0(n12017), .A1(n12019) );
  inv01 U5102 ( .Y(n12039), .A(n12038) );
  nand02 U5103 ( .Y(n12040), .A0(n12021), .A1(n12023) );
  inv01 U5104 ( .Y(n12041), .A(n12040) );
  nand02 U5105 ( .Y(n12042), .A0(n12039), .A1(n12041) );
  inv01 U5106 ( .Y(n12002), .A(n12042) );
  nand02 U5107 ( .Y(n14145), .A0(n12043), .A1(n12044) );
  inv02 U5108 ( .Y(n12045), .A(n14148) );
  inv02 U5109 ( .Y(n12046), .A(n14147) );
  inv02 U5110 ( .Y(n12047), .A(n14146) );
  inv02 U5111 ( .Y(n12048), .A(n13569) );
  inv02 U5112 ( .Y(n12049), .A(n13535) );
  inv02 U5113 ( .Y(n12050), .A(n13573) );
  nand02 U5114 ( .Y(n12051), .A0(n12047), .A1(n12052) );
  nand02 U5115 ( .Y(n12053), .A0(n12048), .A1(n12054) );
  nand02 U5116 ( .Y(n12055), .A0(n12049), .A1(n12056) );
  nand02 U5117 ( .Y(n12057), .A0(n12049), .A1(n12058) );
  nand02 U5118 ( .Y(n12059), .A0(n12050), .A1(n12060) );
  nand02 U5119 ( .Y(n12061), .A0(n12050), .A1(n12062) );
  nand02 U5120 ( .Y(n12063), .A0(n12050), .A1(n12064) );
  nand02 U5121 ( .Y(n12065), .A0(n12050), .A1(n12066) );
  nand02 U5122 ( .Y(n12067), .A0(n12045), .A1(n12046) );
  inv01 U5123 ( .Y(n12052), .A(n12067) );
  nand02 U5124 ( .Y(n12068), .A0(n12045), .A1(n12046) );
  inv01 U5125 ( .Y(n12054), .A(n12068) );
  nand02 U5126 ( .Y(n12069), .A0(n12045), .A1(n12047) );
  inv01 U5127 ( .Y(n12056), .A(n12069) );
  nand02 U5128 ( .Y(n12070), .A0(n12045), .A1(n12048) );
  inv01 U5129 ( .Y(n12058), .A(n12070) );
  nand02 U5130 ( .Y(n12071), .A0(n12046), .A1(n12047) );
  inv01 U5131 ( .Y(n12060), .A(n12071) );
  nand02 U5132 ( .Y(n12072), .A0(n12046), .A1(n12048) );
  inv01 U5133 ( .Y(n12062), .A(n12072) );
  nand02 U5134 ( .Y(n12073), .A0(n12047), .A1(n12049) );
  inv01 U5135 ( .Y(n12064), .A(n12073) );
  nand02 U5136 ( .Y(n12074), .A0(n12048), .A1(n12049) );
  inv01 U5137 ( .Y(n12066), .A(n12074) );
  nand02 U5138 ( .Y(n12075), .A0(n12051), .A1(n12053) );
  inv01 U5139 ( .Y(n12076), .A(n12075) );
  nand02 U5140 ( .Y(n12077), .A0(n12055), .A1(n12057) );
  inv01 U5141 ( .Y(n12078), .A(n12077) );
  nand02 U5142 ( .Y(n12079), .A0(n12076), .A1(n12078) );
  inv01 U5143 ( .Y(n12043), .A(n12079) );
  nand02 U5144 ( .Y(n12080), .A0(n12059), .A1(n12061) );
  inv01 U5145 ( .Y(n12081), .A(n12080) );
  nand02 U5146 ( .Y(n12082), .A0(n12063), .A1(n12065) );
  inv01 U5147 ( .Y(n12083), .A(n12082) );
  nand02 U5148 ( .Y(n12084), .A0(n12081), .A1(n12083) );
  inv01 U5149 ( .Y(n12044), .A(n12084) );
  inv01 U5150 ( .Y(n14381), .A(n12085) );
  inv01 U5151 ( .Y(n12086), .A(s_exp_10a_7_) );
  inv01 U5152 ( .Y(n12087), .A(s_exp_10a_8_) );
  inv01 U5153 ( .Y(n12088), .A(s_exp_10a_6_) );
  inv01 U5154 ( .Y(n12089), .A(n14384) );
  nand02 U5155 ( .Y(n12085), .A0(n12090), .A1(n12091) );
  nand02 U5156 ( .Y(n12092), .A0(n12086), .A1(n12087) );
  inv01 U5157 ( .Y(n12090), .A(n12092) );
  nand02 U5158 ( .Y(n12093), .A0(n12088), .A1(n12089) );
  inv01 U5159 ( .Y(n12091), .A(n12093) );
  nand02 U5160 ( .Y(n14181), .A0(n12094), .A1(n12095) );
  inv02 U5161 ( .Y(n12096), .A(n14165) );
  inv02 U5162 ( .Y(n12097), .A(n14169) );
  inv02 U5163 ( .Y(n12098), .A(n14182) );
  inv02 U5164 ( .Y(n12099), .A(n13573) );
  inv02 U5165 ( .Y(n12100), .A(n13552) );
  inv02 U5166 ( .Y(n12101), .A(n13569) );
  nand02 U5167 ( .Y(n12102), .A0(n12098), .A1(n12103) );
  nand02 U5168 ( .Y(n12104), .A0(n12099), .A1(n12105) );
  nand02 U5169 ( .Y(n12106), .A0(n12100), .A1(n12107) );
  nand02 U5170 ( .Y(n12108), .A0(n12100), .A1(n12109) );
  nand02 U5171 ( .Y(n12110), .A0(n12101), .A1(n12111) );
  nand02 U5172 ( .Y(n12112), .A0(n12101), .A1(n12113) );
  nand02 U5173 ( .Y(n12114), .A0(n12101), .A1(n12115) );
  nand02 U5174 ( .Y(n12116), .A0(n12101), .A1(n12117) );
  nand02 U5175 ( .Y(n12118), .A0(n12096), .A1(n12097) );
  inv01 U5176 ( .Y(n12103), .A(n12118) );
  nand02 U5177 ( .Y(n12119), .A0(n12096), .A1(n12097) );
  inv01 U5178 ( .Y(n12105), .A(n12119) );
  nand02 U5179 ( .Y(n12120), .A0(n12096), .A1(n12098) );
  inv01 U5180 ( .Y(n12107), .A(n12120) );
  nand02 U5181 ( .Y(n12121), .A0(n12096), .A1(n12099) );
  inv01 U5182 ( .Y(n12109), .A(n12121) );
  nand02 U5183 ( .Y(n12122), .A0(n12097), .A1(n12098) );
  inv01 U5184 ( .Y(n12111), .A(n12122) );
  nand02 U5185 ( .Y(n12123), .A0(n12097), .A1(n12099) );
  inv01 U5186 ( .Y(n12113), .A(n12123) );
  nand02 U5187 ( .Y(n12124), .A0(n12098), .A1(n12100) );
  inv01 U5188 ( .Y(n12115), .A(n12124) );
  nand02 U5189 ( .Y(n12125), .A0(n12099), .A1(n12100) );
  inv01 U5190 ( .Y(n12117), .A(n12125) );
  nand02 U5191 ( .Y(n12126), .A0(n12102), .A1(n12104) );
  inv01 U5192 ( .Y(n12127), .A(n12126) );
  nand02 U5193 ( .Y(n12128), .A0(n12106), .A1(n12108) );
  inv01 U5194 ( .Y(n12129), .A(n12128) );
  nand02 U5195 ( .Y(n12130), .A0(n12127), .A1(n12129) );
  inv01 U5196 ( .Y(n12094), .A(n12130) );
  nand02 U5197 ( .Y(n12131), .A0(n12110), .A1(n12112) );
  inv01 U5198 ( .Y(n12132), .A(n12131) );
  nand02 U5199 ( .Y(n12133), .A0(n12114), .A1(n12116) );
  inv01 U5200 ( .Y(n12134), .A(n12133) );
  nand02 U5201 ( .Y(n12135), .A0(n12132), .A1(n12134) );
  inv01 U5202 ( .Y(n12095), .A(n12135) );
  nand02 U5203 ( .Y(n14283), .A0(n12136), .A1(n12137) );
  inv02 U5204 ( .Y(n12138), .A(n13576) );
  inv02 U5205 ( .Y(n12139), .A(n13561) );
  inv02 U5206 ( .Y(n12140), .A(n13557) );
  inv02 U5207 ( .Y(n12141), .A(n14284) );
  inv02 U5208 ( .Y(n12142), .A(n14116) );
  inv02 U5209 ( .Y(n12143), .A(n14285) );
  nand02 U5210 ( .Y(n12144), .A0(n12140), .A1(n12145) );
  nand02 U5211 ( .Y(n12146), .A0(n12141), .A1(n12147) );
  nand02 U5212 ( .Y(n12148), .A0(n12142), .A1(n12149) );
  nand02 U5213 ( .Y(n12150), .A0(n12142), .A1(n12151) );
  nand02 U5214 ( .Y(n12152), .A0(n12143), .A1(n12153) );
  nand02 U5215 ( .Y(n12154), .A0(n12143), .A1(n12155) );
  nand02 U5216 ( .Y(n12156), .A0(n12143), .A1(n12157) );
  nand02 U5217 ( .Y(n12158), .A0(n12143), .A1(n12159) );
  nand02 U5218 ( .Y(n12160), .A0(n12138), .A1(n12139) );
  inv01 U5219 ( .Y(n12145), .A(n12160) );
  nand02 U5220 ( .Y(n12161), .A0(n12138), .A1(n12139) );
  inv01 U5221 ( .Y(n12147), .A(n12161) );
  nand02 U5222 ( .Y(n12162), .A0(n12138), .A1(n12140) );
  inv01 U5223 ( .Y(n12149), .A(n12162) );
  nand02 U5224 ( .Y(n12163), .A0(n12138), .A1(n12141) );
  inv01 U5225 ( .Y(n12151), .A(n12163) );
  nand02 U5226 ( .Y(n12164), .A0(n12139), .A1(n12140) );
  inv01 U5227 ( .Y(n12153), .A(n12164) );
  nand02 U5228 ( .Y(n12165), .A0(n12139), .A1(n12141) );
  inv01 U5229 ( .Y(n12155), .A(n12165) );
  nand02 U5230 ( .Y(n12166), .A0(n12140), .A1(n12142) );
  inv01 U5231 ( .Y(n12157), .A(n12166) );
  nand02 U5232 ( .Y(n12167), .A0(n12141), .A1(n12142) );
  inv01 U5233 ( .Y(n12159), .A(n12167) );
  nand02 U5234 ( .Y(n12168), .A0(n12144), .A1(n12146) );
  inv01 U5235 ( .Y(n12169), .A(n12168) );
  nand02 U5236 ( .Y(n12170), .A0(n12148), .A1(n12150) );
  inv01 U5237 ( .Y(n12171), .A(n12170) );
  nand02 U5238 ( .Y(n12172), .A0(n12169), .A1(n12171) );
  inv01 U5239 ( .Y(n12136), .A(n12172) );
  nand02 U5240 ( .Y(n12173), .A0(n12152), .A1(n12154) );
  inv01 U5241 ( .Y(n12174), .A(n12173) );
  nand02 U5242 ( .Y(n12175), .A0(n12156), .A1(n12158) );
  inv01 U5243 ( .Y(n12176), .A(n12175) );
  nand02 U5244 ( .Y(n12177), .A0(n12174), .A1(n12176) );
  inv01 U5245 ( .Y(n12137), .A(n12177) );
  nand02 U5246 ( .Y(n14359), .A0(n12178), .A1(n12179) );
  inv02 U5247 ( .Y(n12180), .A(n13566) );
  inv02 U5248 ( .Y(n12181), .A(n13560) );
  inv02 U5249 ( .Y(n12182), .A(n13574) );
  inv02 U5250 ( .Y(n12183), .A(n14291) );
  inv02 U5251 ( .Y(n12184), .A(n14187) );
  inv02 U5252 ( .Y(n12185), .A(n14282) );
  nand02 U5253 ( .Y(n12186), .A0(n12182), .A1(n12187) );
  nand02 U5254 ( .Y(n12188), .A0(n12183), .A1(n12189) );
  nand02 U5255 ( .Y(n12190), .A0(n12184), .A1(n12191) );
  nand02 U5256 ( .Y(n12192), .A0(n12184), .A1(n12193) );
  nand02 U5257 ( .Y(n12194), .A0(n12185), .A1(n12195) );
  nand02 U5258 ( .Y(n12196), .A0(n12185), .A1(n12197) );
  nand02 U5259 ( .Y(n12198), .A0(n12185), .A1(n12199) );
  nand02 U5260 ( .Y(n12200), .A0(n12185), .A1(n12201) );
  nand02 U5261 ( .Y(n12202), .A0(n12180), .A1(n12181) );
  inv01 U5262 ( .Y(n12187), .A(n12202) );
  nand02 U5263 ( .Y(n12203), .A0(n12180), .A1(n12181) );
  inv01 U5264 ( .Y(n12189), .A(n12203) );
  nand02 U5265 ( .Y(n12204), .A0(n12180), .A1(n12182) );
  inv01 U5266 ( .Y(n12191), .A(n12204) );
  nand02 U5267 ( .Y(n12205), .A0(n12180), .A1(n12183) );
  inv01 U5268 ( .Y(n12193), .A(n12205) );
  nand02 U5269 ( .Y(n12206), .A0(n12181), .A1(n12182) );
  inv01 U5270 ( .Y(n12195), .A(n12206) );
  nand02 U5271 ( .Y(n12207), .A0(n12181), .A1(n12183) );
  inv01 U5272 ( .Y(n12197), .A(n12207) );
  nand02 U5273 ( .Y(n12208), .A0(n12182), .A1(n12184) );
  inv01 U5274 ( .Y(n12199), .A(n12208) );
  nand02 U5275 ( .Y(n12209), .A0(n12183), .A1(n12184) );
  inv01 U5276 ( .Y(n12201), .A(n12209) );
  nand02 U5277 ( .Y(n12210), .A0(n12186), .A1(n12188) );
  inv01 U5278 ( .Y(n12211), .A(n12210) );
  nand02 U5279 ( .Y(n12212), .A0(n12190), .A1(n12192) );
  inv01 U5280 ( .Y(n12213), .A(n12212) );
  nand02 U5281 ( .Y(n12214), .A0(n12211), .A1(n12213) );
  inv01 U5282 ( .Y(n12178), .A(n12214) );
  nand02 U5283 ( .Y(n12215), .A0(n12194), .A1(n12196) );
  inv01 U5284 ( .Y(n12216), .A(n12215) );
  nand02 U5285 ( .Y(n12217), .A0(n12198), .A1(n12200) );
  inv01 U5286 ( .Y(n12218), .A(n12217) );
  nand02 U5287 ( .Y(n12219), .A0(n12216), .A1(n12218) );
  inv01 U5288 ( .Y(n12179), .A(n12219) );
  inv02 U5289 ( .Y(n14282), .A(n13242) );
  buf02 U5290 ( .Y(n12220), .A(n14390) );
  inv01 U5291 ( .Y(n14378), .A(n12221) );
  inv01 U5292 ( .Y(n12222), .A(s_exp_10b[8]) );
  inv01 U5293 ( .Y(n12223), .A(s_exp_10b[5]) );
  inv01 U5294 ( .Y(n12224), .A(n14379) );
  inv01 U5295 ( .Y(n12225), .A(s_exp_10b[6]) );
  nand02 U5296 ( .Y(n12221), .A0(n12226), .A1(n12227) );
  nand02 U5297 ( .Y(n12228), .A0(n12222), .A1(n12223) );
  inv01 U5298 ( .Y(n12226), .A(n12228) );
  nand02 U5299 ( .Y(n12229), .A0(n12224), .A1(n12225) );
  inv01 U5300 ( .Y(n12227), .A(n12229) );
  inv01 U5301 ( .Y(s_output_o_22_), .A(n12230) );
  nor02 U5302 ( .Y(n12231), .A0(n12280), .A1(n13986) );
  nor02 U5303 ( .Y(n12232), .A0(n12298), .A1(n13985) );
  inv01 U5304 ( .Y(n12233), .A(n13987) );
  nor02 U5305 ( .Y(n12230), .A0(n12233), .A1(n12234) );
  nor02 U5306 ( .Y(n12235), .A0(n12231), .A1(n12232) );
  inv01 U5307 ( .Y(n12234), .A(n12235) );
  nand02 U5308 ( .Y(n13793), .A0(n12236), .A1(n12237) );
  inv01 U5309 ( .Y(n12238), .A(n13809) );
  inv01 U5310 ( .Y(n12239), .A(s_fract_48_i[2]) );
  inv01 U5311 ( .Y(n12240), .A(n13808) );
  inv01 U5312 ( .Y(n12241), .A(n13810) );
  inv01 U5313 ( .Y(n12242), .A(s_fract_48_i[0]) );
  nand02 U5314 ( .Y(n12236), .A0(n12240), .A1(n12243) );
  nand02 U5315 ( .Y(n12237), .A0(n12241), .A1(n12242) );
  nand02 U5316 ( .Y(n12244), .A0(n12238), .A1(n12239) );
  inv01 U5317 ( .Y(n12243), .A(n12244) );
  xor2 U5318 ( .Y(n12245), .A0(s_shr2_4_), .A1(n14395) );
  inv02 U5319 ( .Y(n12246), .A(n12245) );
  inv02 U5320 ( .Y(n13607), .A(n____return5956_4_) );
  inv02 U5321 ( .Y(n13744), .A(n12247) );
  nand02 U5322 ( .Y(n12247), .A0(n10405), .A1(n12248) );
  nand02 U5323 ( .Y(n12249), .A0(n13772), .A1(n13791) );
  inv01 U5324 ( .Y(n12248), .A(n12249) );
  buf02 U5325 ( .Y(n12250), .A(s_fract_48_i[28]) );
  buf02 U5326 ( .Y(n12253), .A(s_fract_48_i[28]) );
  buf02 U5327 ( .Y(n12251), .A(s_fract_48_i[28]) );
  buf02 U5328 ( .Y(n12252), .A(s_fract_48_i[28]) );
  inv02 U5329 ( .Y(n14147), .A(n14359) );
  buf02 U5330 ( .Y(n12254), .A(s_fract_48_i[36]) );
  buf02 U5331 ( .Y(n12257), .A(s_fract_48_i[36]) );
  buf02 U5332 ( .Y(n12255), .A(s_fract_48_i[36]) );
  buf02 U5333 ( .Y(n12256), .A(s_fract_48_i[36]) );
  inv02 U5334 ( .Y(n14085), .A(n14283) );
  inv02 U5335 ( .Y(n13755), .A(n12258) );
  nand02 U5336 ( .Y(n12258), .A0(n10423), .A1(n12259) );
  nand02 U5337 ( .Y(n12260), .A0(n13753), .A1(n13805) );
  inv01 U5338 ( .Y(n12259), .A(n12260) );
  ao22 U5339 ( .Y(n12261), .A0(n14284), .A1(n13576), .B0(n14116), .B1(n13557)
         );
  inv01 U5340 ( .Y(n12262), .A(n12261) );
  nand02 U5341 ( .Y(n12263), .A0(n13535), .A1(n13574) );
  inv02 U5342 ( .Y(n12264), .A(n12263) );
  nand02 U5343 ( .Y(n12265), .A0(n14371), .A1(n11497) );
  inv02 U5344 ( .Y(n12266), .A(n12265) );
  nand02 U5345 ( .Y(n12267), .A0(s_shr2_5_), .A1(n14372) );
  inv02 U5346 ( .Y(n14372), .A(s_shr2_4_) );
  nand02 U5347 ( .Y(n13981), .A0(n12268), .A1(n12269) );
  inv02 U5348 ( .Y(n12270), .A(s_expo1[1]) );
  inv01 U5349 ( .Y(n12271), .A(n____return6651_1_) );
  inv01 U5350 ( .Y(n12272), .A(n13520) );
  nand02 U5351 ( .Y(n12268), .A0(n13520), .A1(n12270) );
  nand02 U5352 ( .Y(n12269), .A0(n12271), .A1(n12272) );
  or04 U5353 ( .Y(n12273), .A0(s_opa_i_11_), .A1(n14005), .A2(s_opa_i_10_), 
        .A3(s_opa_i_0_) );
  inv01 U5354 ( .Y(n12274), .A(n12273) );
  or04 U5355 ( .Y(n12275), .A0(s_frac2a_10_), .A1(n14047), .A2(s_frac2a_0_), 
        .A3(n____return6760) );
  inv01 U5356 ( .Y(n12276), .A(n12275) );
  or04 U5357 ( .Y(n12277), .A0(s_opb_i_11_), .A1(n14009), .A2(s_opb_i_10_), 
        .A3(s_opb_i_0_) );
  inv01 U5358 ( .Y(n12278), .A(n12277) );
  inv01 U5359 ( .Y(n14001), .A(n12279) );
  inv01 U5360 ( .Y(n12280), .A(n13990) );
  inv01 U5361 ( .Y(n12281), .A(s_opa_i_23_) );
  inv01 U5362 ( .Y(n12282), .A(s_opa_i_24_) );
  inv01 U5363 ( .Y(n12283), .A(s_opa_i_25_) );
  nand02 U5364 ( .Y(n12279), .A0(n12284), .A1(n12285) );
  nand02 U5365 ( .Y(n12286), .A0(n12280), .A1(n12281) );
  inv01 U5366 ( .Y(n12284), .A(n12286) );
  nand02 U5367 ( .Y(n12287), .A0(n12282), .A1(n12283) );
  inv01 U5368 ( .Y(n12285), .A(n12287) );
  inv01 U5369 ( .Y(n13945), .A(n12288) );
  inv01 U5370 ( .Y(n12289), .A(n13828) );
  inv01 U5371 ( .Y(n12290), .A(n13827) );
  inv01 U5372 ( .Y(n12291), .A(n12422) );
  inv01 U5373 ( .Y(n12292), .A(n13954) );
  nand02 U5374 ( .Y(n12288), .A0(n12293), .A1(n12294) );
  nand02 U5375 ( .Y(n12295), .A0(n12289), .A1(n12290) );
  inv01 U5376 ( .Y(n12293), .A(n12295) );
  nand02 U5377 ( .Y(n12296), .A0(n12291), .A1(n12292) );
  inv01 U5378 ( .Y(n12294), .A(n12296) );
  inv01 U5379 ( .Y(n14000), .A(n12297) );
  inv01 U5380 ( .Y(n12298), .A(n13991) );
  inv01 U5381 ( .Y(n12299), .A(s_opb_i_23_) );
  inv01 U5382 ( .Y(n12300), .A(s_opb_i_24_) );
  inv01 U5383 ( .Y(n12301), .A(s_opb_i_25_) );
  nand02 U5384 ( .Y(n12297), .A0(n12302), .A1(n12303) );
  nand02 U5385 ( .Y(n12304), .A0(n12298), .A1(n12299) );
  inv01 U5386 ( .Y(n12302), .A(n12304) );
  nand02 U5387 ( .Y(n12305), .A0(n12300), .A1(n12301) );
  inv01 U5388 ( .Y(n12303), .A(n12305) );
  inv02 U5389 ( .Y(s_expo2b[1]), .A(n13981) );
  inv01 U5390 ( .Y(n13773), .A(n12306) );
  inv01 U5391 ( .Y(n12307), .A(n13634) );
  inv01 U5392 ( .Y(n12308), .A(n13633) );
  inv01 U5393 ( .Y(n12309), .A(n13207) );
  inv01 U5394 ( .Y(n12310), .A(n13793) );
  nand02 U5395 ( .Y(n12306), .A0(n12311), .A1(n12312) );
  nand02 U5396 ( .Y(n12313), .A0(n12307), .A1(n12308) );
  inv01 U5397 ( .Y(n12311), .A(n12313) );
  nand02 U5398 ( .Y(n12314), .A0(n12309), .A1(n12310) );
  inv01 U5399 ( .Y(n12312), .A(n12314) );
  nand02 U5400 ( .Y(n13934), .A0(n12315), .A1(n12316) );
  inv02 U5401 ( .Y(n12317), .A(n13848) );
  inv02 U5402 ( .Y(n12318), .A(n13935) );
  inv01 U5403 ( .Y(n12319), .A(n13901) );
  inv01 U5404 ( .Y(n12320), .A(s_fract_48_i[40]) );
  inv01 U5405 ( .Y(n12321), .A(n13745) );
  inv01 U5406 ( .Y(n12322), .A(n12796) );
  nand02 U5407 ( .Y(n12323), .A0(n12319), .A1(n12324) );
  nand02 U5408 ( .Y(n12325), .A0(n12320), .A1(n12326) );
  nand02 U5409 ( .Y(n12327), .A0(n12321), .A1(n12328) );
  nand02 U5410 ( .Y(n12329), .A0(n12322), .A1(n12330) );
  nand02 U5411 ( .Y(n12331), .A0(n12322), .A1(n12332) );
  nand02 U5412 ( .Y(n12333), .A0(n12322), .A1(n12334) );
  nand02 U5413 ( .Y(n12335), .A0(n12317), .A1(n12318) );
  inv01 U5414 ( .Y(n12324), .A(n12335) );
  nand02 U5415 ( .Y(n12336), .A0(n12317), .A1(n12318) );
  inv01 U5416 ( .Y(n12326), .A(n12336) );
  nand02 U5417 ( .Y(n12337), .A0(n12317), .A1(n12318) );
  inv01 U5418 ( .Y(n12328), .A(n12337) );
  nand02 U5419 ( .Y(n12338), .A0(n12317), .A1(n12319) );
  inv01 U5420 ( .Y(n12330), .A(n12338) );
  nand02 U5421 ( .Y(n12339), .A0(n12317), .A1(n12320) );
  inv01 U5422 ( .Y(n12332), .A(n12339) );
  nand02 U5423 ( .Y(n12340), .A0(n12317), .A1(n12321) );
  inv01 U5424 ( .Y(n12334), .A(n12340) );
  nand02 U5425 ( .Y(n12341), .A0(n12323), .A1(n12325) );
  inv01 U5426 ( .Y(n12342), .A(n12341) );
  nand02 U5427 ( .Y(n12343), .A0(n12327), .A1(n12342) );
  inv01 U5428 ( .Y(n12315), .A(n12343) );
  nand02 U5429 ( .Y(n12344), .A0(n12329), .A1(n12331) );
  inv01 U5430 ( .Y(n12345), .A(n12344) );
  nand02 U5431 ( .Y(n12346), .A0(n12333), .A1(n12345) );
  inv01 U5432 ( .Y(n12316), .A(n12346) );
  nand02 U5433 ( .Y(n12347), .A0(n14396), .A1(n13556) );
  buf08 U5434 ( .Y(n13556), .A(n14244) );
  buf02 U5435 ( .Y(n12348), .A(s_fract_48_i[26]) );
  buf02 U5436 ( .Y(n12351), .A(s_fract_48_i[26]) );
  buf02 U5437 ( .Y(n12349), .A(s_fract_48_i[26]) );
  buf02 U5438 ( .Y(n12350), .A(s_fract_48_i[26]) );
  or04 U5439 ( .Y(n12352), .A0(n14004), .A1(s_opa_i_14_), .A2(s_opa_i_16_), 
        .A3(s_opa_i_15_) );
  inv01 U5440 ( .Y(n12353), .A(n12352) );
  or04 U5441 ( .Y(n12354), .A0(n14046), .A1(s_frac2a_13_), .A2(s_frac2a_15_), 
        .A3(s_frac2a_14_) );
  inv01 U5442 ( .Y(n12355), .A(n12354) );
  or04 U5443 ( .Y(n12356), .A0(n14008), .A1(s_opb_i_14_), .A2(s_opb_i_16_), 
        .A3(s_opb_i_15_) );
  inv01 U5444 ( .Y(n12357), .A(n12356) );
  or04 U5445 ( .Y(n12358), .A0(n14003), .A1(s_opa_i_1_), .A2(s_opa_i_21_), 
        .A3(s_opa_i_20_) );
  inv01 U5446 ( .Y(n12359), .A(n12358) );
  or04 U5447 ( .Y(n12360), .A0(n14007), .A1(s_opb_i_1_), .A2(s_opb_i_21_), 
        .A3(s_opb_i_20_) );
  inv01 U5448 ( .Y(n12361), .A(n12360) );
  or04 U5449 ( .Y(n12362), .A0(s_frac2a_20_), .A1(n14045), .A2(s_frac2a_1_), 
        .A3(s_frac2a_19_) );
  inv01 U5450 ( .Y(n12363), .A(n12362) );
  xor2 U5451 ( .Y(n12364), .A0(n10295), .A1(n14353) );
  inv02 U5452 ( .Y(n12365), .A(n12364) );
  inv01 U5453 ( .Y(n13774), .A(n12366) );
  inv01 U5454 ( .Y(n12367), .A(n13209) );
  inv01 U5455 ( .Y(n12368), .A(n13635) );
  inv01 U5456 ( .Y(n12369), .A(n13636) );
  inv01 U5457 ( .Y(n12370), .A(n13787) );
  nand02 U5458 ( .Y(n12366), .A0(n12371), .A1(n12372) );
  nand02 U5459 ( .Y(n12373), .A0(n12367), .A1(n12368) );
  inv01 U5460 ( .Y(n12371), .A(n12373) );
  nand02 U5461 ( .Y(n12374), .A0(n12369), .A1(n12370) );
  inv01 U5462 ( .Y(n12372), .A(n12374) );
  inv01 U5463 ( .Y(n13946), .A(n12375) );
  inv01 U5464 ( .Y(n12376), .A(n13831) );
  inv01 U5465 ( .Y(n12377), .A(n13834) );
  inv01 U5466 ( .Y(n12378), .A(n13833) );
  inv01 U5467 ( .Y(n12379), .A(n13953) );
  nand02 U5468 ( .Y(n12375), .A0(n12380), .A1(n12381) );
  nand02 U5469 ( .Y(n12382), .A0(n12376), .A1(n12377) );
  inv01 U5470 ( .Y(n12380), .A(n12382) );
  nand02 U5471 ( .Y(n12383), .A0(n12378), .A1(n12379) );
  inv01 U5472 ( .Y(n12381), .A(n12383) );
  inv02 U5473 ( .Y(n13644), .A(n12384) );
  nand02 U5474 ( .Y(n12384), .A0(n12385), .A1(n12386) );
  nand02 U5475 ( .Y(n12387), .A0(s_fract_48_i[46]), .A1(n10338) );
  inv01 U5476 ( .Y(n12385), .A(n12387) );
  nand02 U5477 ( .Y(n12388), .A0(n13746), .A1(n13747) );
  inv01 U5478 ( .Y(n12386), .A(n12388) );
  inv02 U5479 ( .Y(n13747), .A(s_fract_48_i[45]) );
  nor02 U5480 ( .Y(n13775), .A0(n12389), .A1(n12390) );
  nor02 U5481 ( .Y(n12391), .A0(n13781), .A1(n13624) );
  inv01 U5482 ( .Y(n12389), .A(n12391) );
  nor02 U5483 ( .Y(n12392), .A0(n13625), .A1(n13622) );
  inv01 U5484 ( .Y(n12390), .A(n12392) );
  inv01 U5485 ( .Y(n13947), .A(n12393) );
  inv01 U5486 ( .Y(n12394), .A(n13816) );
  inv01 U5487 ( .Y(n12395), .A(n13818) );
  inv01 U5488 ( .Y(n12396), .A(n10279) );
  inv01 U5489 ( .Y(n12397), .A(n13950) );
  nand02 U5490 ( .Y(n12393), .A0(n12398), .A1(n12399) );
  nand02 U5491 ( .Y(n12400), .A0(n12394), .A1(n12395) );
  inv01 U5492 ( .Y(n12398), .A(n12400) );
  nand02 U5493 ( .Y(n12401), .A0(n12396), .A1(n12397) );
  inv01 U5494 ( .Y(n12399), .A(n12401) );
  or04 U5495 ( .Y(n12402), .A0(n14002), .A1(s_opa_i_4_), .A2(s_opa_i_6_), .A3(
        s_opa_i_5_) );
  inv01 U5496 ( .Y(n12403), .A(n12402) );
  or04 U5497 ( .Y(n12404), .A0(n14044), .A1(s_frac2a_4_), .A2(s_frac2a_6_), 
        .A3(s_frac2a_5_) );
  inv01 U5498 ( .Y(n12405), .A(n12404) );
  or04 U5499 ( .Y(n12406), .A0(n14006), .A1(s_opb_i_4_), .A2(s_opb_i_6_), .A3(
        s_opb_i_5_) );
  inv01 U5500 ( .Y(n12407), .A(n12406) );
  buf02 U5501 ( .Y(n12408), .A(s_fract_48_i[25]) );
  buf02 U5502 ( .Y(n12411), .A(s_fract_48_i[25]) );
  buf02 U5503 ( .Y(n12409), .A(s_fract_48_i[25]) );
  buf02 U5504 ( .Y(n12410), .A(s_fract_48_i[25]) );
  or04 U5505 ( .Y(n12412), .A0(n13978), .A1(n13976), .A2(n13974), .A3(n13969)
         );
  inv01 U5506 ( .Y(n12413), .A(n12412) );
  inv02 U5507 ( .Y(n13830), .A(n13919) );
  inv02 U5508 ( .Y(n12414), .A(n13960) );
  inv08 U5509 ( .Y(n12415), .A(n12414) );
  inv01 U5510 ( .Y(n12416), .A(n12414) );
  buf02 U5511 ( .Y(n12417), .A(s_fract_48_i[20]) );
  buf02 U5512 ( .Y(n12420), .A(s_fract_48_i[20]) );
  buf02 U5513 ( .Y(n12418), .A(s_fract_48_i[20]) );
  buf02 U5514 ( .Y(n12419), .A(s_fract_48_i[20]) );
  nand02 U5515 ( .Y(n12421), .A0(s_fract_48_i[17]), .A1(n13955) );
  inv02 U5516 ( .Y(n12422), .A(n12421) );
  nor02 U5517 ( .Y(n14013), .A0(n12423), .A1(n12424) );
  nor02 U5518 ( .Y(n12425), .A0(n13979), .A1(n13977) );
  inv02 U5519 ( .Y(n12423), .A(n12425) );
  nor02 U5520 ( .Y(n12426), .A0(n13975), .A1(n13971) );
  inv01 U5521 ( .Y(n12424), .A(n12426) );
  inv02 U5522 ( .Y(n13979), .A(n____return7168_4_) );
  inv01 U5523 ( .Y(n13776), .A(n12427) );
  inv01 U5524 ( .Y(n12428), .A(n12470) );
  inv01 U5525 ( .Y(n12429), .A(n13628) );
  inv01 U5526 ( .Y(n12430), .A(n13626) );
  inv01 U5527 ( .Y(n12431), .A(n13777) );
  nand02 U5528 ( .Y(n12427), .A0(n12432), .A1(n12433) );
  nand02 U5529 ( .Y(n12434), .A0(n12428), .A1(n12429) );
  inv01 U5530 ( .Y(n12432), .A(n12434) );
  nand02 U5531 ( .Y(n12435), .A0(n12430), .A1(n12431) );
  inv01 U5532 ( .Y(n12433), .A(n12435) );
  inv01 U5533 ( .Y(n13948), .A(n12436) );
  inv01 U5534 ( .Y(n12437), .A(n13823) );
  inv01 U5535 ( .Y(n12438), .A(n13820) );
  inv01 U5536 ( .Y(n12439), .A(n13949) );
  nand02 U5537 ( .Y(n12436), .A0(n12440), .A1(n12441) );
  nand02 U5538 ( .Y(n12442), .A0(n12437), .A1(n13908) );
  inv01 U5539 ( .Y(n12440), .A(n12442) );
  nand02 U5540 ( .Y(n12443), .A0(n12438), .A1(n12439) );
  inv01 U5541 ( .Y(n12441), .A(n12443) );
  or03 U5542 ( .Y(n12444), .A0(n13902), .A1(s_fract_48_i[39]), .A2(n13938) );
  inv01 U5543 ( .Y(n12445), .A(n12444) );
  or03 U5544 ( .Y(n12446), .A0(n14366), .A1(s_shr2_5_), .A2(n14340) );
  inv01 U5545 ( .Y(n12447), .A(n12446) );
  inv02 U5546 ( .Y(n12448), .A(n13958) );
  inv08 U5547 ( .Y(n12449), .A(n12448) );
  inv01 U5548 ( .Y(n12450), .A(n12448) );
  or03 U5549 ( .Y(n12451), .A0(n13848), .A1(n13847), .A2(n13849) );
  inv01 U5550 ( .Y(n12452), .A(n12451) );
  inv01 U5551 ( .Y(n13952), .A(n12453) );
  inv01 U5552 ( .Y(n12454), .A(n10575) );
  inv01 U5553 ( .Y(n12455), .A(n10290) );
  inv01 U5554 ( .Y(n12456), .A(n12253) );
  nand02 U5555 ( .Y(n12453), .A0(n12456), .A1(n12457) );
  nand02 U5556 ( .Y(n12458), .A0(n12454), .A1(n12455) );
  inv01 U5557 ( .Y(n12457), .A(n12458) );
  buf02 U5558 ( .Y(n12459), .A(s_fract_48_i[24]) );
  buf02 U5559 ( .Y(n12462), .A(s_fract_48_i[24]) );
  buf02 U5560 ( .Y(n12460), .A(s_fract_48_i[24]) );
  buf02 U5561 ( .Y(n12461), .A(s_fract_48_i[24]) );
  inv01 U5562 ( .Y(n13998), .A(n12463) );
  inv01 U5563 ( .Y(n12464), .A(n10300) );
  inv01 U5564 ( .Y(n12465), .A(s_round) );
  inv01 U5565 ( .Y(n12466), .A(n14489) );
  nand02 U5566 ( .Y(n12463), .A0(n12466), .A1(n12467) );
  nand02 U5567 ( .Y(n12468), .A0(n12464), .A1(n12465) );
  inv01 U5568 ( .Y(n12467), .A(n12468) );
  nand02 U5569 ( .Y(n12469), .A0(s_fract_48_i[23]), .A1(n13778) );
  inv02 U5570 ( .Y(n12470), .A(n12469) );
  or02 U5571 ( .Y(n12471), .A0(n13537), .A1(n13612) );
  inv02 U5572 ( .Y(n12472), .A(n12471) );
  or02 U5573 ( .Y(n12473), .A0(n13537), .A1(n13603) );
  inv02 U5574 ( .Y(n12474), .A(n12473) );
  or02 U5575 ( .Y(n12475), .A0(n13537), .A1(n13606) );
  inv02 U5576 ( .Y(n12476), .A(n12475) );
  or02 U5577 ( .Y(n12477), .A0(n13537), .A1(n13610) );
  inv02 U5578 ( .Y(n12478), .A(n12477) );
  or02 U5579 ( .Y(n12479), .A0(n13537), .A1(n13608) );
  inv02 U5580 ( .Y(n12480), .A(n12479) );
  nand02 U5581 ( .Y(n13999), .A0(n12481), .A1(n12482) );
  inv02 U5582 ( .Y(n12483), .A(n14001) );
  inv02 U5583 ( .Y(n12484), .A(n14000) );
  inv02 U5584 ( .Y(n12485), .A(n10394) );
  inv02 U5585 ( .Y(n12486), .A(n14435) );
  inv02 U5586 ( .Y(n12487), .A(n14434) );
  inv02 U5587 ( .Y(n12488), .A(n10392) );
  inv02 U5588 ( .Y(n12489), .A(n14448) );
  inv02 U5589 ( .Y(n12490), .A(n14447) );
  nand02 U5590 ( .Y(n12491), .A0(n12483), .A1(n12484) );
  nand02 U5591 ( .Y(n12492), .A0(n12483), .A1(n12485) );
  nand02 U5592 ( .Y(n12493), .A0(n12483), .A1(n12486) );
  nand02 U5593 ( .Y(n12494), .A0(n12483), .A1(n12487) );
  nand02 U5594 ( .Y(n12495), .A0(n12484), .A1(n12488) );
  nand02 U5595 ( .Y(n12496), .A0(n12485), .A1(n12488) );
  nand02 U5596 ( .Y(n12497), .A0(n12486), .A1(n12488) );
  nand02 U5597 ( .Y(n12498), .A0(n12487), .A1(n12488) );
  nand02 U5598 ( .Y(n12499), .A0(n12484), .A1(n12489) );
  nand02 U5599 ( .Y(n12500), .A0(n12485), .A1(n12489) );
  nand02 U5600 ( .Y(n12501), .A0(n12486), .A1(n12489) );
  nand02 U5601 ( .Y(n12502), .A0(n12487), .A1(n12489) );
  nand02 U5602 ( .Y(n12503), .A0(n12484), .A1(n12490) );
  nand02 U5603 ( .Y(n12504), .A0(n12485), .A1(n12490) );
  nand02 U5604 ( .Y(n12505), .A0(n12486), .A1(n12490) );
  nand02 U5605 ( .Y(n12506), .A0(n12487), .A1(n12490) );
  nand02 U5606 ( .Y(n12507), .A0(n12491), .A1(n12492) );
  inv01 U5607 ( .Y(n12508), .A(n12507) );
  nand02 U5608 ( .Y(n12509), .A0(n12493), .A1(n12494) );
  inv01 U5609 ( .Y(n12510), .A(n12509) );
  nand02 U5610 ( .Y(n12511), .A0(n12508), .A1(n12510) );
  inv01 U5611 ( .Y(n12512), .A(n12511) );
  nand02 U5612 ( .Y(n12513), .A0(n12495), .A1(n12496) );
  inv01 U5613 ( .Y(n12514), .A(n12513) );
  nand02 U5614 ( .Y(n12515), .A0(n12497), .A1(n12498) );
  inv01 U5615 ( .Y(n12516), .A(n12515) );
  nand02 U5616 ( .Y(n12517), .A0(n12514), .A1(n12516) );
  inv01 U5617 ( .Y(n12518), .A(n12517) );
  nand02 U5618 ( .Y(n12519), .A0(n12512), .A1(n12518) );
  inv01 U5619 ( .Y(n12481), .A(n12519) );
  nand02 U5620 ( .Y(n12520), .A0(n12499), .A1(n12500) );
  inv01 U5621 ( .Y(n12521), .A(n12520) );
  nand02 U5622 ( .Y(n12522), .A0(n12501), .A1(n12502) );
  inv01 U5623 ( .Y(n12523), .A(n12522) );
  nand02 U5624 ( .Y(n12524), .A0(n12521), .A1(n12523) );
  inv01 U5625 ( .Y(n12525), .A(n12524) );
  nand02 U5626 ( .Y(n12526), .A0(n12503), .A1(n12504) );
  inv01 U5627 ( .Y(n12527), .A(n12526) );
  nand02 U5628 ( .Y(n12528), .A0(n12505), .A1(n12506) );
  inv01 U5629 ( .Y(n12529), .A(n12528) );
  nand02 U5630 ( .Y(n12530), .A0(n12527), .A1(n12529) );
  inv01 U5631 ( .Y(n12531), .A(n12530) );
  nand02 U5632 ( .Y(n12532), .A0(n12525), .A1(n12531) );
  inv01 U5633 ( .Y(n12482), .A(n12532) );
  inv01 U5634 ( .Y(n14231), .A(n12533) );
  nor02 U5635 ( .Y(n12534), .A0(n14302), .A1(n13577) );
  nor02 U5636 ( .Y(n12535), .A0(n14301), .A1(n13562) );
  inv01 U5637 ( .Y(n12536), .A(n9896) );
  nor02 U5638 ( .Y(n12533), .A0(n12536), .A1(n12537) );
  nor02 U5639 ( .Y(n12538), .A0(n12534), .A1(n12535) );
  inv01 U5640 ( .Y(n12537), .A(n12538) );
  inv01 U5641 ( .Y(n14186), .A(n12539) );
  nor02 U5642 ( .Y(n12540), .A0(n14326), .A1(n13567) );
  nor02 U5643 ( .Y(n12541), .A0(n14290), .A1(n13575) );
  inv01 U5644 ( .Y(n12542), .A(n9871) );
  nor02 U5645 ( .Y(n12539), .A0(n12542), .A1(n12543) );
  nor02 U5646 ( .Y(n12544), .A0(n12540), .A1(n12541) );
  inv01 U5647 ( .Y(n12543), .A(n12544) );
  inv01 U5648 ( .Y(n14192), .A(n12545) );
  nor02 U5649 ( .Y(n12546), .A0(n13423), .A1(n14204) );
  nor02 U5650 ( .Y(n12547), .A0(n14297), .A1(n13575) );
  inv01 U5651 ( .Y(n12548), .A(n9862) );
  nor02 U5652 ( .Y(n12545), .A0(n12548), .A1(n12549) );
  nor02 U5653 ( .Y(n12550), .A0(n12546), .A1(n12547) );
  inv01 U5654 ( .Y(n12549), .A(n12550) );
  inv01 U5655 ( .Y(n14155), .A(n12551) );
  nor02 U5656 ( .Y(n12552), .A0(n14266), .A1(n13567) );
  nor02 U5657 ( .Y(n12553), .A0(n14228), .A1(n13575) );
  inv01 U5658 ( .Y(n12554), .A(n9788) );
  nor02 U5659 ( .Y(n12551), .A0(n12554), .A1(n12555) );
  nor02 U5660 ( .Y(n12556), .A0(n12552), .A1(n12553) );
  inv01 U5661 ( .Y(n12555), .A(n12556) );
  inv01 U5662 ( .Y(n14197), .A(n12557) );
  nor02 U5663 ( .Y(n12558), .A0(n14254), .A1(n14204) );
  nor02 U5664 ( .Y(n12559), .A0(n14304), .A1(n13575) );
  inv01 U5665 ( .Y(n12560), .A(n14331) );
  nor02 U5666 ( .Y(n12557), .A0(n12560), .A1(n12561) );
  nor02 U5667 ( .Y(n12562), .A0(n12558), .A1(n12559) );
  inv01 U5668 ( .Y(n12561), .A(n12562) );
  inv01 U5669 ( .Y(n14055), .A(n12563) );
  nor02 U5670 ( .Y(n12564), .A0(n14243), .A1(n13577) );
  nor02 U5671 ( .Y(n12565), .A0(n14242), .A1(n13562) );
  inv01 U5672 ( .Y(n12566), .A(n9923) );
  nor02 U5673 ( .Y(n12563), .A0(n12566), .A1(n12567) );
  nor02 U5674 ( .Y(n12568), .A0(n12564), .A1(n12565) );
  inv01 U5675 ( .Y(n12567), .A(n12568) );
  inv01 U5676 ( .Y(n14094), .A(n12569) );
  nor02 U5677 ( .Y(n12570), .A0(n14303), .A1(n13577) );
  nor02 U5678 ( .Y(n12571), .A0(n14302), .A1(n13562) );
  inv01 U5679 ( .Y(n12572), .A(n9860) );
  nor02 U5680 ( .Y(n12569), .A0(n12572), .A1(n12573) );
  nor02 U5681 ( .Y(n12574), .A0(n12570), .A1(n12571) );
  inv01 U5682 ( .Y(n12573), .A(n12574) );
  inv01 U5683 ( .Y(n14076), .A(n12575) );
  nor02 U5684 ( .Y(n12576), .A0(n14275), .A1(n13577) );
  nor02 U5685 ( .Y(n12577), .A0(n14274), .A1(n13562) );
  inv01 U5686 ( .Y(n12578), .A(n9925) );
  nor02 U5687 ( .Y(n12575), .A0(n12578), .A1(n12579) );
  nor02 U5688 ( .Y(n12580), .A0(n12576), .A1(n12577) );
  inv01 U5689 ( .Y(n12579), .A(n12580) );
  inv01 U5690 ( .Y(n14084), .A(n12581) );
  nor02 U5691 ( .Y(n12582), .A0(n14287), .A1(n13577) );
  nor02 U5692 ( .Y(n12583), .A0(n14286), .A1(n13562) );
  inv01 U5693 ( .Y(n12584), .A(n9754) );
  nor02 U5694 ( .Y(n12581), .A0(n12584), .A1(n12585) );
  nor02 U5695 ( .Y(n12586), .A0(n12582), .A1(n12583) );
  inv01 U5696 ( .Y(n12585), .A(n12586) );
  inv01 U5697 ( .Y(n14212), .A(n12587) );
  nor02 U5698 ( .Y(n12588), .A0(n14286), .A1(n13577) );
  nor02 U5699 ( .Y(n12589), .A0(n14322), .A1(n13562) );
  inv01 U5700 ( .Y(n12590), .A(n9866) );
  nor02 U5701 ( .Y(n12587), .A0(n12590), .A1(n12591) );
  nor02 U5702 ( .Y(n12592), .A0(n12588), .A1(n12589) );
  inv01 U5703 ( .Y(n12591), .A(n12592) );
  inv01 U5704 ( .Y(n14205), .A(n12593) );
  nor02 U5705 ( .Y(n12594), .A0(n14272), .A1(n13562) );
  nor02 U5706 ( .Y(n12595), .A0(n14317), .A1(n13558) );
  inv01 U5707 ( .Y(n12596), .A(n9806) );
  nor02 U5708 ( .Y(n12593), .A0(n12596), .A1(n12597) );
  nor02 U5709 ( .Y(n12598), .A0(n12594), .A1(n12595) );
  inv01 U5710 ( .Y(n12597), .A(n12598) );
  inv04 U5711 ( .Y(n13558), .A(n13557) );
  inv01 U5712 ( .Y(n14309), .A(n12599) );
  nor02 U5713 ( .Y(n12600), .A0(n14294), .A1(n13558) );
  nor02 U5714 ( .Y(n12601), .A0(n14328), .A1(n13577) );
  inv01 U5715 ( .Y(n12602), .A(n9846) );
  nor02 U5716 ( .Y(n12599), .A0(n12602), .A1(n12603) );
  nor02 U5717 ( .Y(n12604), .A0(n12600), .A1(n12601) );
  inv01 U5718 ( .Y(n12603), .A(n12604) );
  inv01 U5719 ( .Y(n14088), .A(n12605) );
  nor02 U5720 ( .Y(n12606), .A0(n14294), .A1(n13577) );
  nor02 U5721 ( .Y(n12607), .A0(n14243), .A1(n13558) );
  inv01 U5722 ( .Y(n12608), .A(n14295) );
  nor02 U5723 ( .Y(n12605), .A0(n12608), .A1(n12609) );
  nor02 U5724 ( .Y(n12610), .A0(n12606), .A1(n12607) );
  inv01 U5725 ( .Y(n12609), .A(n12610) );
  inv01 U5726 ( .Y(n14083), .A(n12611) );
  nor02 U5727 ( .Y(n12612), .A0(n13942), .A1(n13582) );
  nor02 U5728 ( .Y(n12613), .A0(n13782), .A1(n13598) );
  inv01 U5729 ( .Y(n12614), .A(n14219) );
  nor02 U5730 ( .Y(n12611), .A0(n12614), .A1(n12615) );
  nor02 U5731 ( .Y(n12616), .A0(n12612), .A1(n12613) );
  inv01 U5732 ( .Y(n12615), .A(n12616) );
  inv01 U5733 ( .Y(n14166), .A(n12617) );
  nor02 U5734 ( .Y(n12618), .A0(n14315), .A1(n13577) );
  nor02 U5735 ( .Y(n12619), .A0(n14275), .A1(n13558) );
  inv01 U5736 ( .Y(n12620), .A(n9830) );
  nor02 U5737 ( .Y(n12617), .A0(n12620), .A1(n12621) );
  nor02 U5738 ( .Y(n12622), .A0(n12618), .A1(n12619) );
  inv01 U5739 ( .Y(n12621), .A(n12622) );
  inv01 U5740 ( .Y(n14220), .A(n12623) );
  nor02 U5741 ( .Y(n12624), .A0(n14287), .A1(n13558) );
  nor02 U5742 ( .Y(n12625), .A0(n14323), .A1(n13577) );
  inv01 U5743 ( .Y(n12626), .A(n9832) );
  nor02 U5744 ( .Y(n12623), .A0(n12626), .A1(n12627) );
  nor02 U5745 ( .Y(n12628), .A0(n12624), .A1(n12625) );
  inv01 U5746 ( .Y(n12627), .A(n12628) );
  inv01 U5747 ( .Y(n14128), .A(n12629) );
  nor02 U5748 ( .Y(n12630), .A0(n13772), .A1(n13580) );
  nor02 U5749 ( .Y(n12631), .A0(n13791), .A1(n13596) );
  inv01 U5750 ( .Y(n12632), .A(n10067) );
  nor02 U5751 ( .Y(n12629), .A0(n12632), .A1(n12633) );
  nor02 U5752 ( .Y(n12634), .A0(n12630), .A1(n12631) );
  inv01 U5753 ( .Y(n12633), .A(n12634) );
  inv02 U5754 ( .Y(n14330), .A(n12635) );
  nor02 U5755 ( .Y(n12636), .A0(n14303), .A1(n13558) );
  nor02 U5756 ( .Y(n12637), .A0(n14370), .A1(n13577) );
  inv01 U5757 ( .Y(n12638), .A(n9907) );
  nor02 U5758 ( .Y(n12635), .A0(n12638), .A1(n12639) );
  nor02 U5759 ( .Y(n12640), .A0(n12636), .A1(n12637) );
  inv01 U5760 ( .Y(n12639), .A(n12640) );
  inv01 U5761 ( .Y(n14075), .A(n12641) );
  nor02 U5762 ( .Y(n12642), .A0(n13806), .A1(n13583) );
  nor02 U5763 ( .Y(n12643), .A0(n13942), .A1(n13599) );
  inv01 U5764 ( .Y(n12644), .A(n9656) );
  nor02 U5765 ( .Y(n12641), .A0(n12644), .A1(n12645) );
  nor02 U5766 ( .Y(n12646), .A0(n12642), .A1(n12643) );
  inv01 U5767 ( .Y(n12645), .A(n12646) );
  inv01 U5768 ( .Y(n14091), .A(n12647) );
  nor02 U5769 ( .Y(n12648), .A0(n13782), .A1(n13583) );
  nor02 U5770 ( .Y(n12649), .A0(n13754), .A1(n13599) );
  inv01 U5771 ( .Y(n12650), .A(n9662) );
  nor02 U5772 ( .Y(n12647), .A0(n12650), .A1(n12651) );
  nor02 U5773 ( .Y(n12652), .A0(n12648), .A1(n12649) );
  inv01 U5774 ( .Y(n12651), .A(n12652) );
  inv01 U5775 ( .Y(n14120), .A(n12653) );
  nor02 U5776 ( .Y(n12654), .A0(n13791), .A1(n13580) );
  nor02 U5777 ( .Y(n12655), .A0(n13745), .A1(n13595) );
  inv01 U5778 ( .Y(n12656), .A(n14149) );
  nor02 U5779 ( .Y(n12653), .A0(n12656), .A1(n12657) );
  nor02 U5780 ( .Y(n12658), .A0(n12654), .A1(n12655) );
  inv01 U5781 ( .Y(n12657), .A(n12658) );
  nand02 U5782 ( .Y(n14136), .A0(n9766), .A1(n12659) );
  inv01 U5783 ( .Y(n12660), .A(n13792) );
  inv01 U5784 ( .Y(n12661), .A(n13595) );
  inv01 U5785 ( .Y(n12662), .A(n13772) );
  nand02 U5786 ( .Y(n12663), .A0(n9630), .A1(n12660) );
  nand02 U5787 ( .Y(n12664), .A0(n12661), .A1(n12662) );
  nand02 U5788 ( .Y(n12665), .A0(n12663), .A1(n12664) );
  inv01 U5789 ( .Y(n12659), .A(n12665) );
  inv02 U5790 ( .Y(n13782), .A(n12923) );
  inv02 U5791 ( .Y(n13772), .A(s_fract_48_i[39]) );
  inv01 U5792 ( .Y(n14168), .A(n12666) );
  nor02 U5793 ( .Y(n12667), .A0(n14279), .A1(n13567) );
  nor02 U5794 ( .Y(n12668), .A0(n14234), .A1(n13575) );
  inv01 U5795 ( .Y(n12669), .A(n9790) );
  nor02 U5796 ( .Y(n12666), .A0(n12669), .A1(n12670) );
  nor02 U5797 ( .Y(n12671), .A0(n12667), .A1(n12668) );
  inv01 U5798 ( .Y(n12670), .A(n12671) );
  inv01 U5799 ( .Y(n14178), .A(n12672) );
  nor02 U5800 ( .Y(n12673), .A0(n14304), .A1(n13567) );
  nor02 U5801 ( .Y(n12674), .A0(n14266), .A1(n13575) );
  inv01 U5802 ( .Y(n12675), .A(n9824) );
  nor02 U5803 ( .Y(n12672), .A0(n12675), .A1(n12676) );
  nor02 U5804 ( .Y(n12677), .A0(n12673), .A1(n12674) );
  inv01 U5805 ( .Y(n12676), .A(n12677) );
  inv01 U5806 ( .Y(n14175), .A(n12678) );
  nor02 U5807 ( .Y(n12679), .A0(n14297), .A1(n13567) );
  nor02 U5808 ( .Y(n12680), .A0(n14249), .A1(n13575) );
  inv01 U5809 ( .Y(n12681), .A(n9808) );
  nor02 U5810 ( .Y(n12678), .A0(n12681), .A1(n12682) );
  nor02 U5811 ( .Y(n12683), .A0(n12679), .A1(n12680) );
  inv01 U5812 ( .Y(n12682), .A(n12683) );
  inv01 U5813 ( .Y(n14110), .A(n12684) );
  nor02 U5814 ( .Y(n12685), .A0(n14208), .A1(n13567) );
  nor02 U5815 ( .Y(n12686), .A0(n14207), .A1(n13575) );
  inv01 U5816 ( .Y(n12687), .A(n9796) );
  nor02 U5817 ( .Y(n12684), .A0(n12687), .A1(n12688) );
  nor02 U5818 ( .Y(n12689), .A0(n12685), .A1(n12686) );
  inv01 U5819 ( .Y(n12688), .A(n12689) );
  inv02 U5820 ( .Y(n13816), .A(n12690) );
  nand02 U5821 ( .Y(n12690), .A0(s_fract_48_i[31]), .A1(n12691) );
  nand02 U5822 ( .Y(n12692), .A0(n10306), .A1(n13794) );
  inv01 U5823 ( .Y(n12691), .A(n12692) );
  inv01 U5824 ( .Y(n14172), .A(n12693) );
  nor02 U5825 ( .Y(n12694), .A0(n14290), .A1(n13567) );
  nor02 U5826 ( .Y(n12695), .A0(n14236), .A1(n13575) );
  inv01 U5827 ( .Y(n12696), .A(n9792) );
  nor02 U5828 ( .Y(n12693), .A0(n12696), .A1(n12697) );
  nor02 U5829 ( .Y(n12698), .A0(n12694), .A1(n12695) );
  inv01 U5830 ( .Y(n12697), .A(n12698) );
  inv01 U5831 ( .Y(n14152), .A(n12699) );
  nor02 U5832 ( .Y(n12700), .A0(n14249), .A1(n13567) );
  nor02 U5833 ( .Y(n12701), .A0(n14224), .A1(n13575) );
  inv01 U5834 ( .Y(n12702), .A(n9780) );
  nor02 U5835 ( .Y(n12699), .A0(n12702), .A1(n12703) );
  nor02 U5836 ( .Y(n12704), .A0(n12700), .A1(n12701) );
  inv01 U5837 ( .Y(n12703), .A(n12704) );
  inv01 U5838 ( .Y(n14142), .A(n12705) );
  nor02 U5839 ( .Y(n12706), .A0(n14234), .A1(n13567) );
  nor02 U5840 ( .Y(n12707), .A0(n14208), .A1(n13575) );
  inv01 U5841 ( .Y(n12708), .A(n9786) );
  nor02 U5842 ( .Y(n12705), .A0(n12708), .A1(n12709) );
  nor02 U5843 ( .Y(n12710), .A0(n12706), .A1(n12707) );
  inv01 U5844 ( .Y(n12709), .A(n12710) );
  inv01 U5845 ( .Y(n14118), .A(n12711) );
  nor02 U5846 ( .Y(n12712), .A0(n14215), .A1(n13567) );
  nor02 U5847 ( .Y(n12713), .A0(n14214), .A1(n13575) );
  inv01 U5848 ( .Y(n12714), .A(n9794) );
  nor02 U5849 ( .Y(n12711), .A0(n12714), .A1(n12715) );
  nor02 U5850 ( .Y(n12716), .A0(n12712), .A1(n12713) );
  inv01 U5851 ( .Y(n12715), .A(n12716) );
  inv02 U5852 ( .Y(n14134), .A(n12717) );
  nor02 U5853 ( .Y(n12718), .A0(n14228), .A1(n13567) );
  nor02 U5854 ( .Y(n12719), .A0(n14227), .A1(n13575) );
  inv01 U5855 ( .Y(n12720), .A(n9798) );
  nor02 U5856 ( .Y(n12717), .A0(n12720), .A1(n12721) );
  nor02 U5857 ( .Y(n12722), .A0(n12718), .A1(n12719) );
  inv01 U5858 ( .Y(n12721), .A(n12722) );
  inv02 U5859 ( .Y(n14182), .A(n12723) );
  nor02 U5860 ( .Y(n12724), .A0(n14313), .A1(n13567) );
  nor02 U5861 ( .Y(n12725), .A0(n14279), .A1(n13575) );
  inv01 U5862 ( .Y(n12726), .A(n9887) );
  nor02 U5863 ( .Y(n12723), .A0(n12726), .A1(n12727) );
  nor02 U5864 ( .Y(n12728), .A0(n12724), .A1(n12725) );
  inv01 U5865 ( .Y(n12727), .A(n12728) );
  inv01 U5866 ( .Y(n14148), .A(n12729) );
  nor02 U5867 ( .Y(n12730), .A0(n14236), .A1(n13567) );
  nor02 U5868 ( .Y(n12731), .A0(n14215), .A1(n13575) );
  inv01 U5869 ( .Y(n12732), .A(n9784) );
  nor02 U5870 ( .Y(n12729), .A0(n12732), .A1(n12733) );
  nor02 U5871 ( .Y(n12734), .A0(n12730), .A1(n12731) );
  inv01 U5872 ( .Y(n12733), .A(n12734) );
  inv02 U5873 ( .Y(n14126), .A(n12735) );
  nor02 U5874 ( .Y(n12736), .A0(n14224), .A1(n13567) );
  nor02 U5875 ( .Y(n12737), .A0(n14223), .A1(n13575) );
  inv01 U5876 ( .Y(n12738), .A(n9802) );
  nor02 U5877 ( .Y(n12735), .A0(n12738), .A1(n12739) );
  nor02 U5878 ( .Y(n12740), .A0(n12736), .A1(n12737) );
  inv01 U5879 ( .Y(n12739), .A(n12740) );
  inv08 U5880 ( .Y(n13567), .A(n13566) );
  nand02 U5881 ( .Y(n14103), .A0(n14143), .A1(n12741) );
  inv01 U5882 ( .Y(n12742), .A(n13745) );
  inv01 U5883 ( .Y(n12743), .A(n13596) );
  inv01 U5884 ( .Y(n12744), .A(n13786) );
  nand02 U5885 ( .Y(n12745), .A0(n9628), .A1(n12742) );
  nand02 U5886 ( .Y(n12746), .A0(n12743), .A1(n12744) );
  nand02 U5887 ( .Y(n12747), .A0(n12745), .A1(n12746) );
  inv01 U5888 ( .Y(n12741), .A(n12747) );
  inv02 U5889 ( .Y(n13831), .A(n12748) );
  nand02 U5890 ( .Y(n12748), .A0(n12749), .A1(n12750) );
  nand02 U5891 ( .Y(n12751), .A0(n10288), .A1(n13941) );
  inv01 U5892 ( .Y(n12749), .A(n12751) );
  nand02 U5893 ( .Y(n12752), .A0(n13782), .A1(n13942) );
  inv01 U5894 ( .Y(n12750), .A(n12752) );
  inv02 U5895 ( .Y(n13942), .A(n12888) );
  buf02 U5896 ( .Y(n12753), .A(n14090) );
  inv02 U5897 ( .Y(n13635), .A(n12754) );
  nand02 U5898 ( .Y(n12754), .A0(n12755), .A1(n12756) );
  nand02 U5899 ( .Y(n12757), .A0(n10292), .A1(n10352) );
  inv01 U5900 ( .Y(n12755), .A(n12757) );
  nand02 U5901 ( .Y(n12758), .A0(n13765), .A1(n13789) );
  inv01 U5902 ( .Y(n12756), .A(n12758) );
  nand02 U5903 ( .Y(n14193), .A0(n12759), .A1(n12760) );
  inv01 U5904 ( .Y(n12761), .A(n13768) );
  inv01 U5905 ( .Y(n12762), .A(n13595) );
  inv01 U5906 ( .Y(n12763), .A(n14342) );
  inv01 U5907 ( .Y(n12764), .A(n13810) );
  nand02 U5908 ( .Y(n12759), .A0(n12761), .A1(n12762) );
  nand02 U5909 ( .Y(n12760), .A0(n12763), .A1(n12764) );
  inv01 U5910 ( .Y(n14342), .A(n14109) );
  nand02 U5911 ( .Y(n14093), .A0(n10063), .A1(n12765) );
  inv01 U5912 ( .Y(n12766), .A(n13583) );
  inv01 U5913 ( .Y(n12767), .A(n13754) );
  inv01 U5914 ( .Y(n12768), .A(n13599) );
  inv01 U5915 ( .Y(n12769), .A(n13807) );
  nand02 U5916 ( .Y(n12770), .A0(n12766), .A1(n12767) );
  nand02 U5917 ( .Y(n12771), .A0(n12768), .A1(n12769) );
  nand02 U5918 ( .Y(n12772), .A0(n12770), .A1(n12771) );
  inv01 U5919 ( .Y(n12765), .A(n12772) );
  inv02 U5920 ( .Y(s_exp_10a_6_), .A(n10507) );
  inv01 U5921 ( .Y(n12773), .A(s_exp_10a_8_) );
  inv02 U5922 ( .Y(n12774), .A(n12773) );
  nand02 U5923 ( .Y(n14285), .A0(n10069), .A1(n12775) );
  inv01 U5924 ( .Y(n12776), .A(n13583) );
  inv01 U5925 ( .Y(n12777), .A(n13745) );
  inv01 U5926 ( .Y(n12778), .A(n13599) );
  inv01 U5927 ( .Y(n12779), .A(n13791) );
  nand02 U5928 ( .Y(n12780), .A0(n12776), .A1(n12777) );
  nand02 U5929 ( .Y(n12781), .A0(n12778), .A1(n12779) );
  nand02 U5930 ( .Y(n12782), .A0(n12780), .A1(n12781) );
  inv01 U5931 ( .Y(n12775), .A(n12782) );
  inv02 U5932 ( .Y(n13791), .A(s_fract_48_i[40]) );
  inv01 U5933 ( .Y(n14276), .A(n12783) );
  nor02 U5934 ( .Y(n12784), .A0(n13792), .A1(n13583) );
  nor02 U5935 ( .Y(n12785), .A0(n13930), .A1(n13599) );
  inv01 U5936 ( .Y(n12786), .A(n9680) );
  nor02 U5937 ( .Y(n12783), .A0(n12786), .A1(n12787) );
  nor02 U5938 ( .Y(n12788), .A0(n12784), .A1(n12785) );
  inv01 U5939 ( .Y(n12787), .A(n12788) );
  inv01 U5940 ( .Y(n14245), .A(n12789) );
  nor02 U5941 ( .Y(n12790), .A0(n13791), .A1(n13583) );
  nor02 U5942 ( .Y(n12791), .A0(n13772), .A1(n13599) );
  inv01 U5943 ( .Y(n12792), .A(n9690) );
  nor02 U5944 ( .Y(n12789), .A0(n12792), .A1(n12793) );
  nor02 U5945 ( .Y(n12794), .A0(n12790), .A1(n12791) );
  inv01 U5946 ( .Y(n12793), .A(n12794) );
  or02 U5947 ( .Y(n12795), .A0(s_fract_48_i[45]), .A1(s_fract_48_i[46]) );
  inv02 U5948 ( .Y(n12796), .A(n12795) );
  buf02 U5949 ( .Y(n12797), .A(n14057) );
  inv02 U5950 ( .Y(n12798), .A(n12848) );
  nand02 U5951 ( .Y(n14345), .A0(n10083), .A1(n12799) );
  inv01 U5952 ( .Y(n12800), .A(n13583) );
  inv01 U5953 ( .Y(n12801), .A(n13785) );
  inv01 U5954 ( .Y(n12802), .A(n13599) );
  inv01 U5955 ( .Y(n12803), .A(n13786) );
  nand02 U5956 ( .Y(n12804), .A0(n12800), .A1(n12801) );
  nand02 U5957 ( .Y(n12805), .A0(n12802), .A1(n12803) );
  nand02 U5958 ( .Y(n12806), .A0(n12804), .A1(n12805) );
  inv01 U5959 ( .Y(n12799), .A(n12806) );
  inv02 U5960 ( .Y(n13786), .A(n10396) );
  inv01 U5961 ( .Y(n12807), .A(s_exp_10a_7_) );
  inv02 U5962 ( .Y(n12808), .A(n12807) );
  buf02 U5963 ( .Y(n12809), .A(n14067) );
  inv02 U5964 ( .Y(n13976), .A(n12810) );
  inv01 U5965 ( .Y(n12811), .A(n13520) );
  nor02 U5966 ( .Y(n12812), .A0(s_expo1[5]), .A1(n12811) );
  nor02 U5967 ( .Y(n12813), .A0(n13520), .A1(n____return6651_5_) );
  nor02 U5968 ( .Y(n12810), .A0(n12812), .A1(n12813) );
  inv02 U5969 ( .Y(n13978), .A(n12814) );
  inv01 U5970 ( .Y(n12815), .A(s_frac2a_46_) );
  nor02 U5971 ( .Y(n12816), .A0(s_expo1[4]), .A1(n12815) );
  nor02 U5972 ( .Y(n12817), .A0(s_frac2a_46_), .A1(n____return6651_4_) );
  nor02 U5973 ( .Y(n12814), .A0(n12816), .A1(n12817) );
  inv02 U5974 ( .Y(n13974), .A(n12818) );
  inv01 U5975 ( .Y(n12819), .A(n13520) );
  nor02 U5976 ( .Y(n12820), .A0(s_expo1[6]), .A1(n12819) );
  nor02 U5977 ( .Y(n12821), .A0(n13520), .A1(n____return6651_6_) );
  nor02 U5978 ( .Y(n12818), .A0(n12820), .A1(n12821) );
  inv02 U5979 ( .Y(n13969), .A(n12822) );
  inv01 U5980 ( .Y(n12823), .A(s_frac2a_46_) );
  nor02 U5981 ( .Y(n12824), .A0(s_expo1[7]), .A1(n12823) );
  nor02 U5982 ( .Y(n12825), .A0(s_frac2a_46_), .A1(n____return6651_7_) );
  nor02 U5983 ( .Y(n12822), .A0(n12824), .A1(n12825) );
  buf02 U5984 ( .Y(n12826), .A(n13983) );
  buf02 U5985 ( .Y(n12827), .A(n14200) );
  buf02 U5986 ( .Y(n12828), .A(n14200) );
  inv02 U5987 ( .Y(n13657), .A(n12829) );
  nand02 U5988 ( .Y(n12829), .A0(s_fract_48_i[30]), .A1(n12830) );
  nand02 U5989 ( .Y(n12831), .A0(n13502), .A1(n12919) );
  inv01 U5990 ( .Y(n12830), .A(n12831) );
  inv02 U5991 ( .Y(s_expo2b[0]), .A(n12826) );
  ao221 U5992 ( .Y(n12832), .A0(n14256), .A1(n13566), .B0(n14267), .B1(n13574), 
        .C0(n14347) );
  inv01 U5993 ( .Y(n12833), .A(n12832) );
  ao221 U5994 ( .Y(n12834), .A0(n14250), .A1(n13574), .B0(n14240), .B1(n13566), 
        .C0(n14341) );
  inv01 U5995 ( .Y(n12835), .A(n12834) );
  nand02 U5996 ( .Y(n14371), .A0(n12836), .A1(n12837) );
  inv01 U5997 ( .Y(n12838), .A(s_shr2_5_) );
  inv01 U5998 ( .Y(n12839), .A(n14367) );
  inv01 U5999 ( .Y(n12840), .A(n13592) );
  nand02 U6000 ( .Y(n12836), .A0(n12838), .A1(n12839) );
  nand02 U6001 ( .Y(n12837), .A0(n12838), .A1(n12840) );
  or02 U6002 ( .Y(n12841), .A0(n10375), .A1(s_fract_48_i[4]) );
  inv02 U6003 ( .Y(n12842), .A(n12841) );
  buf02 U6004 ( .Y(n12843), .A(n14386) );
  buf02 U6005 ( .Y(n12844), .A(n14386) );
  nand02 U6006 ( .Y(n14233), .A0(n12845), .A1(n12846) );
  inv02 U6007 ( .Y(n12847), .A(n13566) );
  inv02 U6008 ( .Y(n12848), .A(n14209) );
  inv02 U6009 ( .Y(n12849), .A(n13574) );
  inv02 U6010 ( .Y(n12850), .A(n14280) );
  inv02 U6011 ( .Y(n12851), .A(n14158) );
  inv02 U6012 ( .Y(n12852), .A(n14269) );
  nand02 U6013 ( .Y(n12853), .A0(n12849), .A1(n12854) );
  nand02 U6014 ( .Y(n12855), .A0(n12850), .A1(n12856) );
  nand02 U6015 ( .Y(n12857), .A0(n12851), .A1(n12858) );
  nand02 U6016 ( .Y(n12859), .A0(n12851), .A1(n12860) );
  nand02 U6017 ( .Y(n12861), .A0(n12852), .A1(n12862) );
  nand02 U6018 ( .Y(n12863), .A0(n12852), .A1(n12864) );
  nand02 U6019 ( .Y(n12865), .A0(n12852), .A1(n12866) );
  nand02 U6020 ( .Y(n12867), .A0(n12852), .A1(n12868) );
  nand02 U6021 ( .Y(n12869), .A0(n12847), .A1(n12848) );
  inv01 U6022 ( .Y(n12854), .A(n12869) );
  nand02 U6023 ( .Y(n12870), .A0(n12847), .A1(n12848) );
  inv01 U6024 ( .Y(n12856), .A(n12870) );
  nand02 U6025 ( .Y(n12871), .A0(n12847), .A1(n12849) );
  inv01 U6026 ( .Y(n12858), .A(n12871) );
  nand02 U6027 ( .Y(n12872), .A0(n12847), .A1(n12850) );
  inv01 U6028 ( .Y(n12860), .A(n12872) );
  nand02 U6029 ( .Y(n12873), .A0(n12848), .A1(n12849) );
  inv01 U6030 ( .Y(n12862), .A(n12873) );
  nand02 U6031 ( .Y(n12874), .A0(n12848), .A1(n12850) );
  inv01 U6032 ( .Y(n12864), .A(n12874) );
  nand02 U6033 ( .Y(n12875), .A0(n12849), .A1(n12851) );
  inv01 U6034 ( .Y(n12866), .A(n12875) );
  nand02 U6035 ( .Y(n12876), .A0(n12850), .A1(n12851) );
  inv01 U6036 ( .Y(n12868), .A(n12876) );
  nand02 U6037 ( .Y(n12877), .A0(n12853), .A1(n12855) );
  inv01 U6038 ( .Y(n12878), .A(n12877) );
  nand02 U6039 ( .Y(n12879), .A0(n12857), .A1(n12859) );
  inv01 U6040 ( .Y(n12880), .A(n12879) );
  nand02 U6041 ( .Y(n12881), .A0(n12878), .A1(n12880) );
  inv01 U6042 ( .Y(n12845), .A(n12881) );
  nand02 U6043 ( .Y(n12882), .A0(n12861), .A1(n12863) );
  inv01 U6044 ( .Y(n12883), .A(n12882) );
  nand02 U6045 ( .Y(n12884), .A0(n12865), .A1(n12867) );
  inv01 U6046 ( .Y(n12885), .A(n12884) );
  nand02 U6047 ( .Y(n12886), .A0(n12883), .A1(n12885) );
  inv01 U6048 ( .Y(n12846), .A(n12886) );
  buf02 U6049 ( .Y(n12887), .A(s_fract_48_i[9]) );
  buf02 U6050 ( .Y(n12889), .A(s_fract_48_i[9]) );
  buf02 U6051 ( .Y(n12888), .A(s_fract_48_i[9]) );
  ao221 U6052 ( .Y(n12890), .A0(n14247), .A1(n13576), .B0(n14248), .B1(n13557), 
        .C0(n14337) );
  inv02 U6053 ( .Y(n12891), .A(n12890) );
  nand02 U6054 ( .Y(n14068), .A0(n12892), .A1(n12893) );
  inv02 U6055 ( .Y(n12894), .A(n14262) );
  inv01 U6056 ( .Y(n12895), .A(n13557) );
  inv01 U6057 ( .Y(n12896), .A(n13576) );
  inv01 U6058 ( .Y(n12897), .A(n14259) );
  inv01 U6059 ( .Y(n12898), .A(n14261) );
  nand02 U6060 ( .Y(n12899), .A0(n12896), .A1(n12900) );
  nand02 U6061 ( .Y(n12901), .A0(n12897), .A1(n12902) );
  nand02 U6062 ( .Y(n12903), .A0(n12898), .A1(n12904) );
  nand02 U6063 ( .Y(n12905), .A0(n12898), .A1(n12906) );
  nand02 U6064 ( .Y(n12907), .A0(n12894), .A1(n12895) );
  inv01 U6065 ( .Y(n12900), .A(n12907) );
  nand02 U6066 ( .Y(n12908), .A0(n12894), .A1(n12895) );
  inv01 U6067 ( .Y(n12902), .A(n12908) );
  nand02 U6068 ( .Y(n12909), .A0(n12894), .A1(n12896) );
  inv01 U6069 ( .Y(n12904), .A(n12909) );
  nand02 U6070 ( .Y(n12910), .A0(n12894), .A1(n12897) );
  inv01 U6071 ( .Y(n12906), .A(n12910) );
  nand02 U6072 ( .Y(n12911), .A0(n12899), .A1(n12901) );
  inv01 U6073 ( .Y(n12892), .A(n12911) );
  nand02 U6074 ( .Y(n12912), .A0(n12903), .A1(n12905) );
  inv01 U6075 ( .Y(n12893), .A(n12912) );
  ao221 U6076 ( .Y(n12913), .A0(n14289), .A1(n13576), .B0(n14324), .B1(n13557), 
        .C0(n14362) );
  inv02 U6077 ( .Y(n12914), .A(n12913) );
  buf08 U6078 ( .Y(n13557), .A(n14246) );
  inv02 U6079 ( .Y(s_expo2b[3]), .A(n9905) );
  buf08 U6080 ( .Y(n12915), .A(n13980) );
  inv02 U6081 ( .Y(n13973), .A(n12915) );
  ao221 U6082 ( .Y(n12916), .A0(n14277), .A1(n13576), .B0(n14278), .B1(n13557), 
        .C0(n14355) );
  inv02 U6083 ( .Y(n12917), .A(n12916) );
  nand02 U6084 ( .Y(n12918), .A0(n13952), .A1(n9632) );
  inv02 U6085 ( .Y(n12919), .A(n12918) );
  or02 U6086 ( .Y(n12920), .A0(n13563), .A1(n13577) );
  inv02 U6087 ( .Y(n12921), .A(n12920) );
  buf02 U6088 ( .Y(n12922), .A(s_fract_48_i[8]) );
  buf02 U6089 ( .Y(n12925), .A(s_fract_48_i[8]) );
  buf02 U6090 ( .Y(n12923), .A(s_fract_48_i[8]) );
  buf02 U6091 ( .Y(n12924), .A(s_fract_48_i[8]) );
  or02 U6092 ( .Y(n12926), .A0(n12267), .A1(n13577) );
  inv02 U6093 ( .Y(n12927), .A(n12926) );
  inv02 U6094 ( .Y(n13938), .A(n12928) );
  inv01 U6095 ( .Y(n12929), .A(n13746) );
  inv01 U6096 ( .Y(n12930), .A(n13785) );
  inv01 U6097 ( .Y(n12931), .A(n13786) );
  inv01 U6098 ( .Y(n12932), .A(n12796) );
  nor02 U6099 ( .Y(n12928), .A0(n12933), .A1(n12934) );
  nor02 U6100 ( .Y(n12935), .A0(n12929), .A1(n12930) );
  inv01 U6101 ( .Y(n12933), .A(n12935) );
  nor02 U6102 ( .Y(n12936), .A0(n12931), .A1(n12932) );
  inv01 U6103 ( .Y(n12934), .A(n12936) );
  inv02 U6104 ( .Y(n14324), .A(n12937) );
  nor02 U6105 ( .Y(n12938), .A0(n13796), .A1(n13583) );
  nor02 U6106 ( .Y(n12939), .A0(n13794), .A1(n13599) );
  inv01 U6107 ( .Y(n12940), .A(n9949) );
  nor02 U6108 ( .Y(n12937), .A0(n12940), .A1(n12941) );
  nor02 U6109 ( .Y(n12942), .A0(n12938), .A1(n12939) );
  inv01 U6110 ( .Y(n12941), .A(n12942) );
  inv02 U6111 ( .Y(n14261), .A(n12943) );
  nor02 U6112 ( .Y(n12944), .A0(n13797), .A1(n13582) );
  nor02 U6113 ( .Y(n12945), .A0(n13798), .A1(n13598) );
  inv01 U6114 ( .Y(n12946), .A(n9676) );
  nor02 U6115 ( .Y(n12943), .A0(n12946), .A1(n12947) );
  nor02 U6116 ( .Y(n12948), .A0(n12944), .A1(n12945) );
  inv01 U6117 ( .Y(n12947), .A(n12948) );
  inv02 U6118 ( .Y(n14286), .A(n14324) );
  inv02 U6119 ( .Y(n14302), .A(n14261) );
  inv02 U6120 ( .Y(n14194), .A(n12949) );
  nor02 U6121 ( .Y(n12950), .A0(n13749), .A1(n13580) );
  nor02 U6122 ( .Y(n12951), .A0(n13784), .A1(n13596) );
  inv01 U6123 ( .Y(n12952), .A(n10065) );
  nor02 U6124 ( .Y(n12949), .A0(n12952), .A1(n12953) );
  nor02 U6125 ( .Y(n12954), .A0(n12950), .A1(n12951) );
  inv01 U6126 ( .Y(n12953), .A(n12954) );
  inv02 U6127 ( .Y(n14189), .A(n12955) );
  nor02 U6128 ( .Y(n12956), .A0(n13784), .A1(n13580) );
  nor02 U6129 ( .Y(n12957), .A0(n13937), .A1(n13595) );
  inv01 U6130 ( .Y(n12958), .A(n9708) );
  nor02 U6131 ( .Y(n12955), .A0(n12958), .A1(n12959) );
  nor02 U6132 ( .Y(n12960), .A0(n12956), .A1(n12957) );
  inv01 U6133 ( .Y(n12959), .A(n12960) );
  inv02 U6134 ( .Y(n14183), .A(n12961) );
  nor02 U6135 ( .Y(n12962), .A0(n13937), .A1(n13580) );
  nor02 U6136 ( .Y(n12963), .A0(n13800), .A1(n13596) );
  inv01 U6137 ( .Y(n12964), .A(n9742) );
  nor02 U6138 ( .Y(n12961), .A0(n12964), .A1(n12965) );
  nor02 U6139 ( .Y(n12966), .A0(n12962), .A1(n12963) );
  inv01 U6140 ( .Y(n12965), .A(n12966) );
  inv02 U6141 ( .Y(n14249), .A(n14194) );
  inv02 U6142 ( .Y(n13784), .A(n12418) );
  inv02 U6143 ( .Y(n14236), .A(n14189) );
  inv02 U6144 ( .Y(n13937), .A(n10724) );
  inv02 U6145 ( .Y(n14234), .A(n14183) );
  inv02 U6146 ( .Y(n14203), .A(n12967) );
  nor02 U6147 ( .Y(n12968), .A0(n13801), .A1(n13580) );
  nor02 U6148 ( .Y(n12969), .A0(n13749), .A1(n13595) );
  inv01 U6149 ( .Y(n12970), .A(n14305) );
  nor02 U6150 ( .Y(n12967), .A0(n12970), .A1(n12971) );
  nor02 U6151 ( .Y(n12972), .A0(n12968), .A1(n12969) );
  inv01 U6152 ( .Y(n12971), .A(n12972) );
  inv02 U6153 ( .Y(n14266), .A(n14203) );
  inv02 U6154 ( .Y(n14229), .A(n12973) );
  nor02 U6155 ( .Y(n12974), .A0(n13804), .A1(n13580) );
  nor02 U6156 ( .Y(n12975), .A0(n13803), .A1(n13595) );
  inv01 U6157 ( .Y(n12976), .A(n9684) );
  nor02 U6158 ( .Y(n12973), .A0(n12976), .A1(n12977) );
  nor02 U6159 ( .Y(n12978), .A0(n12974), .A1(n12975) );
  inv01 U6160 ( .Y(n12977), .A(n12978) );
  inv02 U6161 ( .Y(n14288), .A(n12979) );
  nor02 U6162 ( .Y(n12980), .A0(n13930), .A1(n13582) );
  nor02 U6163 ( .Y(n12981), .A0(n13790), .A1(n13598) );
  inv01 U6164 ( .Y(n12982), .A(n14363) );
  nor02 U6165 ( .Y(n12979), .A0(n12982), .A1(n12983) );
  nor02 U6166 ( .Y(n12984), .A0(n12980), .A1(n12981) );
  inv01 U6167 ( .Y(n12983), .A(n12984) );
  inv02 U6168 ( .Y(n14304), .A(n14229) );
  inv02 U6169 ( .Y(n14225), .A(n12985) );
  nor02 U6170 ( .Y(n12986), .A0(n13803), .A1(n13580) );
  nor02 U6171 ( .Y(n12987), .A0(n13779), .A1(n13596) );
  inv01 U6172 ( .Y(n12988), .A(n10031) );
  nor02 U6173 ( .Y(n12985), .A0(n12988), .A1(n12989) );
  nor02 U6174 ( .Y(n12990), .A0(n12986), .A1(n12987) );
  inv01 U6175 ( .Y(n12989), .A(n12990) );
  inv02 U6176 ( .Y(n14211), .A(n12991) );
  nor02 U6177 ( .Y(n12992), .A0(n13802), .A1(n13580) );
  nor02 U6178 ( .Y(n12993), .A0(n13801), .A1(n13596) );
  inv01 U6179 ( .Y(n12994), .A(n14314) );
  nor02 U6180 ( .Y(n12991), .A0(n12994), .A1(n12995) );
  nor02 U6181 ( .Y(n12996), .A0(n12992), .A1(n12993) );
  inv01 U6182 ( .Y(n12995), .A(n12996) );
  inv02 U6183 ( .Y(n14216), .A(n12997) );
  nor02 U6184 ( .Y(n12998), .A0(n13779), .A1(n13580) );
  nor02 U6185 ( .Y(n12999), .A0(n13802), .A1(n13595) );
  inv01 U6186 ( .Y(n13000), .A(n9963) );
  nor02 U6187 ( .Y(n12997), .A0(n13000), .A1(n13001) );
  nor02 U6188 ( .Y(n13002), .A0(n12998), .A1(n12999) );
  inv01 U6189 ( .Y(n13001), .A(n13002) );
  inv02 U6190 ( .Y(n14297), .A(n14225) );
  inv02 U6191 ( .Y(n14279), .A(n14211) );
  inv02 U6192 ( .Y(n14290), .A(n14216) );
  inv02 U6193 ( .Y(n14318), .A(n13003) );
  nor02 U6194 ( .Y(n13004), .A0(n14104), .A1(n13582) );
  nor02 U6195 ( .Y(n13005), .A0(n13747), .A1(n13598) );
  inv01 U6196 ( .Y(n13006), .A(n9638) );
  nor02 U6197 ( .Y(n13003), .A0(n13006), .A1(n13007) );
  nor02 U6198 ( .Y(n13008), .A0(n13004), .A1(n13005) );
  inv01 U6199 ( .Y(n13007), .A(n13008) );
  or02 U6200 ( .Y(n13009), .A0(n14340), .A1(n13769) );
  inv02 U6201 ( .Y(n13010), .A(n13009) );
  inv02 U6202 ( .Y(n14169), .A(n13011) );
  nor02 U6203 ( .Y(n13012), .A0(n13767), .A1(n13580) );
  nor02 U6204 ( .Y(n13013), .A0(n13927), .A1(n13596) );
  inv01 U6205 ( .Y(n13014), .A(n9710) );
  nor02 U6206 ( .Y(n13011), .A0(n13014), .A1(n13015) );
  nor02 U6207 ( .Y(n13016), .A0(n13012), .A1(n13013) );
  inv01 U6208 ( .Y(n13015), .A(n13016) );
  inv02 U6209 ( .Y(n14176), .A(n13017) );
  nor02 U6210 ( .Y(n13018), .A0(n13799), .A1(n13580) );
  nor02 U6211 ( .Y(n13019), .A0(n13766), .A1(n13596) );
  inv01 U6212 ( .Y(n13020), .A(n14251) );
  nor02 U6213 ( .Y(n13017), .A0(n13020), .A1(n13021) );
  nor02 U6214 ( .Y(n13022), .A0(n13018), .A1(n13019) );
  inv01 U6215 ( .Y(n13021), .A(n13022) );
  inv02 U6216 ( .Y(n14208), .A(n14169) );
  inv02 U6217 ( .Y(n14224), .A(n14176) );
  inv02 U6218 ( .Y(n14316), .A(n13023) );
  nor02 U6219 ( .Y(n13024), .A0(n13927), .A1(n13582) );
  nor02 U6220 ( .Y(n13025), .A0(n13767), .A1(n13598) );
  inv01 U6221 ( .Y(n13026), .A(n10001) );
  nor02 U6222 ( .Y(n13023), .A0(n13026), .A1(n13027) );
  nor02 U6223 ( .Y(n13028), .A0(n13024), .A1(n13025) );
  inv01 U6224 ( .Y(n13027), .A(n13028) );
  inv02 U6225 ( .Y(n14296), .A(n13029) );
  nor02 U6226 ( .Y(n13030), .A0(n13789), .A1(n13582) );
  nor02 U6227 ( .Y(n13031), .A0(n13765), .A1(n13598) );
  inv01 U6228 ( .Y(n13032), .A(n9682) );
  nor02 U6229 ( .Y(n13029), .A0(n13032), .A1(n13033) );
  nor02 U6230 ( .Y(n13034), .A0(n13030), .A1(n13031) );
  inv01 U6231 ( .Y(n13033), .A(n13034) );
  inv02 U6232 ( .Y(n14173), .A(n13035) );
  nor02 U6233 ( .Y(n13036), .A0(n13766), .A1(n13580) );
  nor02 U6234 ( .Y(n13037), .A0(n13767), .A1(n13595) );
  inv01 U6235 ( .Y(n13038), .A(n9983) );
  nor02 U6236 ( .Y(n13035), .A0(n13038), .A1(n13039) );
  nor02 U6237 ( .Y(n13040), .A0(n13036), .A1(n13037) );
  inv01 U6238 ( .Y(n13039), .A(n13040) );
  inv02 U6239 ( .Y(n14180), .A(n13041) );
  nor02 U6240 ( .Y(n13042), .A0(n13800), .A1(n13580) );
  nor02 U6241 ( .Y(n13043), .A0(n13799), .A1(n13595) );
  inv01 U6242 ( .Y(n13044), .A(n9670) );
  nor02 U6243 ( .Y(n13041), .A0(n13044), .A1(n13045) );
  nor02 U6244 ( .Y(n13046), .A0(n13042), .A1(n13043) );
  inv01 U6245 ( .Y(n13045), .A(n13046) );
  inv02 U6246 ( .Y(n14275), .A(n14316) );
  inv02 U6247 ( .Y(n13927), .A(n12349) );
  inv02 U6248 ( .Y(n14243), .A(n14296) );
  inv02 U6249 ( .Y(n14215), .A(n14173) );
  inv02 U6250 ( .Y(n13767), .A(n12409) );
  inv02 U6251 ( .Y(n14228), .A(n14180) );
  inv02 U6252 ( .Y(n14064), .A(n13047) );
  nor02 U6253 ( .Y(n13048), .A0(n13799), .A1(n13582) );
  nor02 U6254 ( .Y(n13049), .A0(n13800), .A1(n13598) );
  inv01 U6255 ( .Y(n13050), .A(n9692) );
  nor02 U6256 ( .Y(n13047), .A0(n13050), .A1(n13051) );
  nor02 U6257 ( .Y(n13052), .A0(n13048), .A1(n13049) );
  inv01 U6258 ( .Y(n13051), .A(n13052) );
  inv02 U6259 ( .Y(n13957), .A(n13961) );
  inv02 U6260 ( .Y(n14303), .A(n14064) );
  inv02 U6261 ( .Y(n13800), .A(s_fract_48_i[22]) );
  inv02 U6262 ( .Y(n13799), .A(s_fract_48_i[23]) );
  inv02 U6263 ( .Y(n14059), .A(n13053) );
  nor02 U6264 ( .Y(n13054), .A0(n14239), .A1(n13575) );
  nor02 U6265 ( .Y(n13055), .A0(n13423), .A1(n13567) );
  nor02 U6266 ( .Y(n13056), .A0(n13393), .A1(n14199) );
  nor02 U6267 ( .Y(n13053), .A0(n13056), .A1(n13057) );
  nor02 U6268 ( .Y(n13058), .A0(n13054), .A1(n13055) );
  inv01 U6269 ( .Y(n13057), .A(n13058) );
  inv02 U6270 ( .Y(n14077), .A(n13059) );
  nor02 U6271 ( .Y(n13060), .A0(n14273), .A1(n13558) );
  nor02 U6272 ( .Y(n13061), .A0(n14272), .A1(n13577) );
  nor02 U6273 ( .Y(n13062), .A0(n13562), .A1(n14271) );
  nor02 U6274 ( .Y(n13059), .A0(n13062), .A1(n13063) );
  nor02 U6275 ( .Y(n13064), .A0(n13060), .A1(n13061) );
  inv01 U6276 ( .Y(n13063), .A(n13064) );
  inv02 U6277 ( .Y(n14050), .A(n13065) );
  nor02 U6278 ( .Y(n13066), .A0(n13766), .A1(n13583) );
  nor02 U6279 ( .Y(n13067), .A0(n13799), .A1(n13599) );
  inv01 U6280 ( .Y(n13068), .A(n9642) );
  nor02 U6281 ( .Y(n13065), .A0(n13068), .A1(n13069) );
  nor02 U6282 ( .Y(n13070), .A0(n13066), .A1(n13067) );
  inv01 U6283 ( .Y(n13069), .A(n13070) );
  inv02 U6284 ( .Y(n14069), .A(n13071) );
  nor02 U6285 ( .Y(n13072), .A0(n14199), .A1(n14255) );
  nor02 U6286 ( .Y(n13073), .A0(n14254), .A1(n13567) );
  nor02 U6287 ( .Y(n13074), .A0(n14253), .A1(n13575) );
  nor02 U6288 ( .Y(n13071), .A0(n13074), .A1(n13075) );
  nor02 U6289 ( .Y(n13076), .A0(n13072), .A1(n13073) );
  inv01 U6290 ( .Y(n13075), .A(n13076) );
  inv02 U6291 ( .Y(n14165), .A(n13077) );
  nor02 U6292 ( .Y(n13078), .A0(n14272), .A1(n13558) );
  nor02 U6293 ( .Y(n13079), .A0(n14317), .A1(n13577) );
  inv01 U6294 ( .Y(n13080), .A(n9873) );
  nor02 U6295 ( .Y(n13077), .A0(n13080), .A1(n13081) );
  nor02 U6296 ( .Y(n13082), .A0(n13078), .A1(n13079) );
  inv01 U6297 ( .Y(n13081), .A(n13082) );
  inv02 U6298 ( .Y(n14294), .A(n14050) );
  inv02 U6299 ( .Y(n13766), .A(n12460) );
  inv02 U6300 ( .Y(n14317), .A(n14276) );
  inv02 U6301 ( .Y(n14272), .A(n14356) );
  inv02 U6302 ( .Y(n14325), .A(n13083) );
  nor02 U6303 ( .Y(n13084), .A0(n13767), .A1(n13583) );
  nor02 U6304 ( .Y(n13085), .A0(n13766), .A1(n13599) );
  inv01 U6305 ( .Y(n13086), .A(n10029) );
  nor02 U6306 ( .Y(n13083), .A0(n13086), .A1(n13087) );
  nor02 U6307 ( .Y(n13088), .A0(n13084), .A1(n13085) );
  inv01 U6308 ( .Y(n13087), .A(n13088) );
  inv02 U6309 ( .Y(n14287), .A(n14325) );
  inv02 U6310 ( .Y(n14129), .A(n13089) );
  nor02 U6311 ( .Y(n13090), .A0(n13763), .A1(n13580) );
  nor02 U6312 ( .Y(n13091), .A0(n13790), .A1(n13596) );
  inv01 U6313 ( .Y(n13092), .A(n9979) );
  nor02 U6314 ( .Y(n13089), .A0(n13092), .A1(n13093) );
  nor02 U6315 ( .Y(n13094), .A0(n13090), .A1(n13091) );
  inv01 U6316 ( .Y(n13093), .A(n13094) );
  inv02 U6317 ( .Y(n14137), .A(n13095) );
  nor02 U6318 ( .Y(n13096), .A0(n13795), .A1(n13580) );
  nor02 U6319 ( .Y(n13097), .A0(n13763), .A1(n13595) );
  inv01 U6320 ( .Y(n13098), .A(n14179) );
  nor02 U6321 ( .Y(n13095), .A0(n13098), .A1(n13099) );
  nor02 U6322 ( .Y(n13100), .A0(n13096), .A1(n13097) );
  inv01 U6323 ( .Y(n13099), .A(n13100) );
  nand02 U6324 ( .Y(n14121), .A0(n9768), .A1(n13101) );
  inv01 U6325 ( .Y(n13102), .A(n13790) );
  inv01 U6326 ( .Y(n13103), .A(n13595) );
  inv01 U6327 ( .Y(n13104), .A(n13930) );
  nand02 U6328 ( .Y(n13105), .A0(n9629), .A1(n13102) );
  nand02 U6329 ( .Y(n13106), .A0(n13103), .A1(n13104) );
  nand02 U6330 ( .Y(n13107), .A0(n13105), .A1(n13106) );
  inv01 U6331 ( .Y(n13101), .A(n13107) );
  inv02 U6332 ( .Y(n13930), .A(n10830) );
  inv02 U6333 ( .Y(n13790), .A(n12255) );
  inv02 U6334 ( .Y(n14237), .A(n13108) );
  nor02 U6335 ( .Y(n13109), .A0(n13805), .A1(n13580) );
  nor02 U6336 ( .Y(n13110), .A0(n13756), .A1(n13595) );
  inv01 U6337 ( .Y(n13111), .A(n9666) );
  nor02 U6338 ( .Y(n13108), .A0(n13111), .A1(n13112) );
  nor02 U6339 ( .Y(n13113), .A0(n13109), .A1(n13110) );
  inv01 U6340 ( .Y(n13112), .A(n13113) );
  inv02 U6341 ( .Y(n14235), .A(n13114) );
  nor02 U6342 ( .Y(n13115), .A0(n13756), .A1(n13580) );
  nor02 U6343 ( .Y(n13116), .A0(n13804), .A1(n13596) );
  inv01 U6344 ( .Y(n13117), .A(n9716) );
  nor02 U6345 ( .Y(n13114), .A0(n13117), .A1(n13118) );
  nor02 U6346 ( .Y(n13119), .A0(n13115), .A1(n13116) );
  inv01 U6347 ( .Y(n13118), .A(n13119) );
  inv02 U6348 ( .Y(n14117), .A(n13120) );
  nor02 U6349 ( .Y(n13121), .A0(n14319), .A1(n14204) );
  nor02 U6350 ( .Y(n13122), .A0(n14326), .A1(n13575) );
  inv01 U6351 ( .Y(n13123), .A(n9864) );
  nor02 U6352 ( .Y(n13120), .A0(n13123), .A1(n13124) );
  nor02 U6353 ( .Y(n13125), .A0(n13121), .A1(n13122) );
  inv01 U6354 ( .Y(n13124), .A(n13125) );
  inv02 U6355 ( .Y(n14326), .A(n14237) );
  inv02 U6356 ( .Y(n14114), .A(n13126) );
  nor02 U6357 ( .Y(n13127), .A0(n14310), .A1(n14204) );
  nor02 U6358 ( .Y(n13128), .A0(n14313), .A1(n13575) );
  inv01 U6359 ( .Y(n13129), .A(n9875) );
  nor02 U6360 ( .Y(n13126), .A0(n13129), .A1(n13130) );
  nor02 U6361 ( .Y(n13131), .A0(n13127), .A1(n13128) );
  inv01 U6362 ( .Y(n13130), .A(n13131) );
  inv02 U6363 ( .Y(n14313), .A(n14235) );
  inv02 U6364 ( .Y(n14185), .A(n13132) );
  nor02 U6365 ( .Y(n13133), .A0(n14322), .A1(n13558) );
  nor02 U6366 ( .Y(n13134), .A0(n14321), .A1(n13577) );
  inv01 U6367 ( .Y(n13135), .A(n9965) );
  nor02 U6368 ( .Y(n13132), .A0(n13135), .A1(n13136) );
  nor02 U6369 ( .Y(n13137), .A0(n13133), .A1(n13134) );
  inv01 U6370 ( .Y(n13136), .A(n13137) );
  inv02 U6371 ( .Y(n14322), .A(n14285) );
  inv02 U6372 ( .Y(n14099), .A(n13138) );
  nor02 U6373 ( .Y(n13139), .A0(n13930), .A1(n13580) );
  nor02 U6374 ( .Y(n13140), .A0(n13792), .A1(n13596) );
  inv01 U6375 ( .Y(n13141), .A(n9720) );
  nor02 U6376 ( .Y(n13138), .A0(n13141), .A1(n13142) );
  nor02 U6377 ( .Y(n13143), .A0(n13139), .A1(n13140) );
  inv01 U6378 ( .Y(n13142), .A(n13143) );
  inv02 U6379 ( .Y(n14061), .A(n13144) );
  nor02 U6380 ( .Y(n13145), .A0(n13805), .A1(n13582) );
  nor02 U6381 ( .Y(n13146), .A0(n13753), .A1(n13598) );
  inv01 U6382 ( .Y(n13147), .A(n9672) );
  nor02 U6383 ( .Y(n13144), .A0(n13147), .A1(n13148) );
  nor02 U6384 ( .Y(n13149), .A0(n13145), .A1(n13146) );
  inv01 U6385 ( .Y(n13148), .A(n13149) );
  inv02 U6386 ( .Y(n13792), .A(s_fract_48_i[38]) );
  inv02 U6387 ( .Y(n14196), .A(n13150) );
  nor02 U6388 ( .Y(n13151), .A0(n14257), .A1(n14338) );
  nor02 U6389 ( .Y(n13152), .A0(n14258), .A1(n13562) );
  inv01 U6390 ( .Y(n13153), .A(n14368) );
  nor02 U6391 ( .Y(n13150), .A0(n13153), .A1(n13154) );
  nor02 U6392 ( .Y(n13155), .A0(n13151), .A1(n13152) );
  inv01 U6393 ( .Y(n13154), .A(n13155) );
  inv02 U6394 ( .Y(n14191), .A(n13156) );
  nor02 U6395 ( .Y(n13157), .A0(n13417), .A1(n13562) );
  nor02 U6396 ( .Y(n13158), .A0(n14293), .A1(n13558) );
  inv01 U6397 ( .Y(n13159), .A(n9804) );
  nor02 U6398 ( .Y(n13156), .A0(n13159), .A1(n13160) );
  nor02 U6399 ( .Y(n13161), .A0(n13157), .A1(n13158) );
  inv01 U6400 ( .Y(n13160), .A(n13161) );
  inv02 U6401 ( .Y(n14089), .A(n13162) );
  nor02 U6402 ( .Y(n13163), .A0(n14241), .A1(n13562) );
  nor02 U6403 ( .Y(n13164), .A0(n14293), .A1(n13577) );
  nor02 U6404 ( .Y(n13165), .A0(n13417), .A1(n13558) );
  nor02 U6405 ( .Y(n13162), .A0(n13165), .A1(n13166) );
  nor02 U6406 ( .Y(n13167), .A0(n13163), .A1(n13164) );
  inv01 U6407 ( .Y(n13166), .A(n13167) );
  inv02 U6408 ( .Y(n14293), .A(n14245) );
  inv02 U6409 ( .Y(n14265), .A(n13168) );
  nor02 U6410 ( .Y(n13169), .A0(n13772), .A1(n13582) );
  nor02 U6411 ( .Y(n13170), .A0(n13792), .A1(n13598) );
  inv01 U6412 ( .Y(n13171), .A(n9646) );
  nor02 U6413 ( .Y(n13168), .A0(n13171), .A1(n13172) );
  nor02 U6414 ( .Y(n13173), .A0(n13169), .A1(n13170) );
  inv01 U6415 ( .Y(n13172), .A(n13173) );
  inv02 U6416 ( .Y(n14073), .A(n13174) );
  nor02 U6417 ( .Y(n13175), .A0(n13804), .A1(n13583) );
  nor02 U6418 ( .Y(n13176), .A0(n13756), .A1(n13599) );
  inv01 U6419 ( .Y(n13177), .A(n9678) );
  nor02 U6420 ( .Y(n13174), .A0(n13177), .A1(n13178) );
  nor02 U6421 ( .Y(n13179), .A0(n13175), .A1(n13176) );
  inv01 U6422 ( .Y(n13178), .A(n13179) );
  inv02 U6423 ( .Y(n13821), .A(n13180) );
  inv01 U6424 ( .Y(n13181), .A(n13772) );
  inv01 U6425 ( .Y(n13182), .A(n13902) );
  inv01 U6426 ( .Y(n13183), .A(n13938) );
  nand02 U6427 ( .Y(n13180), .A0(n13183), .A1(n13184) );
  nand02 U6428 ( .Y(n13185), .A0(n13181), .A1(n13182) );
  inv01 U6429 ( .Y(n13184), .A(n13185) );
  inv02 U6430 ( .Y(n14065), .A(n13186) );
  nor02 U6431 ( .Y(n13187), .A0(n13753), .A1(n13583) );
  nor02 U6432 ( .Y(n13188), .A0(n13806), .A1(n13599) );
  inv01 U6433 ( .Y(n13189), .A(n9748) );
  nor02 U6434 ( .Y(n13186), .A0(n13189), .A1(n13190) );
  nor02 U6435 ( .Y(n13191), .A0(n13187), .A1(n13188) );
  inv01 U6436 ( .Y(n13190), .A(n13191) );
  inv02 U6437 ( .Y(n13804), .A(s_fract_48_i[14]) );
  inv02 U6438 ( .Y(n14095), .A(n13192) );
  nor02 U6439 ( .Y(n13193), .A0(n14301), .A1(n13577) );
  nor02 U6440 ( .Y(n13194), .A0(n14258), .A1(n13558) );
  nor02 U6441 ( .Y(n13195), .A0(n14257), .A1(n13562) );
  nor02 U6442 ( .Y(n13192), .A0(n13195), .A1(n13196) );
  nor02 U6443 ( .Y(n13197), .A0(n13193), .A1(n13194) );
  inv01 U6444 ( .Y(n13196), .A(n13197) );
  inv02 U6445 ( .Y(n14258), .A(n14345) );
  inv02 U6446 ( .Y(n14301), .A(n14265) );
  inv02 U6447 ( .Y(n14080), .A(n13198) );
  nor02 U6448 ( .Y(n13199), .A0(n13756), .A1(n13582) );
  nor02 U6449 ( .Y(n13200), .A0(n13805), .A1(n13598) );
  inv01 U6450 ( .Y(n13201), .A(n9746) );
  nor02 U6451 ( .Y(n13198), .A0(n13201), .A1(n13202) );
  nor02 U6452 ( .Y(n13203), .A0(n13199), .A1(n13200) );
  inv01 U6453 ( .Y(n13202), .A(n13203) );
  inv02 U6454 ( .Y(n13805), .A(s_fract_48_i[12]) );
  or02 U6455 ( .Y(n13204), .A0(n13715), .A1(n13761) );
  inv02 U6456 ( .Y(n13205), .A(n13204) );
  nand03 U6457 ( .Y(n13206), .A0(n13511), .A1(n13768), .A2(n13770) );
  inv02 U6458 ( .Y(n13207), .A(n13206) );
  nand02 U6459 ( .Y(n13208), .A0(s_fract_48_i[31]), .A1(n13788) );
  inv02 U6460 ( .Y(n13209), .A(n13208) );
  buf02 U6461 ( .Y(n13210), .A(n14311) );
  inv02 U6462 ( .Y(n14353), .A(s_shr2_2_) );
  nor02 U6463 ( .Y(n13211), .A0(n13582), .A1(n14398) );
  inv04 U6464 ( .Y(n14398), .A(s_shr3) );
  inv02 U6465 ( .Y(n14255), .A(n12827) );
  inv02 U6466 ( .Y(n14240), .A(n13212) );
  nor02 U6467 ( .Y(n13213), .A0(n13754), .A1(n13580) );
  nor02 U6468 ( .Y(n13214), .A0(n13782), .A1(n13595) );
  inv01 U6469 ( .Y(n13215), .A(n9738) );
  nor02 U6470 ( .Y(n13212), .A0(n13215), .A1(n13216) );
  nor02 U6471 ( .Y(n13217), .A0(n13213), .A1(n13214) );
  inv01 U6472 ( .Y(n13216), .A(n13217) );
  inv02 U6473 ( .Y(n14248), .A(n13218) );
  nor02 U6474 ( .Y(n13219), .A0(n13790), .A1(n13582) );
  nor02 U6475 ( .Y(n13220), .A0(n13763), .A1(n13598) );
  inv01 U6476 ( .Y(n13221), .A(n10047) );
  nor02 U6477 ( .Y(n13218), .A0(n13221), .A1(n13222) );
  nor02 U6478 ( .Y(n13223), .A0(n13219), .A1(n13220) );
  inv01 U6479 ( .Y(n13222), .A(n13223) );
  inv02 U6480 ( .Y(n14278), .A(n13224) );
  nor02 U6481 ( .Y(n13225), .A0(n13795), .A1(n13582) );
  nor02 U6482 ( .Y(n13226), .A0(n13796), .A1(n13598) );
  inv01 U6483 ( .Y(n13227), .A(n9921) );
  nor02 U6484 ( .Y(n13224), .A0(n13227), .A1(n13228) );
  nor02 U6485 ( .Y(n13229), .A0(n13225), .A1(n13226) );
  inv01 U6486 ( .Y(n13228), .A(n13229) );
  inv02 U6487 ( .Y(n13754), .A(n10287) );
  inv02 U6488 ( .Y(n13763), .A(n10820) );
  inv02 U6489 ( .Y(n14256), .A(n13230) );
  nor02 U6490 ( .Y(n13231), .A0(n13807), .A1(n13580) );
  nor02 U6491 ( .Y(n13232), .A0(n13754), .A1(n13595) );
  inv01 U6492 ( .Y(n13233), .A(n9668) );
  nor02 U6493 ( .Y(n13230), .A0(n13233), .A1(n13234) );
  nor02 U6494 ( .Y(n13235), .A0(n13231), .A1(n13232) );
  inv01 U6495 ( .Y(n13234), .A(n13235) );
  inv02 U6496 ( .Y(n13807), .A(s_fract_48_i[6]) );
  inv02 U6497 ( .Y(n14284), .A(n13236) );
  nor02 U6498 ( .Y(n13237), .A0(n13747), .A1(n13583) );
  nor02 U6499 ( .Y(n13238), .A0(n13746), .A1(n13599) );
  inv01 U6500 ( .Y(n13239), .A(n9686) );
  nor02 U6501 ( .Y(n13236), .A0(n13239), .A1(n13240) );
  nor02 U6502 ( .Y(n13241), .A0(n13237), .A1(n13238) );
  inv01 U6503 ( .Y(n13240), .A(n13241) );
  nor02 U6504 ( .Y(n13243), .A0(n13811), .A1(n13580) );
  nor02 U6505 ( .Y(n13244), .A0(n13917), .A1(n13595) );
  inv01 U6506 ( .Y(n13245), .A(n9898) );
  nor02 U6507 ( .Y(n13242), .A0(n13245), .A1(n13246) );
  nor02 U6508 ( .Y(n13247), .A0(n13243), .A1(n13244) );
  inv02 U6509 ( .Y(n13246), .A(n13247) );
  inv02 U6510 ( .Y(n14132), .A(n13248) );
  nor02 U6511 ( .Y(n13249), .A0(n13769), .A1(n13582) );
  nor02 U6512 ( .Y(n13250), .A0(n14104), .A1(n13598) );
  inv01 U6513 ( .Y(n13251), .A(n10061) );
  nor02 U6514 ( .Y(n13248), .A0(n13251), .A1(n13252) );
  nor02 U6515 ( .Y(n13253), .A0(n13249), .A1(n13250) );
  inv01 U6516 ( .Y(n13252), .A(n13253) );
  inv02 U6517 ( .Y(n14269), .A(n13254) );
  nor02 U6518 ( .Y(n13255), .A0(n13917), .A1(n13580) );
  nor02 U6519 ( .Y(n13256), .A0(n13807), .A1(n13596) );
  inv01 U6520 ( .Y(n13257), .A(n9902) );
  nor02 U6521 ( .Y(n13254), .A0(n13257), .A1(n13258) );
  nor02 U6522 ( .Y(n13259), .A0(n13255), .A1(n13256) );
  inv01 U6523 ( .Y(n13258), .A(n13259) );
  inv02 U6524 ( .Y(n14257), .A(n14132) );
  inv02 U6525 ( .Y(n14104), .A(s_fract_48_i[46]) );
  inv02 U6526 ( .Y(n13917), .A(n10376) );
  inv02 U6527 ( .Y(n14150), .A(n13260) );
  nor02 U6528 ( .Y(n13261), .A0(n13789), .A1(n13580) );
  nor02 U6529 ( .Y(n13262), .A0(n13928), .A1(n13595) );
  inv01 U6530 ( .Y(n13263), .A(n9652) );
  nor02 U6531 ( .Y(n13260), .A0(n13263), .A1(n13264) );
  nor02 U6532 ( .Y(n13265), .A0(n13261), .A1(n13262) );
  inv01 U6533 ( .Y(n13264), .A(n13265) );
  inv02 U6534 ( .Y(n14153), .A(n13266) );
  nor02 U6535 ( .Y(n13267), .A0(n13765), .A1(n13580) );
  nor02 U6536 ( .Y(n13268), .A0(n13789), .A1(n13596) );
  inv01 U6537 ( .Y(n13269), .A(n9674) );
  nor02 U6538 ( .Y(n13266), .A0(n13269), .A1(n13270) );
  nor02 U6539 ( .Y(n13271), .A0(n13267), .A1(n13268) );
  inv01 U6540 ( .Y(n13270), .A(n13271) );
  inv02 U6541 ( .Y(n14156), .A(n13272) );
  nor02 U6542 ( .Y(n13273), .A0(n13927), .A1(n13580) );
  nor02 U6543 ( .Y(n13274), .A0(n13765), .A1(n13595) );
  inv01 U6544 ( .Y(n13275), .A(n9722) );
  nor02 U6545 ( .Y(n13272), .A0(n13275), .A1(n13276) );
  nor02 U6546 ( .Y(n13277), .A0(n13273), .A1(n13274) );
  inv01 U6547 ( .Y(n13276), .A(n13277) );
  inv02 U6548 ( .Y(n14144), .A(n13278) );
  nor02 U6549 ( .Y(n13279), .A0(n13928), .A1(n13580) );
  nor02 U6550 ( .Y(n13280), .A0(n13798), .A1(n13596) );
  inv01 U6551 ( .Y(n13281), .A(n9718) );
  nor02 U6552 ( .Y(n13278), .A0(n13281), .A1(n13282) );
  nor02 U6553 ( .Y(n13283), .A0(n13279), .A1(n13280) );
  inv01 U6554 ( .Y(n13282), .A(n13283) );
  inv02 U6555 ( .Y(n13928), .A(n10291) );
  inv02 U6556 ( .Y(n13789), .A(n12251) );
  inv02 U6557 ( .Y(n13765), .A(n10573) );
  inv02 U6558 ( .Y(n14291), .A(n13284) );
  nor02 U6559 ( .Y(n13285), .A0(n13782), .A1(n13580) );
  nor02 U6560 ( .Y(n13286), .A0(n13942), .A1(n13596) );
  inv01 U6561 ( .Y(n13287), .A(n9648) );
  nor02 U6562 ( .Y(n13284), .A0(n13287), .A1(n13288) );
  nor02 U6563 ( .Y(n13289), .A0(n13285), .A1(n13286) );
  inv01 U6564 ( .Y(n13288), .A(n13289) );
  inv02 U6565 ( .Y(n14267), .A(n13290) );
  nor02 U6566 ( .Y(n13291), .A0(n13806), .A1(n13580) );
  nor02 U6567 ( .Y(n13292), .A0(n13753), .A1(n13596) );
  inv01 U6568 ( .Y(n13293), .A(n9752) );
  nor02 U6569 ( .Y(n13290), .A0(n13293), .A1(n13294) );
  nor02 U6570 ( .Y(n13295), .A0(n13291), .A1(n13292) );
  inv01 U6571 ( .Y(n13294), .A(n13295) );
  inv02 U6572 ( .Y(n14280), .A(n13296) );
  nor02 U6573 ( .Y(n13297), .A0(n13942), .A1(n13580) );
  nor02 U6574 ( .Y(n13298), .A0(n13806), .A1(n13596) );
  inv01 U6575 ( .Y(n13299), .A(n9750) );
  nor02 U6576 ( .Y(n13296), .A0(n13299), .A1(n13300) );
  nor02 U6577 ( .Y(n13301), .A0(n13297), .A1(n13298) );
  inv01 U6578 ( .Y(n13300), .A(n13301) );
  inv02 U6579 ( .Y(n13806), .A(s_fract_48_i[10]) );
  inv02 U6580 ( .Y(n14247), .A(n13302) );
  nor02 U6581 ( .Y(n13303), .A0(n13794), .A1(n13583) );
  nor02 U6582 ( .Y(n13304), .A0(n13797), .A1(n13599) );
  inv01 U6583 ( .Y(n13305), .A(n9660) );
  nor02 U6584 ( .Y(n13302), .A0(n13305), .A1(n13306) );
  nor02 U6585 ( .Y(n13307), .A0(n13303), .A1(n13304) );
  inv01 U6586 ( .Y(n13306), .A(n13307) );
  inv02 U6587 ( .Y(n14250), .A(n13308) );
  nor02 U6588 ( .Y(n13309), .A0(n13753), .A1(n13580) );
  nor02 U6589 ( .Y(n13310), .A0(n13805), .A1(n13596) );
  inv01 U6590 ( .Y(n13311), .A(n9724) );
  nor02 U6591 ( .Y(n13308), .A0(n13311), .A1(n13312) );
  nor02 U6592 ( .Y(n13313), .A0(n13309), .A1(n13310) );
  inv01 U6593 ( .Y(n13312), .A(n13313) );
  inv02 U6594 ( .Y(n14289), .A(n13314) );
  nor02 U6595 ( .Y(n13315), .A0(n13928), .A1(n13582) );
  nor02 U6596 ( .Y(n13316), .A0(n13789), .A1(n13598) );
  inv01 U6597 ( .Y(n13317), .A(n9688) );
  nor02 U6598 ( .Y(n13314), .A0(n13317), .A1(n13318) );
  nor02 U6599 ( .Y(n13319), .A0(n13315), .A1(n13316) );
  inv01 U6600 ( .Y(n13318), .A(n13319) );
  inv02 U6601 ( .Y(n14277), .A(n13320) );
  nor02 U6602 ( .Y(n13321), .A0(n13798), .A1(n13583) );
  nor02 U6603 ( .Y(n13322), .A0(n13928), .A1(n13599) );
  inv01 U6604 ( .Y(n13323), .A(n9712) );
  nor02 U6605 ( .Y(n13320), .A0(n13323), .A1(n13324) );
  nor02 U6606 ( .Y(n13325), .A0(n13321), .A1(n13322) );
  inv01 U6607 ( .Y(n13324), .A(n13325) );
  inv02 U6608 ( .Y(n13798), .A(s_fract_48_i[30]) );
  inv02 U6609 ( .Y(n14264), .A(n13326) );
  nor02 U6610 ( .Y(n13327), .A0(n13763), .A1(n13583) );
  nor02 U6611 ( .Y(n13328), .A0(n13795), .A1(n13599) );
  inv01 U6612 ( .Y(n13329), .A(n9664) );
  nor02 U6613 ( .Y(n13326), .A0(n13329), .A1(n13330) );
  nor02 U6614 ( .Y(n13331), .A0(n13327), .A1(n13328) );
  inv01 U6615 ( .Y(n13330), .A(n13331) );
  inv02 U6616 ( .Y(n14081), .A(n13332) );
  nor02 U6617 ( .Y(n13333), .A0(n13937), .A1(n13582) );
  nor02 U6618 ( .Y(n13334), .A0(n13784), .A1(n13598) );
  inv01 U6619 ( .Y(n13335), .A(n10033) );
  nor02 U6620 ( .Y(n13332), .A0(n13335), .A1(n13336) );
  nor02 U6621 ( .Y(n13337), .A0(n13333), .A1(n13334) );
  inv01 U6622 ( .Y(n13336), .A(n13337) );
  inv02 U6623 ( .Y(n14070), .A(n13338) );
  nor02 U6624 ( .Y(n13339), .A0(n13749), .A1(n13583) );
  nor02 U6625 ( .Y(n13340), .A0(n13801), .A1(n13599) );
  inv01 U6626 ( .Y(n13341), .A(n9654) );
  nor02 U6627 ( .Y(n13338), .A0(n13341), .A1(n13342) );
  nor02 U6628 ( .Y(n13343), .A0(n13339), .A1(n13340) );
  inv01 U6629 ( .Y(n13342), .A(n13343) );
  inv02 U6630 ( .Y(n13795), .A(s_fract_48_i[34]) );
  inv02 U6631 ( .Y(n13801), .A(s_fract_48_i[18]) );
  inv02 U6632 ( .Y(n13749), .A(n10720) );
  inv02 U6633 ( .Y(n14138), .A(n13344) );
  nor02 U6634 ( .Y(n13345), .A0(n13798), .A1(n13580) );
  nor02 U6635 ( .Y(n13346), .A0(n13797), .A1(n13595) );
  inv01 U6636 ( .Y(n13347), .A(n9640) );
  nor02 U6637 ( .Y(n13344), .A0(n13347), .A1(n13348) );
  nor02 U6638 ( .Y(n13349), .A0(n13345), .A1(n13346) );
  inv01 U6639 ( .Y(n13348), .A(n13349) );
  inv02 U6640 ( .Y(n14122), .A(n13350) );
  nor02 U6641 ( .Y(n13351), .A0(n13794), .A1(n13580) );
  nor02 U6642 ( .Y(n13352), .A0(n13796), .A1(n13595) );
  inv01 U6643 ( .Y(n13353), .A(n14188) );
  nor02 U6644 ( .Y(n13350), .A0(n13353), .A1(n13354) );
  nor02 U6645 ( .Y(n13355), .A0(n13351), .A1(n13352) );
  inv01 U6646 ( .Y(n13354), .A(n13355) );
  inv02 U6647 ( .Y(n14130), .A(n13356) );
  nor02 U6648 ( .Y(n13357), .A0(n13797), .A1(n13580) );
  nor02 U6649 ( .Y(n13358), .A0(n13794), .A1(n13596) );
  inv01 U6650 ( .Y(n13359), .A(n9947) );
  nor02 U6651 ( .Y(n13356), .A0(n13359), .A1(n13360) );
  nor02 U6652 ( .Y(n13361), .A0(n13357), .A1(n13358) );
  inv01 U6653 ( .Y(n13360), .A(n13361) );
  inv02 U6654 ( .Y(n13796), .A(s_fract_48_i[33]) );
  inv02 U6655 ( .Y(n13797), .A(s_fract_48_i[31]) );
  inv02 U6656 ( .Y(n14072), .A(n13362) );
  nor02 U6657 ( .Y(n13363), .A0(n13800), .A1(n13583) );
  nor02 U6658 ( .Y(n13364), .A0(n13937), .A1(n13599) );
  inv01 U6659 ( .Y(n13365), .A(n9650) );
  nor02 U6660 ( .Y(n13362), .A0(n13365), .A1(n13366) );
  nor02 U6661 ( .Y(n13367), .A0(n13363), .A1(n13364) );
  inv01 U6662 ( .Y(n13366), .A(n13367) );
  inv02 U6663 ( .Y(n14259), .A(n13368) );
  nor02 U6664 ( .Y(n13369), .A0(n13765), .A1(n13583) );
  nor02 U6665 ( .Y(n13370), .A0(n13927), .A1(n13599) );
  inv01 U6666 ( .Y(n13371), .A(n9714) );
  nor02 U6667 ( .Y(n13368), .A0(n13371), .A1(n13372) );
  nor02 U6668 ( .Y(n13373), .A0(n13369), .A1(n13370) );
  inv01 U6669 ( .Y(n13372), .A(n13373) );
  inv02 U6670 ( .Y(n14054), .A(n13374) );
  nor02 U6671 ( .Y(n13375), .A0(n13784), .A1(n13583) );
  nor02 U6672 ( .Y(n13376), .A0(n13749), .A1(n13599) );
  inv01 U6673 ( .Y(n13377), .A(n9997) );
  nor02 U6674 ( .Y(n13374), .A0(n13377), .A1(n13378) );
  nor02 U6675 ( .Y(n13379), .A0(n13375), .A1(n13376) );
  inv01 U6676 ( .Y(n13378), .A(n13379) );
  inv02 U6677 ( .Y(n14112), .A(n13380) );
  nor02 U6678 ( .Y(n13381), .A0(n13796), .A1(n13580) );
  nor02 U6679 ( .Y(n13382), .A0(n13795), .A1(n13596) );
  inv01 U6680 ( .Y(n13383), .A(n9694) );
  nor02 U6681 ( .Y(n13380), .A0(n13383), .A1(n13384) );
  nor02 U6682 ( .Y(n13385), .A0(n13381), .A1(n13382) );
  inv01 U6683 ( .Y(n13384), .A(n13385) );
  inv02 U6684 ( .Y(n14063), .A(n13386) );
  nor02 U6685 ( .Y(n13387), .A0(n13803), .A1(n13582) );
  nor02 U6686 ( .Y(n13388), .A0(n13804), .A1(n13598) );
  inv01 U6687 ( .Y(n13389), .A(n9740) );
  nor02 U6688 ( .Y(n13386), .A0(n13389), .A1(n13390) );
  nor02 U6689 ( .Y(n13391), .A0(n13387), .A1(n13388) );
  inv01 U6690 ( .Y(n13390), .A(n13391) );
  inv02 U6691 ( .Y(n13803), .A(s_fract_48_i[15]) );
  buf02 U6692 ( .Y(n13392), .A(n14193) );
  inv02 U6693 ( .Y(n13393), .A(n13392) );
  inv02 U6694 ( .Y(n13394), .A(n13392) );
  inv02 U6695 ( .Y(n14254), .A(n14348) );
  inv02 U6696 ( .Y(n14052), .A(n13395) );
  nor02 U6697 ( .Y(n13396), .A0(n13779), .A1(n13582) );
  nor02 U6698 ( .Y(n13397), .A0(n13803), .A1(n13598) );
  inv01 U6699 ( .Y(n13398), .A(n9658) );
  nor02 U6700 ( .Y(n13395), .A0(n13398), .A1(n13399) );
  nor02 U6701 ( .Y(n13400), .A0(n13396), .A1(n13397) );
  inv01 U6702 ( .Y(n13399), .A(n13400) );
  nor02 U6703 ( .Y(n13402), .A0(n13801), .A1(n13583) );
  nor02 U6704 ( .Y(n13403), .A0(n13802), .A1(n13599) );
  inv01 U6705 ( .Y(n13404), .A(n14351) );
  nor02 U6706 ( .Y(n13401), .A0(n13404), .A1(n13405) );
  nor02 U6707 ( .Y(n13406), .A0(n13402), .A1(n13403) );
  inv01 U6708 ( .Y(n13405), .A(n13406) );
  inv02 U6709 ( .Y(n14082), .A(n13407) );
  nor02 U6710 ( .Y(n13408), .A0(n13802), .A1(n13582) );
  nor02 U6711 ( .Y(n13409), .A0(n13779), .A1(n13598) );
  inv01 U6712 ( .Y(n13410), .A(n14358) );
  nor02 U6713 ( .Y(n13407), .A0(n13410), .A1(n13411) );
  nor02 U6714 ( .Y(n13412), .A0(n13408), .A1(n13409) );
  inv01 U6715 ( .Y(n13411), .A(n13412) );
  inv02 U6716 ( .Y(n13802), .A(s_fract_48_i[17]) );
  inv02 U6717 ( .Y(n13941), .A(n13413) );
  nand02 U6718 ( .Y(n13413), .A0(n10421), .A1(n13414) );
  nand02 U6719 ( .Y(n13415), .A0(n13806), .A1(n13753) );
  inv01 U6720 ( .Y(n13414), .A(n13415) );
  buf02 U6721 ( .Y(n13416), .A(n14339) );
  inv02 U6722 ( .Y(n13417), .A(n13416) );
  inv02 U6723 ( .Y(n13418), .A(n13416) );
  inv02 U6724 ( .Y(n13419), .A(n13762) );
  inv02 U6725 ( .Y(n13420), .A(n13419) );
  inv02 U6726 ( .Y(n13421), .A(n13419) );
  buf02 U6727 ( .Y(n13422), .A(n14343) );
  inv02 U6728 ( .Y(n13423), .A(n13422) );
  or02 U6729 ( .Y(n13424), .A0(s_fract_48_i[1]), .A1(s_fract_48_i[0]) );
  inv02 U6730 ( .Y(n13425), .A(n13424) );
  inv02 U6731 ( .Y(n13426), .A(n13748) );
  inv02 U6732 ( .Y(n13427), .A(n13426) );
  inv02 U6733 ( .Y(n13428), .A(n13426) );
  inv02 U6734 ( .Y(n13429), .A(n13936) );
  inv02 U6735 ( .Y(n13430), .A(n13429) );
  inv02 U6736 ( .Y(n13431), .A(n13429) );
  nand02 U6737 ( .Y(n13432), .A0(n12445), .A1(n13792) );
  inv02 U6738 ( .Y(n13433), .A(n13432) );
  inv02 U6739 ( .Y(n14387), .A(n13434) );
  inv01 U6740 ( .Y(n13435), .A(n14391) );
  inv01 U6741 ( .Y(n13436), .A(n12220) );
  inv01 U6742 ( .Y(n13437), .A(n14389) );
  nand02 U6743 ( .Y(n13434), .A0(n13437), .A1(n13438) );
  nand02 U6744 ( .Y(n13439), .A0(n13435), .A1(n13436) );
  inv01 U6745 ( .Y(n13438), .A(n13439) );
  inv02 U6746 ( .Y(n14391), .A(s_exp_10_i_3_) );
  inv02 U6747 ( .Y(n13752), .A(n13440) );
  nand02 U6748 ( .Y(n13440), .A0(n13205), .A1(n13441) );
  nand02 U6749 ( .Y(n13442), .A0(n13425), .A1(n13807) );
  inv01 U6750 ( .Y(n13441), .A(n13442) );
  xor2 U6751 ( .Y(n13443), .A0(n14388), .A1(s_exp_10_i_5_) );
  inv04 U6752 ( .Y(n13444), .A(n9774) );
  xor2 U6753 ( .Y(n13445), .A0(n13769), .A1(s_exp_10_i_0_) );
  inv02 U6754 ( .Y(n13446), .A(n13445) );
  inv01 U6755 ( .Y(n13447), .A(n13445) );
  inv02 U6756 ( .Y(n14158), .A(n13448) );
  nor02 U6757 ( .Y(n13449), .A0(n13810), .A1(n13580) );
  nor02 U6758 ( .Y(n13450), .A0(n14308), .A1(n13595) );
  inv01 U6759 ( .Y(n13451), .A(n9904) );
  nor02 U6760 ( .Y(n13448), .A0(n13451), .A1(n13452) );
  nor02 U6761 ( .Y(n13453), .A0(n13449), .A1(n13450) );
  inv01 U6762 ( .Y(n13452), .A(n13453) );
  inv02 U6763 ( .Y(n14310), .A(n14158) );
  inv02 U6764 ( .Y(n14308), .A(s_fract_48_i[2]) );
  inv02 U6765 ( .Y(n13810), .A(s_fract_48_i[1]) );
  xor2 U6766 ( .Y(n13454), .A0(n12220), .A1(s_exp_10_i_2_) );
  inv01 U6767 ( .Y(n13455), .A(n13454) );
  inv02 U6768 ( .Y(n13456), .A(n13454) );
  xor2 U6769 ( .Y(n13457), .A0(n14391), .A1(n10329) );
  inv01 U6770 ( .Y(n13458), .A(n13457) );
  inv02 U6771 ( .Y(n13459), .A(n13457) );
  xor2 U6772 ( .Y(n13460), .A0(n14392), .A1(s_exp_10_i_1_) );
  inv01 U6773 ( .Y(n13461), .A(n13460) );
  inv02 U6774 ( .Y(n13462), .A(n13460) );
  inv02 U6775 ( .Y(n14187), .A(n13463) );
  nor02 U6776 ( .Y(n13464), .A0(n14308), .A1(n14342) );
  nor02 U6777 ( .Y(n13465), .A0(n13810), .A1(n13595) );
  nor02 U6778 ( .Y(n13466), .A0(n13580), .A1(n13768) );
  nor02 U6779 ( .Y(n13463), .A0(n13466), .A1(n13467) );
  nor02 U6780 ( .Y(n13468), .A0(n13464), .A1(n13465) );
  inv01 U6781 ( .Y(n13467), .A(n13468) );
  inv02 U6782 ( .Y(n14319), .A(n14187) );
  inv02 U6783 ( .Y(n13768), .A(s_fract_48_i[0]) );
  inv02 U6784 ( .Y(n13469), .A(n13968) );
  inv02 U6785 ( .Y(n13470), .A(n13469) );
  inv02 U6786 ( .Y(n13471), .A(n13469) );
  inv02 U6787 ( .Y(n13472), .A(n13967) );
  inv02 U6788 ( .Y(n13473), .A(n13472) );
  inv02 U6789 ( .Y(n13474), .A(n13472) );
  inv02 U6790 ( .Y(n14124), .A(n13476) );
  nor02 U6791 ( .Y(n13477), .A0(n13769), .A1(n13598) );
  nor02 U6792 ( .Y(n13478), .A0(n13747), .A1(n14340) );
  nor02 U6793 ( .Y(n13479), .A0(n14104), .A1(n13518) );
  nor02 U6794 ( .Y(n13476), .A0(n13479), .A1(n13480) );
  nor02 U6795 ( .Y(n13481), .A0(n13477), .A1(n13478) );
  inv01 U6796 ( .Y(n13480), .A(n13481) );
  inv02 U6797 ( .Y(n14241), .A(n14124) );
  inv02 U6798 ( .Y(n13751), .A(n13482) );
  inv01 U6799 ( .Y(n13483), .A(n10286) );
  inv01 U6800 ( .Y(n13484), .A(n12887) );
  inv01 U6801 ( .Y(n13485), .A(n12925) );
  nand02 U6802 ( .Y(n13482), .A0(n13485), .A1(n13486) );
  nand02 U6803 ( .Y(n13487), .A0(n13483), .A1(n13484) );
  inv01 U6804 ( .Y(n13486), .A(n13487) );
  inv02 U6805 ( .Y(n13770), .A(n13488) );
  nand02 U6806 ( .Y(n13488), .A0(n13916), .A1(n13489) );
  nand02 U6807 ( .Y(n13490), .A0(n13205), .A1(n13810) );
  inv01 U6808 ( .Y(n13489), .A(n13490) );
  inv08 U6809 ( .Y(n13564), .A(n13563) );
  inv02 U6810 ( .Y(n13916), .A(n13515) );
  inv02 U6811 ( .Y(n13750), .A(n13491) );
  inv01 U6812 ( .Y(n13492), .A(n10722) );
  inv01 U6813 ( .Y(n13493), .A(n10726) );
  inv01 U6814 ( .Y(n13494), .A(n12417) );
  nand02 U6815 ( .Y(n13491), .A0(n13494), .A1(n13495) );
  nand02 U6816 ( .Y(n13496), .A0(n13492), .A1(n13493) );
  inv01 U6817 ( .Y(n13495), .A(n13496) );
  inv02 U6818 ( .Y(n14116), .A(n13497) );
  nor02 U6819 ( .Y(n13498), .A0(n14104), .A1(n14340) );
  nor02 U6820 ( .Y(n13499), .A0(n13769), .A1(n13518) );
  nor02 U6821 ( .Y(n13497), .A0(n13498), .A1(n13499) );
  inv02 U6822 ( .Y(n14340), .A(n13592) );
  nand02 U6823 ( .Y(n13501), .A0(n13778), .A1(n13799) );
  inv02 U6824 ( .Y(n13502), .A(n13501) );
  inv02 U6825 ( .Y(n13771), .A(n13503) );
  inv01 U6826 ( .Y(n13504), .A(n10821) );
  inv01 U6827 ( .Y(n13505), .A(n10829) );
  inv01 U6828 ( .Y(n13506), .A(n12254) );
  nand02 U6829 ( .Y(n13503), .A0(n13506), .A1(n13507) );
  nand02 U6830 ( .Y(n13508), .A0(n13504), .A1(n13505) );
  inv01 U6831 ( .Y(n13507), .A(n13508) );
  nand02 U6832 ( .Y(n13509), .A0(n13929), .A1(n13798) );
  inv04 U6833 ( .Y(n13510), .A(n13509) );
  buf02 U6834 ( .Y(n13511), .A(s_fract_48_i[47]) );
  buf02 U6835 ( .Y(n13514), .A(s_fract_48_i[47]) );
  buf02 U6836 ( .Y(n13512), .A(s_fract_48_i[47]) );
  buf02 U6837 ( .Y(n13513), .A(s_fract_48_i[47]) );
  nand02 U6838 ( .Y(n13515), .A0(n13941), .A1(n13516) );
  nand02 U6839 ( .Y(n13517), .A0(n13751), .A1(n13807) );
  inv01 U6840 ( .Y(n13516), .A(n13517) );
  inv04 U6841 ( .Y(n13520), .A(n13519) );
  inv02 U6842 ( .Y(n14375), .A(n13521) );
  inv01 U6843 ( .Y(n13522), .A(n14376) );
  inv01 U6844 ( .Y(n13523), .A(n13537) );
  inv01 U6845 ( .Y(n13524), .A(n13617) );
  nand02 U6846 ( .Y(n13521), .A0(n13524), .A1(n13525) );
  nand02 U6847 ( .Y(n13526), .A0(n13522), .A1(n13523) );
  inv01 U6848 ( .Y(n13525), .A(n13526) );
  inv04 U6849 ( .Y(n13794), .A(n10883) );
  inv04 U6850 ( .Y(n13779), .A(n10569) );
  inv04 U6851 ( .Y(n13769), .A(n13512) );
  inv04 U6852 ( .Y(n13785), .A(s_fract_48_i[43]) );
  inv04 U6853 ( .Y(n13756), .A(n10502) );
  buf04 U6854 ( .Y(n13561), .A(n14263) );
  buf08 U6855 ( .Y(n13576), .A(n14260) );
  inv04 U6856 ( .Y(n13745), .A(s_fract_48_i[41]) );
  inv04 U6857 ( .Y(n13966), .A(n13528) );
  inv01 U6858 ( .Y(n13529), .A(n13617) );
  inv01 U6859 ( .Y(n13530), .A(s_exp_10b[8]) );
  inv01 U6860 ( .Y(n13531), .A(n13537) );
  nand02 U6861 ( .Y(n13528), .A0(n13531), .A1(n13532) );
  nand02 U6862 ( .Y(n13533), .A0(n13529), .A1(n13530) );
  inv01 U6863 ( .Y(n13532), .A(n13533) );
  buf08 U6864 ( .Y(n13566), .A(n14270) );
  buf02 U6865 ( .Y(n13534), .A(n13746) );
  inv04 U6866 ( .Y(n13746), .A(s_fract_48_i[44]) );
  buf02 U6867 ( .Y(n13536), .A(n14113) );
  inv04 U6868 ( .Y(n13537), .A(n13616) );
  inv02 U6869 ( .Y(n13616), .A(n13956) );
  inv02 U6870 ( .Y(n13538), .A(n14060) );
  inv02 U6871 ( .Y(n13539), .A(n13538) );
  buf08 U6872 ( .Y(n13542), .A(n14210) );
  buf02 U6873 ( .Y(n13543), .A(n14111) );
  buf02 U6874 ( .Y(n13544), .A(n14111) );
  inv02 U6875 ( .Y(n13546), .A(n14053) );
  inv02 U6876 ( .Y(n13550), .A(n14098) );
  inv02 U6877 ( .Y(n14338), .A(n13556) );
  inv08 U6878 ( .Y(n13560), .A(n14199) );
  inv08 U6879 ( .Y(n13562), .A(n13561) );
  inv04 U6880 ( .Y(n14199), .A(n12798) );
  buf16 U6881 ( .Y(n13565), .A(n14058) );
  inv08 U6882 ( .Y(n13569), .A(n13568) );
  inv08 U6883 ( .Y(n13570), .A(n13972) );
  inv08 U6884 ( .Y(n13571), .A(n13970) );
  inv12 U6885 ( .Y(n13575), .A(n13574) );
  inv12 U6886 ( .Y(n13577), .A(n13576) );
  buf16 U6887 ( .Y(n13578), .A(n10368) );
  buf12 U6888 ( .Y(n13579), .A(n14163) );
  nand02 U6889 ( .Y(n13581), .A0(s_shr2_1_), .A1(s_shr2_0_) );
  buf16 U6890 ( .Y(n13582), .A(n14161) );
  buf16 U6891 ( .Y(n13583), .A(n13581) );
  nor02 U6892 ( .Y(n13584), .A0(s_shl2_1_), .A1(s_shl2_0_) );
  nor02 U6893 ( .Y(n13585), .A0(s_shl2_1_), .A1(s_shl2_0_) );
  inv04 U6894 ( .Y(n13586), .A(n13589) );
  inv02 U6895 ( .Y(n13587), .A(n13584) );
  inv04 U6896 ( .Y(n13588), .A(n13587) );
  inv02 U6897 ( .Y(n13589), .A(n13585) );
  inv04 U6898 ( .Y(n13590), .A(n13589) );
  inv02 U6899 ( .Y(n13591), .A(n14162) );
  inv12 U6900 ( .Y(n13592), .A(n10162) );
  buf12 U6901 ( .Y(n13593), .A(n14108) );
  or02 U6902 ( .Y(n13594), .A0(n14360), .A1(s_shl2_1_) );
  buf16 U6903 ( .Y(n13595), .A(n14105) );
  buf12 U6904 ( .Y(n13596), .A(n13594) );
  or02 U6905 ( .Y(n13597), .A0(n14399), .A1(s_shr2_0_) );
  buf16 U6906 ( .Y(n13598), .A(n14160) );
  buf12 U6907 ( .Y(n13599), .A(n13597) );
  inv01 U6908 ( .Y(n13725), .A(n13624) );
  inv01 U6909 ( .Y(n13724), .A(n13626) );
  nor02 U6910 ( .Y(n13723), .A0(n12470), .A1(n13628) );
  inv01 U6911 ( .Y(n13722), .A(n13629) );
  inv01 U6912 ( .Y(n13734), .A(n13207) );
  nor02 U6913 ( .Y(n13733), .A0(n13209), .A1(n13633) );
  nor02 U6914 ( .Y(n13732), .A0(n13639), .A1(n13638) );
  inv01 U6915 ( .Y(n13731), .A(n13640) );
  nor02 U6916 ( .Y(n13742), .A0(n13644), .A1(n10331) );
  nor02 U6917 ( .Y(n13741), .A0(n13645), .A1(n10363) );
  inv01 U6918 ( .Y(n13740), .A(n10273) );
  inv01 U6919 ( .Y(n13739), .A(n13649) );
  nor02 U6920 ( .Y(n13760), .A0(n13657), .A1(n13655) );
  inv01 U6921 ( .Y(n13759), .A(n13658) );
  inv01 U6922 ( .Y(n13758), .A(n13659) );
  inv01 U6923 ( .Y(n13702), .A(n13622) );
  inv01 U6924 ( .Y(n13701), .A(n12470) );
  inv01 U6925 ( .Y(n13700), .A(n13629) );
  nand03 U6926 ( .Y(n13698), .A0(n13705), .A1(n13706), .A2(n13704) );
  inv01 U6927 ( .Y(n13706), .A(n13207) );
  nor02 U6928 ( .Y(n13705), .A0(n13209), .A1(n13636) );
  nor02 U6929 ( .Y(n13704), .A0(n13639), .A1(n13635) );
  nand03 U6930 ( .Y(n13697), .A0(n13708), .A1(n13709), .A2(n13707) );
  nor02 U6931 ( .Y(n13709), .A0(n13644), .A1(n13662) );
  nor02 U6932 ( .Y(n13708), .A0(n10363), .A1(n13643) );
  nor02 U6933 ( .Y(n13707), .A0(n10273), .A1(n13648) );
  and02 U6934 ( .Y(n13600), .A0(n13715), .A1(n13425) );
  nor02 U6935 ( .Y(n13712), .A0(n13657), .A1(n13653) );
  inv01 U6936 ( .Y(n13711), .A(n13656) );
  inv01 U6937 ( .Y(n13710), .A(n13659) );
  nand03 U6938 ( .Y(n13680), .A0(n13682), .A1(n13683), .A2(n13681) );
  inv01 U6939 ( .Y(n13683), .A(n13622) );
  nor02 U6940 ( .Y(n13682), .A0(n13625), .A1(n13626) );
  nor02 U6941 ( .Y(n13681), .A0(n13629), .A1(n13630) );
  inv01 U6942 ( .Y(n13687), .A(n13207) );
  nor02 U6943 ( .Y(n13686), .A0(n13635), .A1(n13209) );
  nor02 U6944 ( .Y(n13685), .A0(n13637), .A1(n13638) );
  nor02 U6945 ( .Y(n13684), .A0(n13640), .A1(n13641) );
  inv01 U6946 ( .Y(n13691), .A(n13644) );
  nor02 U6947 ( .Y(n13690), .A0(n13645), .A1(n13646) );
  nor02 U6948 ( .Y(n13689), .A0(n13648), .A1(n10273) );
  inv01 U6949 ( .Y(n13688), .A(n13650) );
  nand03 U6950 ( .Y(n13677), .A0(n13693), .A1(n13694), .A2(n13692) );
  inv01 U6951 ( .Y(n13693), .A(n13661) );
  nor02 U6952 ( .Y(n13692), .A0(n10331), .A1(n13662) );
  nand03 U6953 ( .Y(n13666), .A0(n10356), .A1(n13668), .A2(n13667) );
  inv01 U6954 ( .Y(n13668), .A(n13623) );
  inv01 U6955 ( .Y(n13667), .A(n13630) );
  nand02 U6956 ( .Y(n13665), .A0(n13669), .A1(n13670) );
  nor02 U6957 ( .Y(n13670), .A0(n13635), .A1(n13209) );
  inv01 U6958 ( .Y(n13669), .A(n13638) );
  nand03 U6959 ( .Y(n13664), .A0(n13672), .A1(n13673), .A2(n13671) );
  nor02 U6960 ( .Y(n13673), .A0(n13643), .A1(n10363) );
  inv01 U6961 ( .Y(n13672), .A(n13647) );
  nor02 U6962 ( .Y(n13671), .A0(n13649), .A1(n13650) );
  nand02 U6963 ( .Y(n13663), .A0(n13674), .A1(n13675) );
  inv01 U6964 ( .Y(n13674), .A(n13660) );
  nor02 U6965 ( .Y(n13632), .A0(n13637), .A1(n13639) );
  nor02 U6966 ( .Y(n13631), .A0(n13640), .A1(n13641) );
  inv01 U6967 ( .Y(n13620), .A(n13642) );
  inv01 U6968 ( .Y(n13642), .A(n13644) );
  nand03 U6969 ( .Y(n13619), .A0(n13652), .A1(n10365), .A2(n13651) );
  nor02 U6970 ( .Y(n13651), .A0(n13662), .A1(n10331) );
  nand03 U6971 ( .Y(n13907), .A0(n13909), .A1(n13910), .A2(n13908) );
  nor02 U6972 ( .Y(n13910), .A0(n13816), .A1(n13817) );
  nor02 U6973 ( .Y(n13909), .A0(n10158), .A1(n13821) );
  inv01 U6974 ( .Y(n13908), .A(n13824) );
  nor02 U6975 ( .Y(n13915), .A0(n13828), .A1(n10367) );
  nor02 U6976 ( .Y(n13914), .A0(n13830), .A1(n13829) );
  inv01 U6977 ( .Y(n13913), .A(n13831) );
  inv01 U6978 ( .Y(n13912), .A(n13835) );
  nor02 U6979 ( .Y(n13925), .A0(n13840), .A1(n10399) );
  inv01 U6980 ( .Y(n13924), .A(n13841) );
  inv01 U6981 ( .Y(n13923), .A(n13843) );
  inv01 U6982 ( .Y(n13922), .A(n13770) );
  nand03 U6983 ( .Y(n13904), .A0(n13933), .A1(n13934), .A2(n13932) );
  inv01 U6984 ( .Y(n13933), .A(n13847) );
  nor02 U6985 ( .Y(n13932), .A0(n10390), .A1(n13851) );
  nor02 U6986 ( .Y(n13892), .A0(n13816), .A1(n10279) );
  inv01 U6987 ( .Y(n13891), .A(n13818) );
  inv01 U6988 ( .Y(n13890), .A(n13821) );
  inv01 U6989 ( .Y(n13896), .A(n12422) );
  nor02 U6990 ( .Y(n13894), .A0(n13831), .A1(n13833) );
  inv01 U6991 ( .Y(n13893), .A(n13835) );
  nand03 U6992 ( .Y(n13887), .A0(n13898), .A1(n10373), .A2(n13897) );
  inv01 U6993 ( .Y(n13898), .A(n13844) );
  nor02 U6994 ( .Y(n13897), .A0(n13770), .A1(n10301) );
  nand03 U6995 ( .Y(n13886), .A0(n13900), .A1(n10200), .A2(n13899) );
  and04 U6996 ( .Y(n13601), .A0(n10395), .A1(n12796), .A2(n13785), .A3(n13746)
         );
  nor02 U6997 ( .Y(n13900), .A0(n13849), .A1(n13847) );
  nor02 U6998 ( .Y(n13899), .A0(n10390), .A1(n13853) );
  inv01 U6999 ( .Y(n13876), .A(n13816) );
  inv01 U7000 ( .Y(n13875), .A(n13818) );
  nor02 U7001 ( .Y(n13874), .A0(n13820), .A1(n13822) );
  nand03 U7002 ( .Y(n13872), .A0(n13878), .A1(n13879), .A2(n13877) );
  nor02 U7003 ( .Y(n13879), .A0(n13827), .A1(n12422) );
  nor02 U7004 ( .Y(n13878), .A0(n13829), .A1(n13830) );
  inv01 U7005 ( .Y(n13877), .A(n13834) );
  inv01 U7006 ( .Y(n13882), .A(n13840) );
  inv01 U7007 ( .Y(n13881), .A(n13842) );
  nor02 U7008 ( .Y(n13880), .A0(n10301), .A1(n10367) );
  nand03 U7009 ( .Y(n13870), .A0(n13884), .A1(n12452), .A2(n13883) );
  inv01 U7010 ( .Y(n13884), .A(n13852) );
  inv01 U7011 ( .Y(n13883), .A(n13855) );
  nand02 U7012 ( .Y(n13860), .A0(n13861), .A1(n13862) );
  nor02 U7013 ( .Y(n13862), .A0(n13817), .A1(n10279) );
  inv01 U7014 ( .Y(n13861), .A(n13819) );
  nand03 U7015 ( .Y(n13859), .A0(n13864), .A1(n13865), .A2(n13863) );
  nor02 U7016 ( .Y(n13865), .A0(n13827), .A1(n12422) );
  nor02 U7017 ( .Y(n13864), .A0(n13829), .A1(n13830) );
  inv01 U7018 ( .Y(n13863), .A(n13835) );
  nand02 U7019 ( .Y(n13858), .A0(n13866), .A1(n13867) );
  nor02 U7020 ( .Y(n13867), .A0(n13838), .A1(n13839) );
  inv01 U7021 ( .Y(n13866), .A(n13841) );
  nand02 U7022 ( .Y(n13857), .A0(n13868), .A1(n12452) );
  nor02 U7023 ( .Y(n13868), .A0(n13855), .A1(n10399) );
  inv01 U7024 ( .Y(n13815), .A(n10386) );
  nand03 U7025 ( .Y(n13814), .A0(n10354), .A1(n13826), .A2(n13825) );
  inv01 U7026 ( .Y(n13826), .A(n13828) );
  inv01 U7027 ( .Y(n13825), .A(n13834) );
  nand02 U7028 ( .Y(n13813), .A0(n13836), .A1(n13837) );
  inv01 U7029 ( .Y(n13837), .A(n13770) );
  nor02 U7030 ( .Y(n13836), .A0(n10301), .A1(n10367) );
  nand02 U7031 ( .Y(n13812), .A0(n10277), .A1(n13846) );
  nor02 U7032 ( .Y(n13846), .A0(n13850), .A1(n13851) );
  nand02 U7033 ( .Y(n13604), .A0(n13616), .A1(n13617) );
  inv01 U7034 ( .Y(v_count3287_5_), .A(n13618) );
  nand04 U7035 ( .Y(n13621), .A0(n13631), .A1(n13632), .A2(n12369), .A3(n10460) );
  inv01 U7036 ( .Y(v_count3287_4_), .A(n10646) );
  inv01 U7037 ( .Y(v_count3287_3_), .A(n13676) );
  nand04 U7038 ( .Y(n13679), .A0(n13684), .A1(n13685), .A2(n13686), .A3(n13687) );
  nand04 U7039 ( .Y(n13678), .A0(n13688), .A1(n13689), .A2(n13690), .A3(n13691) );
  inv01 U7040 ( .Y(v_count3287_2_), .A(n13695) );
  nand04 U7041 ( .Y(n13699), .A0(n13700), .A1(n13701), .A2(n13702), .A3(n13703) );
  nand04 U7042 ( .Y(n13696), .A0(n13710), .A1(n13711), .A2(n13712), .A3(n13713) );
  inv01 U7043 ( .Y(v_count3287_1_), .A(n13717) );
  nand04 U7044 ( .Y(n13721), .A0(n13722), .A1(n13723), .A2(n13724), .A3(n13725) );
  inv01 U7045 ( .Y(n13623), .A(n13726) );
  inv01 U7046 ( .Y(n13627), .A(n13728) );
  inv01 U7047 ( .Y(n13630), .A(n13729) );
  inv01 U7048 ( .Y(n13629), .A(n13730) );
  nand04 U7049 ( .Y(n13720), .A0(n13731), .A1(n13732), .A2(n13733), .A3(n13734) );
  and02 U7050 ( .Y(n13650), .A0(n12459), .A1(n13502) );
  inv01 U7051 ( .Y(n13638), .A(n13735) );
  inv01 U7052 ( .Y(n13640), .A(n13737) );
  inv01 U7053 ( .Y(n13637), .A(n13738) );
  nand04 U7054 ( .Y(n13719), .A0(n13739), .A1(n13740), .A2(n13741), .A3(n13742) );
  and02 U7055 ( .Y(n13662), .A0(s_fract_48_i[44]), .A1(n10339) );
  and03 U7056 ( .Y(n13643), .A0(n13428), .A1(n13749), .A2(n12418) );
  and03 U7057 ( .Y(n13645), .A0(n13751), .A1(n13752), .A2(s_fract_48_i[10]) );
  and03 U7058 ( .Y(n13648), .A0(n10423), .A1(n13753), .A2(s_fract_48_i[12]) );
  and03 U7059 ( .Y(n13646), .A0(n13752), .A1(n13754), .A2(n12922) );
  and02 U7060 ( .Y(n13649), .A0(s_fract_48_i[18]), .A1(n13757) );
  and02 U7061 ( .Y(n13647), .A0(n10570), .A1(n10477) );
  nand04 U7062 ( .Y(n13718), .A0(n13758), .A1(n13759), .A2(n13760), .A3(n10344) );
  and03 U7063 ( .Y(n13716), .A0(n13205), .A1(n13425), .A2(s_fract_48_i[6]) );
  and02 U7064 ( .Y(n13654), .A0(n10882), .A1(n10481) );
  and03 U7065 ( .Y(n13653), .A0(n13421), .A1(n13763), .A2(n12255) );
  and02 U7066 ( .Y(n13655), .A0(s_fract_48_i[34]), .A1(n13764) );
  and03 U7067 ( .Y(n13656), .A0(n10352), .A1(n13765), .A2(n12251) );
  and04 U7068 ( .Y(n13658), .A0(n12349), .A1(n13502), .A2(n13766), .A3(n13767)
         );
  and03 U7069 ( .Y(n13660), .A0(n13768), .A1(n13769), .A2(n13770) );
  and03 U7070 ( .Y(n13659), .A0(n13771), .A1(n13420), .A2(s_fract_48_i[38]) );
  and03 U7071 ( .Y(n13661), .A0(n10405), .A1(n13772), .A2(s_fract_48_i[40]) );
  nand04 U7072 ( .Y(v_count3287_0_), .A0(n13773), .A1(n13774), .A2(n13775), 
        .A3(n13776) );
  and02 U7073 ( .Y(n13628), .A0(n10721), .A1(n13428) );
  and02 U7074 ( .Y(n13626), .A0(n10416), .A1(n10423) );
  nand03 U7075 ( .Y(n13777), .A0(n13730), .A1(n13729), .A2(n13728) );
  nand03 U7076 ( .Y(n13728), .A0(n10477), .A1(n13779), .A2(s_fract_48_i[17])
         );
  nand03 U7077 ( .Y(n13729), .A0(n13502), .A1(n13766), .A2(n12409) );
  nand02 U7078 ( .Y(n13730), .A0(s_fract_48_i[15]), .A1(n13780) );
  and02 U7079 ( .Y(n13622), .A0(n10504), .A1(n13755) );
  and04 U7080 ( .Y(n13625), .A0(n12887), .A1(n13752), .A2(n13754), .A3(n13782)
         );
  and02 U7081 ( .Y(n13624), .A0(n10289), .A1(n13752) );
  nand03 U7082 ( .Y(n13781), .A0(n13727), .A1(n13668), .A2(n13737) );
  nand02 U7083 ( .Y(n13737), .A0(n10506), .A1(n13783) );
  nand04 U7084 ( .Y(n13726), .A0(n10724), .A1(n13427), .A2(n13749), .A3(n13784) );
  nand03 U7085 ( .Y(n13727), .A0(n10338), .A1(n13746), .A2(s_fract_48_i[45])
         );
  and02 U7086 ( .Y(n13743), .A0(n13783), .A1(n13785) );
  and03 U7087 ( .Y(n13783), .A0(n13745), .A1(n13786), .A2(n13744) );
  and04 U7088 ( .Y(n13636), .A0(n10830), .A1(n13420), .A2(n13763), .A3(n13790)
         );
  nand03 U7089 ( .Y(n13787), .A0(n13736), .A1(n13738), .A2(n13735) );
  nand02 U7090 ( .Y(n13735), .A0(n10574), .A1(n10352) );
  nand02 U7091 ( .Y(n13738), .A0(s_fract_48_i[41]), .A1(n13744) );
  nand02 U7092 ( .Y(n13736), .A0(s_fract_48_i[39]), .A1(n10405) );
  and03 U7093 ( .Y(n13634), .A0(n10481), .A1(n13794), .A2(s_fract_48_i[33]) );
  and02 U7094 ( .Y(n13633), .A0(n10822), .A1(n13421) );
  and02 U7095 ( .Y(n13762), .A0(n13764), .A1(n13795) );
  and03 U7096 ( .Y(n13764), .A0(n13794), .A1(n13796), .A2(n10481) );
  and03 U7097 ( .Y(n13788), .A0(n12919), .A1(n13798), .A2(n13502) );
  and03 U7098 ( .Y(n13778), .A0(n13428), .A1(n13800), .A2(n13750) );
  and02 U7099 ( .Y(n13748), .A0(n13757), .A1(n13801) );
  and03 U7100 ( .Y(n13757), .A0(n13779), .A1(n13802), .A2(n10477) );
  and03 U7101 ( .Y(n13780), .A0(n13756), .A1(n13804), .A2(n13755) );
  aoi21 U7102 ( .Y(n13809), .A0(n10378), .A1(n13811), .B0(s_fract_48_i[3]) );
  inv01 U7103 ( .Y(n13808), .A(n13425) );
  nand04 U7104 ( .Y(n13873), .A0(n10386), .A1(n13874), .A2(n13875), .A3(n13876) );
  nand04 U7105 ( .Y(n13871), .A0(n13880), .A1(n10427), .A2(n13881), .A3(n13882) );
  nand04 U7106 ( .Y(n13889), .A0(n12437), .A1(n13890), .A2(n13891), .A3(n13892) );
  nand04 U7107 ( .Y(n13888), .A0(n13893), .A1(n13894), .A2(n13895), .A3(n13896) );
  inv01 U7108 ( .Y(n13817), .A(n10299) );
  nand04 U7109 ( .Y(n13906), .A0(n13915), .A1(n13913), .A2(n13914), .A3(n13912) );
  inv01 U7110 ( .Y(n13829), .A(n10374) );
  inv01 U7111 ( .Y(n13832), .A(n13920) );
  inv01 U7112 ( .Y(n13835), .A(n13921) );
  nand04 U7113 ( .Y(n13905), .A0(n13925), .A1(n13923), .A2(n13924), .A3(n13922) );
  and02 U7114 ( .Y(n13839), .A0(n10833), .A1(n12351) );
  and04 U7115 ( .Y(n13856), .A0(n13926), .A1(n12460), .A2(n13767), .A3(n13927)
         );
  and02 U7116 ( .Y(n13840), .A0(n10306), .A1(n10884) );
  and03 U7117 ( .Y(n13841), .A0(n12250), .A1(n13928), .A2(n13510) );
  and02 U7118 ( .Y(n13838), .A0(n13929), .A1(s_fract_48_i[30]) );
  and03 U7119 ( .Y(n13843), .A0(n12256), .A1(n13930), .A2(n13433) );
  and02 U7120 ( .Y(n13842), .A0(s_fract_48_i[38]), .A1(n12445) );
  and03 U7121 ( .Y(n13844), .A0(n13433), .A1(s_fract_48_i[34]), .A2(n13771) );
  and04 U7122 ( .Y(n13845), .A0(s_fract_48_i[2]), .A1(n13916), .A2(n12842), 
        .A3(n13931) );
  nand02 U7123 ( .Y(n13935), .A0(n13534), .A1(n13785) );
  and03 U7124 ( .Y(n13848), .A0(n13431), .A1(n13937), .A2(n12419) );
  inv01 U7125 ( .Y(n13901), .A(n13938) );
  and02 U7126 ( .Y(n13847), .A0(n10568), .A1(n10479) );
  and03 U7127 ( .Y(n13849), .A0(n13431), .A1(n13750), .A2(s_fract_48_i[18]) );
  and02 U7128 ( .Y(n13850), .A0(s_fract_48_i[14]), .A1(n13939) );
  and03 U7129 ( .Y(n13853), .A0(n10421), .A1(n13753), .A2(s_fract_48_i[10]) );
  and03 U7130 ( .Y(n13851), .A0(n10475), .A1(n13756), .A2(s_fract_48_i[12]) );
  and03 U7131 ( .Y(n13854), .A0(n13941), .A1(n13942), .A2(n12924) );
  and02 U7132 ( .Y(n13855), .A0(s_fract_48_i[22]), .A1(n13943) );
  and03 U7133 ( .Y(n13852), .A0(n13941), .A1(n13751), .A2(s_fract_48_i[6]) );
  and02 U7134 ( .Y(s_zeros1047_0_), .A0(n13944), .A1(n13769) );
  nand04 U7135 ( .Y(n13944), .A0(n13945), .A1(n13946), .A2(n13947), .A3(n13948) );
  and03 U7136 ( .Y(n13823), .A0(n13916), .A1(n13205), .A2(s_fract_48_i[1]) );
  inv01 U7137 ( .Y(n13761), .A(n13714) );
  nor02 U7138 ( .Y(n13714), .A0(s_fract_48_i[3]), .A1(s_fract_48_i[2]) );
  inv01 U7139 ( .Y(n13715), .A(n12842) );
  and03 U7140 ( .Y(n13824), .A0(n13916), .A1(n12842), .A2(s_fract_48_i[3]) );
  and04 U7141 ( .Y(n13820), .A0(n10820), .A1(n13433), .A2(n13790), .A3(n13930)
         );
  or03 U7142 ( .Y(n13949), .A0(n13821), .A1(n13822), .A2(n13819) );
  and02 U7143 ( .Y(n13819), .A0(n10293), .A1(n13510) );
  and02 U7144 ( .Y(n13822), .A0(n10831), .A1(n13433) );
  and02 U7145 ( .Y(n13818), .A0(s_fract_48_i[33]), .A1(n13951) );
  and02 U7146 ( .Y(n13926), .A0(n13510), .A1(n13952) );
  nand02 U7147 ( .Y(n13950), .A0(n13921), .A1(n10299) );
  nand04 U7148 ( .Y(n13911), .A0(n10573), .A1(n13510), .A2(n13789), .A3(n13928) );
  nand03 U7149 ( .Y(n13921), .A0(n13510), .A1(n12919), .A2(s_fract_48_i[23])
         );
  and02 U7150 ( .Y(n13834), .A0(n10377), .A1(n13916) );
  and02 U7151 ( .Y(n13833), .A0(n12888), .A1(n13941) );
  nand03 U7152 ( .Y(n13953), .A0(n13895), .A1(n13920), .A2(n10374) );
  nand04 U7153 ( .Y(n13918), .A0(n10720), .A1(n13430), .A2(n13784), .A3(n13937) );
  nand02 U7154 ( .Y(n13920), .A0(n10503), .A1(n10474) );
  nand03 U7155 ( .Y(n13919), .A0(n10479), .A1(n13779), .A2(s_fract_48_i[15])
         );
  and02 U7156 ( .Y(n13828), .A0(n10418), .A1(n10421) );
  and02 U7157 ( .Y(n13940), .A0(n13939), .A1(n13804) );
  and03 U7158 ( .Y(n13939), .A0(n13803), .A1(n13779), .A2(n10479) );
  and02 U7159 ( .Y(n13827), .A0(n10725), .A1(n13431) );
  and03 U7160 ( .Y(n13955), .A0(n13750), .A1(n13801), .A2(n13430) );
  and02 U7161 ( .Y(n13936), .A0(n13943), .A1(n13800) );
  and03 U7162 ( .Y(n13943), .A0(n12919), .A1(n13799), .A2(n13510) );
  and03 U7163 ( .Y(n13929), .A0(n13797), .A1(n13794), .A2(n10306) );
  and03 U7164 ( .Y(n13951), .A0(n13433), .A1(n13795), .A2(n13771) );
  nand02 U7165 ( .Y(n13902), .A0(n13745), .A1(n13791) );
  ao21 U7166 ( .Y(s_shr25775_5_), .A0(n9756), .A1(n13537), .B0(n13957) );
  ao21 U7167 ( .Y(s_shr25775_4_), .A0(n9636), .A1(n13537), .B0(n13957) );
  ao21 U7168 ( .Y(s_shr25775_3_), .A0(n9758), .A1(n13537), .B0(n13957) );
  ao21 U7169 ( .Y(s_shr25775_2_), .A0(n9634), .A1(n13537), .B0(n13957) );
  ao21 U7170 ( .Y(s_shr25775_1_), .A0(n9760), .A1(n13537), .B0(n13957) );
  nand02 U7171 ( .Y(s_shr25775_0_), .A0(n9800), .A1(n13961) );
  nand02 U7172 ( .Y(n13961), .A0(n9877), .A1(n13537) );
  nand02 U7173 ( .Y(n13963), .A0(n10401), .A1(n____return5956_5_) );
  nor02 U7174 ( .Y(n13958), .A0(n13959), .A1(n13609) );
  inv01 U7175 ( .Y(n13609), .A(n____return5956_3_) );
  nand02 U7176 ( .Y(n13959), .A0(n12416), .A1(n____return5956_2_) );
  nor02 U7177 ( .Y(n13960), .A0(n13962), .A1(n13613) );
  inv01 U7178 ( .Y(n13613), .A(n____return5956_1_) );
  nand02 U7179 ( .Y(n13962), .A0(n____return5956_0_), .A1(n13511) );
  nor02 U7180 ( .Y(n13965), .A0(n13616), .A1(n13615) );
  ao21 U7181 ( .Y(n13964), .A0(n13537), .A1(n13615), .B0(n13966) );
  ao22 U7182 ( .Y(s_output_o_9_), .A0(n13570), .A1(n14418), .B0(n13571), .B1(
        n14400) );
  ao22 U7183 ( .Y(s_output_o_8_), .A0(n14400), .A1(n13570), .B0(n13571), .B1(
        n14401) );
  ao22 U7184 ( .Y(s_output_o_7_), .A0(n13570), .A1(n14401), .B0(n13571), .B1(
        n14402) );
  ao22 U7185 ( .Y(s_output_o_6_), .A0(n13570), .A1(n14402), .B0(n13571), .B1(
        n14403) );
  ao22 U7186 ( .Y(s_output_o_5_), .A0(n13570), .A1(n14403), .B0(n13571), .B1(
        n14404) );
  ao22 U7187 ( .Y(s_output_o_4_), .A0(n13570), .A1(n14404), .B0(n13571), .B1(
        n14405) );
  ao22 U7188 ( .Y(s_output_o_3_), .A0(n13570), .A1(n14405), .B0(n13571), .B1(
        n14406) );
  ao22 U7189 ( .Y(s_output_o_2_), .A0(n13570), .A1(n14406), .B0(n13571), .B1(
        n14408) );
  ao221 U7190 ( .Y(s_output_o_26_), .A0(s_expo2b[3]), .A1(n13471), .B0(
        n____return7168_3_), .B1(n13474), .C0(n12915) );
  ao221 U7191 ( .Y(s_output_o_25_), .A0(s_expo2b[2]), .A1(n13471), .B0(
        n____return7168_2_), .B1(n13474), .C0(n12915) );
  ao22 U7192 ( .Y(s_output_o_21_), .A0(n13570), .A1(s_frac_rnd_22_), .B0(
        n13571), .B1(n14407) );
  ao22 U7193 ( .Y(s_output_o_20_), .A0(n13570), .A1(n14407), .B0(n13571), .B1(
        n14409) );
  ao22 U7194 ( .Y(s_output_o_1_), .A0(n13570), .A1(n14408), .B0(n13571), .B1(
        s_frac_rnd_1_) );
  ao22 U7195 ( .Y(s_output_o_19_), .A0(n13570), .A1(n14409), .B0(n13571), .B1(
        n14410) );
  ao22 U7196 ( .Y(s_output_o_18_), .A0(n13570), .A1(n14410), .B0(n13571), .B1(
        n14411) );
  ao22 U7197 ( .Y(s_output_o_17_), .A0(n13570), .A1(n14411), .B0(n13571), .B1(
        n14412) );
  ao22 U7198 ( .Y(s_output_o_16_), .A0(n13570), .A1(n14412), .B0(n13571), .B1(
        n14413) );
  ao22 U7199 ( .Y(s_output_o_15_), .A0(n13570), .A1(n14413), .B0(n13571), .B1(
        n14414) );
  ao22 U7200 ( .Y(s_output_o_14_), .A0(n13570), .A1(n14414), .B0(n13571), .B1(
        n14415) );
  ao22 U7201 ( .Y(s_output_o_13_), .A0(n13570), .A1(n14415), .B0(n13571), .B1(
        n14416) );
  ao22 U7202 ( .Y(s_output_o_12_), .A0(n13570), .A1(n14416), .B0(n13571), .B1(
        n14417) );
  ao22 U7203 ( .Y(s_output_o_11_), .A0(n13570), .A1(n14417), .B0(n13571), .B1(
        n14419) );
  ao22 U7204 ( .Y(s_output_o_10_), .A0(n13570), .A1(n14419), .B0(n13571), .B1(
        n14418) );
  nor02 U7205 ( .Y(n13968), .A0(n13993), .A1(n13994) );
  inv01 U7206 ( .Y(n13992), .A(s_frac_rnd_1_) );
  nor02 U7207 ( .Y(n13967), .A0(n13993), .A1(n13995) );
  ao21 U7208 ( .Y(n13993), .A0(n10285), .A1(n10303), .B0(n12915) );
  nand02 U7209 ( .Y(n13980), .A0(n13996), .A1(n13997) );
  inv01 U7210 ( .Y(n13988), .A(n13999) );
  nand04 U7211 ( .Y(n13990), .A0(n12274), .A1(n12353), .A2(n12359), .A3(n12403) );
  nand03 U7212 ( .Y(n14002), .A0(n14437), .A1(n14438), .A2(n14436) );
  nand03 U7213 ( .Y(n14003), .A0(n14440), .A1(n14441), .A2(n14439) );
  nand03 U7214 ( .Y(n14004), .A0(n14443), .A1(n14444), .A2(n14442) );
  nand02 U7215 ( .Y(n14005), .A0(n14445), .A1(n14446) );
  nand04 U7216 ( .Y(n13991), .A0(n12278), .A1(n12357), .A2(n12361), .A3(n12407) );
  nand03 U7217 ( .Y(n14006), .A0(n14424), .A1(n14425), .A2(n14423) );
  nand03 U7218 ( .Y(n14007), .A0(n14427), .A1(n14428), .A2(n14426) );
  nand03 U7219 ( .Y(n14008), .A0(n14430), .A1(n14431), .A2(n14429) );
  nand02 U7220 ( .Y(n14009), .A0(n14432), .A1(n14433) );
  nand02 U7221 ( .Y(n13997), .A0(n9931), .A1(n13996) );
  inv01 U7222 ( .Y(n13996), .A(n13989) );
  nand02 U7223 ( .Y(n13989), .A0(n13986), .A1(n13985) );
  nand02 U7224 ( .Y(n13985), .A0(n10692), .A1(n10863) );
  nand02 U7225 ( .Y(n13986), .A0(n10690), .A1(n10861) );
  inv01 U7226 ( .Y(n13994), .A(n13995) );
  nand02 U7227 ( .Y(n13995), .A0(s_shr3), .A1(n10304) );
  nand04 U7228 ( .Y(n14011), .A0(s_expo2b[3]), .A1(s_expo2b[1]), .A2(n10409), 
        .A3(n12413) );
  nand04 U7229 ( .Y(n14010), .A0(n____return7168_3_), .A1(n____return7168_2_), 
        .A2(n10425), .A3(n14013) );
  inv01 U7230 ( .Y(n13971), .A(n____return7168_7_) );
  inv01 U7231 ( .Y(n13975), .A(n____return7168_6_) );
  inv01 U7232 ( .Y(n13977), .A(n____return7168_5_) );
  inv01 U7233 ( .Y(n13984), .A(n____return7168_0_) );
  inv01 U7234 ( .Y(n13982), .A(n____return7168_1_) );
  mux21 U7235 ( .Y(s_frac_rnd7043_9_), .A0(n14014), .A1(n14465), .S0(n13578)
         );
  inv01 U7236 ( .Y(n14014), .A(n____return7070_9_) );
  mux21 U7237 ( .Y(s_frac_rnd7043_8_), .A0(n14016), .A1(n14466), .S0(n13578)
         );
  inv01 U7238 ( .Y(n14016), .A(n____return7070_8_) );
  mux21 U7239 ( .Y(s_frac_rnd7043_7_), .A0(n14017), .A1(n14467), .S0(n13578)
         );
  inv01 U7240 ( .Y(n14017), .A(n____return7070_7_) );
  mux21 U7241 ( .Y(s_frac_rnd7043_6_), .A0(n14018), .A1(n14468), .S0(n13578)
         );
  inv01 U7242 ( .Y(n14018), .A(n____return7070_6_) );
  mux21 U7243 ( .Y(s_frac_rnd7043_5_), .A0(n14019), .A1(n14469), .S0(n13578)
         );
  inv01 U7244 ( .Y(n14019), .A(n____return7070_5_) );
  mux21 U7245 ( .Y(s_frac_rnd7043_4_), .A0(n14020), .A1(n14470), .S0(n13578)
         );
  inv01 U7246 ( .Y(n14020), .A(n____return7070_4_) );
  mux21 U7247 ( .Y(s_frac_rnd7043_3_), .A0(n14021), .A1(n14471), .S0(n13578)
         );
  inv01 U7248 ( .Y(n14021), .A(n____return7070_3_) );
  mux21 U7249 ( .Y(s_frac_rnd7043_2_), .A0(n14022), .A1(n14472), .S0(n13578)
         );
  inv01 U7250 ( .Y(n14022), .A(n____return7070_2_) );
  mux21 U7251 ( .Y(s_frac_rnd7043_24_), .A0(n14023), .A1(n14473), .S0(n13578)
         );
  inv01 U7252 ( .Y(n14023), .A(n____return7070_24_) );
  inv01 U7253 ( .Y(s_frac_rnd7043_23_), .A(n14024) );
  mux21 U7254 ( .Y(n14024), .A0(n7072_23_), .A1(n13520), .S0(n13578) );
  mux21 U7255 ( .Y(s_frac_rnd7043_22_), .A0(n14025), .A1(n14474), .S0(n13578)
         );
  inv01 U7256 ( .Y(n14025), .A(n____return7070_22_) );
  mux21 U7257 ( .Y(s_frac_rnd7043_21_), .A0(n14026), .A1(n14475), .S0(n13578)
         );
  inv01 U7258 ( .Y(n14026), .A(n____return7070_21_) );
  mux21 U7259 ( .Y(s_frac_rnd7043_20_), .A0(n14027), .A1(n14476), .S0(n13578)
         );
  inv01 U7260 ( .Y(n14027), .A(n____return7070_20_) );
  mux21 U7261 ( .Y(s_frac_rnd7043_1_), .A0(n14028), .A1(n14477), .S0(n13578)
         );
  inv01 U7262 ( .Y(n14028), .A(n____return7070_1_) );
  mux21 U7263 ( .Y(s_frac_rnd7043_19_), .A0(n14029), .A1(n14478), .S0(n13578)
         );
  inv01 U7264 ( .Y(n14029), .A(n____return7070_19_) );
  mux21 U7265 ( .Y(s_frac_rnd7043_18_), .A0(n14030), .A1(n14479), .S0(n13578)
         );
  inv01 U7266 ( .Y(n14030), .A(n____return7070_18_) );
  mux21 U7267 ( .Y(s_frac_rnd7043_17_), .A0(n14031), .A1(n14480), .S0(n13578)
         );
  inv01 U7268 ( .Y(n14031), .A(n____return7070_17_) );
  mux21 U7269 ( .Y(s_frac_rnd7043_16_), .A0(n14032), .A1(n14481), .S0(n13578)
         );
  inv01 U7270 ( .Y(n14032), .A(n____return7070_16_) );
  mux21 U7271 ( .Y(s_frac_rnd7043_15_), .A0(n14033), .A1(n14482), .S0(n13578)
         );
  inv01 U7272 ( .Y(n14033), .A(n____return7070_15_) );
  mux21 U7273 ( .Y(s_frac_rnd7043_14_), .A0(n14034), .A1(n14483), .S0(n13578)
         );
  inv01 U7274 ( .Y(n14034), .A(n____return7070_14_) );
  mux21 U7275 ( .Y(s_frac_rnd7043_13_), .A0(n14035), .A1(n14484), .S0(n13578)
         );
  inv01 U7276 ( .Y(n14035), .A(n____return7070_13_) );
  mux21 U7277 ( .Y(s_frac_rnd7043_12_), .A0(n14036), .A1(n14485), .S0(n13578)
         );
  inv01 U7278 ( .Y(n14036), .A(n____return7070_12_) );
  mux21 U7279 ( .Y(s_frac_rnd7043_11_), .A0(n14037), .A1(n14486), .S0(n13578)
         );
  inv01 U7280 ( .Y(n14037), .A(n____return7070_11_) );
  mux21 U7281 ( .Y(s_frac_rnd7043_10_), .A0(n14038), .A1(n14487), .S0(n13578)
         );
  inv01 U7282 ( .Y(n14038), .A(n____return7070_10_) );
  inv01 U7283 ( .Y(s_frac_rnd7043_0_), .A(n14039) );
  mux21 U7284 ( .Y(n14039), .A0(n____return7070_0_), .A1(s_frac2a_23_), .S0(
        n13578) );
  mux21 U7285 ( .Y(n14015), .A0(n14040), .A1(n14041), .S0(s_rmode_i_1_) );
  nor02 U7286 ( .Y(n14041), .A0(n13998), .A1(n9782) );
  nand04 U7287 ( .Y(n14042), .A0(n12276), .A1(n12355), .A2(n12363), .A3(n12405) );
  nand03 U7288 ( .Y(n14044), .A0(n14491), .A1(n14492), .A2(n14490) );
  nand02 U7289 ( .Y(n14045), .A0(n14493), .A1(n14494) );
  nand03 U7290 ( .Y(n14046), .A0(n14496), .A1(n14497), .A2(n14495) );
  nand02 U7291 ( .Y(n14047), .A0(n14498), .A1(n14499) );
  inv01 U7292 ( .Y(n14043), .A(n14489) );
  nand03 U7293 ( .Y(s_frac2a6207_9_), .A0(n10127), .A1(n10231), .A2(n14048) );
  nand03 U7294 ( .Y(s_frac2a6207_8_), .A0(n10137), .A1(n10168), .A2(n14062) );
  inv01 U7295 ( .Y(n14066), .A(n14068) );
  nand03 U7296 ( .Y(s_frac2a6207_7_), .A0(n10135), .A1(n10237), .A2(n14071) );
  nand03 U7297 ( .Y(s_frac2a6207_6_), .A0(n10117), .A1(n10247), .A2(n14079) );
  nand03 U7298 ( .Y(s_frac2a6207_5_), .A0(n10109), .A1(n10235), .A2(n14087) );
  nand03 U7299 ( .Y(s_frac2a6207_4_), .A0(n10107), .A1(n10233), .A2(n14092) );
  nand02 U7300 ( .Y(s_frac2a6207_47_), .A0(n14096), .A1(n14097) );
  nand03 U7301 ( .Y(s_frac2a6207_46_), .A0(n10202), .A1(n10170), .A2(n14115)
         );
  nand03 U7302 ( .Y(s_frac2a6207_45_), .A0(n10113), .A1(n10172), .A2(n14123)
         );
  nand03 U7303 ( .Y(s_frac2a6207_44_), .A0(n10115), .A1(n10174), .A2(n14131)
         );
  nand03 U7304 ( .Y(s_frac2a6207_43_), .A0(n10160), .A1(n10251), .A2(n14139)
         );
  nand03 U7305 ( .Y(s_frac2a6207_42_), .A0(n10143), .A1(n10239), .A2(n14145)
         );
  nand03 U7306 ( .Y(s_frac2a6207_41_), .A0(n10157), .A1(n10245), .A2(n14151)
         );
  nand03 U7307 ( .Y(s_frac2a6207_40_), .A0(n10155), .A1(n10243), .A2(n14154)
         );
  nand03 U7308 ( .Y(s_frac2a6207_3_), .A0(n10119), .A1(n10184), .A2(n14157) );
  nand03 U7309 ( .Y(s_frac2a6207_39_), .A0(n10151), .A1(n10197), .A2(n14167)
         );
  nand03 U7310 ( .Y(s_frac2a6207_38_), .A0(n10153), .A1(n14170), .A2(n14171)
         );
  nand03 U7311 ( .Y(s_frac2a6207_37_), .A0(n10145), .A1(n10178), .A2(n14174)
         );
  nand03 U7312 ( .Y(s_frac2a6207_36_), .A0(n10149), .A1(n10180), .A2(n14177)
         );
  nand03 U7313 ( .Y(s_frac2a6207_35_), .A0(n10131), .A1(n10253), .A2(n14181)
         );
  nand03 U7314 ( .Y(s_frac2a6207_34_), .A0(n10133), .A1(n10249), .A2(n14184)
         );
  nand03 U7315 ( .Y(s_frac2a6207_33_), .A0(n10129), .A1(n10257), .A2(n14190)
         );
  nand03 U7316 ( .Y(s_frac2a6207_32_), .A0(n10121), .A1(n10166), .A2(n14195)
         );
  nor02 U7317 ( .Y(n14098), .A0(n13527), .A1(n14199) );
  and03 U7318 ( .Y(n14113), .A0(n12447), .A1(n14202), .A2(s_shl2_5_) );
  nor02 U7319 ( .Y(n14102), .A0(n13527), .A1(n13567) );
  nor02 U7320 ( .Y(n14111), .A0(n14204), .A1(n13527) );
  ao221 U7321 ( .Y(s_frac2a6207_31_), .A0(n14114), .A1(n13573), .B0(n14205), 
        .B1(n13569), .C0(n14206) );
  ao22 U7322 ( .Y(n14206), .A0(n12921), .A1(n13010), .B0(n13565), .B1(n14110)
         );
  inv01 U7323 ( .Y(n14207), .A(n14144) );
  ao221 U7324 ( .Y(s_frac2a6207_30_), .A0(n14117), .A1(n13573), .B0(n14212), 
        .B1(n13569), .C0(n14213) );
  ao22 U7325 ( .Y(n14213), .A0(n12921), .A1(n14116), .B0(n13565), .B1(n14118)
         );
  inv01 U7326 ( .Y(n14214), .A(n14150) );
  nand03 U7327 ( .Y(s_frac2a6207_2_), .A0(n10164), .A1(n10176), .A2(n14217) );
  inv01 U7328 ( .Y(n14223), .A(n14153) );
  inv01 U7329 ( .Y(n14227), .A(n14156) );
  inv01 U7330 ( .Y(n14226), .A(n14231) );
  inv01 U7331 ( .Y(n14141), .A(n14233) );
  ao221 U7332 ( .Y(s_frac2a6207_25_), .A0(n14152), .A1(n13565), .B0(n14055), 
        .B1(n13569), .C0(n14238) );
  ao22 U7333 ( .Y(n14238), .A0(n13564), .A1(n12797), .B0(n13573), .B1(n14059)
         );
  inv01 U7334 ( .Y(n14239), .A(n14240) );
  oai22 U7335 ( .Y(n14057), .A0(n14241), .A1(n13558), .B0(n13418), .B1(n13577)
         );
  inv01 U7336 ( .Y(n14242), .A(n14248) );
  inv01 U7337 ( .Y(n14253), .A(n14256) );
  oai22 U7338 ( .Y(n14067), .A0(n14257), .A1(n13558), .B0(n14258), .B1(n13577)
         );
  ao22 U7339 ( .Y(n14262), .A0(n13561), .A1(n14264), .B0(n13556), .B1(n14265)
         );
  inv01 U7340 ( .Y(n14252), .A(n14155) );
  ao221 U7341 ( .Y(s_frac2a6207_23_), .A0(n14168), .A1(n13565), .B0(n14076), 
        .B1(n13569), .C0(n14268) );
  ao22 U7342 ( .Y(n14268), .A0(n13564), .A1(n14077), .B0(n13573), .B1(n10858)
         );
  ao22 U7343 ( .Y(n14078), .A0(n14269), .A1(n13574), .B0(n14158), .B1(n13566)
         );
  inv01 U7344 ( .Y(n14274), .A(n14278) );
  ao221 U7345 ( .Y(s_frac2a6207_22_), .A0(n14172), .A1(n13565), .B0(n14084), 
        .B1(n13569), .C0(n14281) );
  ao22 U7346 ( .Y(n14281), .A0(n13564), .A1(n14085), .B0(n13573), .B1(n10859)
         );
  ao22 U7347 ( .Y(n14086), .A0(n14282), .A1(n13574), .B0(n14187), .B1(n13566)
         );
  ao221 U7348 ( .Y(s_frac2a6207_21_), .A0(n14175), .A1(n13565), .B0(n14088), 
        .B1(n13569), .C0(n14292) );
  ao22 U7349 ( .Y(n14292), .A0(n13564), .A1(n14089), .B0(n13573), .B1(n12753)
         );
  oai22 U7350 ( .Y(n14090), .A0(n13394), .A1(n13567), .B0(n13423), .B1(n13575)
         );
  ao221 U7351 ( .Y(s_frac2a6207_20_), .A0(n14178), .A1(n13565), .B0(n14094), 
        .B1(n13569), .C0(n14298) );
  ao22 U7352 ( .Y(n14298), .A0(n13564), .A1(n14095), .B0(n13573), .B1(n10275)
         );
  nand03 U7353 ( .Y(s_frac2a6207_1_), .A0(n10139), .A1(n10190), .A2(n14306) );
  inv01 U7354 ( .Y(n14315), .A(n14072) );
  inv01 U7355 ( .Y(n14312), .A(n14165) );
  inv01 U7356 ( .Y(n14323), .A(n14081) );
  inv01 U7357 ( .Y(n14320), .A(n14186) );
  inv01 U7358 ( .Y(n14328), .A(n14054) );
  inv01 U7359 ( .Y(n14327), .A(n14192) );
  inv01 U7360 ( .Y(n14329), .A(n14197) );
  nand02 U7361 ( .Y(n14311), .A0(n13573), .A1(n13574) );
  nand02 U7362 ( .Y(n14221), .A0(s_shl2_4_), .A1(n14332) );
  nand03 U7363 ( .Y(s_frac2a6207_15_), .A0(n10125), .A1(n10192), .A2(n14333)
         );
  nand03 U7364 ( .Y(s_frac2a6207_14_), .A0(n10123), .A1(n10255), .A2(n14334)
         );
  nand03 U7365 ( .Y(s_frac2a6207_13_), .A0(n10186), .A1(n10241), .A2(n14335)
         );
  inv01 U7366 ( .Y(n14336), .A(n12891) );
  inv01 U7367 ( .Y(n14125), .A(n12835) );
  nand03 U7368 ( .Y(s_frac2a6207_12_), .A0(n10194), .A1(n10206), .A2(n14344)
         );
  inv01 U7369 ( .Y(n14133), .A(n12833) );
  nor02 U7370 ( .Y(n14210), .A0(n14299), .A1(n14300) );
  nand03 U7371 ( .Y(s_frac2a6207_11_), .A0(n10141), .A1(n14349), .A2(n11053)
         );
  nand02 U7372 ( .Y(n14232), .A0(n9879), .A1(n14352) );
  inv01 U7373 ( .Y(n14273), .A(n14318) );
  inv01 U7374 ( .Y(n14271), .A(n13010) );
  inv01 U7375 ( .Y(n14349), .A(n14354) );
  nand03 U7376 ( .Y(s_frac2a6207_10_), .A0(n10111), .A1(n10188), .A2(n14357)
         );
  nor02 U7377 ( .Y(n14060), .A0(n13568), .A1(n13577) );
  inv01 U7378 ( .Y(n14146), .A(n12262) );
  nor02 U7379 ( .Y(n14270), .A0(n14300), .A1(s_shl2_3_) );
  nor02 U7380 ( .Y(n14209), .A0(n14299), .A1(s_shl2_2_) );
  inv01 U7381 ( .Y(n14299), .A(s_shl2_3_) );
  and02 U7382 ( .Y(n14108), .A0(s_shl2_1_), .A1(s_shl2_0_) );
  nand02 U7383 ( .Y(n14106), .A0(s_shl2_1_), .A1(n14360) );
  or02 U7384 ( .Y(n14105), .A0(n14360), .A1(s_shl2_1_) );
  inv01 U7385 ( .Y(n14360), .A(s_shl2_0_) );
  inv01 U7386 ( .Y(n14058), .A(n14198) );
  inv01 U7387 ( .Y(n14361), .A(n12914) );
  inv01 U7388 ( .Y(n14321), .A(n14288) );
  nand03 U7389 ( .Y(s_frac2a6207_0_), .A0(n10147), .A1(n10182), .A2(n14364) );
  nor02 U7390 ( .Y(n14200), .A0(n13768), .A1(n14342) );
  nor02 U7391 ( .Y(n14109), .A0(s_shl2_1_), .A1(s_shl2_0_) );
  nor02 U7392 ( .Y(n14100), .A0(n13527), .A1(n13575) );
  nor02 U7393 ( .Y(n14201), .A0(s_shl2_3_), .A1(s_shl2_2_) );
  nand02 U7394 ( .Y(n14198), .A0(n9627), .A1(n14202) );
  inv01 U7395 ( .Y(n14202), .A(s_shl2_4_) );
  nor02 U7396 ( .Y(n14332), .A0(n14365), .A1(s_shl2_5_) );
  inv01 U7397 ( .Y(n14365), .A(n12447) );
  inv01 U7398 ( .Y(n14366), .A(n14367) );
  nor02 U7399 ( .Y(n14051), .A0(n13568), .A1(n13558) );
  inv01 U7400 ( .Y(n14370), .A(n14070) );
  nand02 U7401 ( .Y(n14230), .A0(s_shr2_4_), .A1(n14371) );
  nor02 U7402 ( .Y(n14049), .A0(n13568), .A1(n14338) );
  nor02 U7403 ( .Y(n14053), .A0(n13568), .A1(n13562) );
  nand02 U7404 ( .Y(n14222), .A0(n14371), .A1(n14372) );
  nor02 U7405 ( .Y(n14367), .A0(n13577), .A1(s_shr2_4_) );
  nor02 U7406 ( .Y(n14260), .A0(s_shr2_3_), .A1(s_shr2_2_) );
  nor02 U7407 ( .Y(n14162), .A0(s_shr2_1_), .A1(s_shr2_0_) );
  mux21 U7408 ( .Y(n14373), .A0(n6653_8_), .A1(s_expo1[8]), .S0(s_frac2a_46_)
         );
  inv01 U7409 ( .Y(s_expo2b[7]), .A(n13969) );
  inv01 U7410 ( .Y(s_expo2b[6]), .A(n13974) );
  inv01 U7411 ( .Y(s_expo2b[5]), .A(n13976) );
  inv01 U7412 ( .Y(s_expo2b[4]), .A(n13978) );
  mux21 U7413 ( .Y(n14374), .A0(n____return6651_3_), .A1(s_expo1[3]), .S0(
        n13520) );
  mux21 U7414 ( .Y(n14012), .A0(n____return6651_2_), .A1(s_expo1[2]), .S0(
        s_frac2a_46_) );
  mux21 U7415 ( .Y(n13983), .A0(n____return6651_0_), .A1(s_expo1[0]), .S0(
        n13520) );
  ao21 U7416 ( .Y(s_expo15773_7_), .A0(s_exp_10b[7]), .A1(n13966), .B0(n14375)
         );
  ao21 U7417 ( .Y(s_expo15773_6_), .A0(s_exp_10b[6]), .A1(n13966), .B0(n14375)
         );
  ao21 U7418 ( .Y(s_expo15773_5_), .A0(s_exp_10b[5]), .A1(n13966), .B0(n14375)
         );
  ao21 U7419 ( .Y(s_expo15773_4_), .A0(s_exp_10b[4]), .A1(n13966), .B0(n14375)
         );
  ao21 U7420 ( .Y(s_expo15773_3_), .A0(s_exp_10b[3]), .A1(n13966), .B0(n14375)
         );
  ao21 U7421 ( .Y(s_expo15773_2_), .A0(s_exp_10b[2]), .A1(n13966), .B0(n14375)
         );
  ao21 U7422 ( .Y(s_expo15773_1_), .A0(s_exp_10b[1]), .A1(n13966), .B0(n14375)
         );
  inv01 U7423 ( .Y(n14376), .A(s_exp_10b[8]) );
  or02 U7424 ( .Y(s_expo15773_0_), .A0(n13602), .A1(s_exp_10b[0]) );
  or02 U7425 ( .Y(n14379), .A0(s_exp_10b[7]), .A1(s_exp_10b[4]) );
  nor02 U7426 ( .Y(U1086_U4_Z_6), .A0(n13616), .A1(n10507) );
  inv01 U7427 ( .Y(n13603), .A(s_zeros[5]) );
  inv01 U7428 ( .Y(n13606), .A(s_zeros[4]) );
  inv01 U7429 ( .Y(n13608), .A(s_zeros[3]) );
  inv01 U7430 ( .Y(n13610), .A(s_zeros[2]) );
  inv01 U7431 ( .Y(n13612), .A(s_zeros[1]) );
  nand02 U7432 ( .Y(U1086_U3_Z_0), .A0(n13616), .A1(n13614) );
  inv01 U7433 ( .Y(n13614), .A(s_zeros[0]) );
  ao21 U7434 ( .Y(n13956), .A0(n10835), .A1(n14381), .B0(s_exp_10a_9_) );
  xor2 U7435 ( .Y(s_exp_10a_9_), .A0(n14382), .A1(n14500) );
  nand02 U7436 ( .Y(n14382), .A0(n10473), .A1(s_exp_10_i_8_) );
  xor2 U7437 ( .Y(s_exp_10a_7_), .A0(s_exp_10_i_7_), .A1(n14385) );
  and02 U7438 ( .Y(n14385), .A0(s_exp_10_i_6_), .A1(n12844) );
  xor2 U7439 ( .Y(s_exp_10a_8_), .A0(s_exp_10_i_8_), .A1(n10473) );
  and03 U7440 ( .Y(n14383), .A0(n12844), .A1(s_exp_10_i_6_), .A2(s_exp_10_i_7_) );
  xnor2 U7441 ( .Y(n14380), .A0(n12843), .A1(s_exp_10_i_6_) );
  and03 U7442 ( .Y(n14386), .A0(s_exp_10_i_4_), .A1(n14387), .A2(s_exp_10_i_5_) );
  or02 U7443 ( .Y(n14384), .A0(n13475), .A1(n13444) );
  nand02 U7444 ( .Y(n14388), .A0(s_exp_10_i_4_), .A1(n14387) );
  xor2 U7445 ( .Y(s_exp_10a_4_), .A0(s_exp_10_i_4_), .A1(n14387) );
  nand02 U7446 ( .Y(n14392), .A0(n13511), .A1(s_exp_10_i_0_) );
  inv01 U7447 ( .Y(n14389), .A(s_exp_10_i_2_) );
  nand03 U7448 ( .Y(n14390), .A0(s_exp_10_i_1_), .A1(s_exp_10_i_0_), .A2(
        n13512) );
  nand02 U7449 ( .Y(n____return6722_5_), .A0(n14393), .A1(n12267) );
  nand02 U7450 ( .Y(n14346), .A0(s_shr2_5_), .A1(n14372) );
  mux21 U7451 ( .Y(n14393), .A0(n14394), .A1(n12347), .S0(s_shr2_5_) );
  nor02 U7452 ( .Y(n14394), .A0(n14372), .A1(n12347) );
  nand02 U7453 ( .Y(n14395), .A0(n14396), .A1(n13556) );
  nor02 U7454 ( .Y(n14244), .A0(n14352), .A1(n14353) );
  nand02 U7455 ( .Y(n____return6722_3_), .A0(n14397), .A1(n13562) );
  nor02 U7456 ( .Y(n14263), .A0(n14352), .A1(s_shr2_2_) );
  mux21 U7457 ( .Y(n14397), .A0(s_shr2_3_), .A1(n13557), .S0(n13211) );
  nor02 U7458 ( .Y(n14246), .A0(n14353), .A1(s_shr2_3_) );
  nor02 U7459 ( .Y(n14396), .A0(n13582), .A1(n14398) );
  nand02 U7460 ( .Y(n14161), .A0(s_shr2_1_), .A1(s_shr2_0_) );
  nand02 U7461 ( .Y(n____return6722_1_), .A0(n9810), .A1(n13598) );
  or02 U7462 ( .Y(n14160), .A0(n14399), .A1(s_shr2_0_) );
  inv01 U7463 ( .Y(n14163), .A(n13518) );
  nand02 U7464 ( .Y(n14164), .A0(s_shr2_0_), .A1(n14399) );
  inv01 U7465 ( .Y(n14399), .A(s_shr2_1_) );
  post_norm_mul_DW01_inc_9_0 add_233_plus_plus ( .A(s_expo2b), .SUM({n7170_8_, 
        n____return7168_7_, n____return7168_6_, n____return7168_5_, 
        n____return7168_4_, n____return7168_3_, n____return7168_2_, 
        n____return7168_1_, n____return7168_0_}) );
  post_norm_mul_DW01_inc_25_0 add_222_plus_plus ( .A({s_frac2a_47_, n13520, 
        s_frac2a_45_, s_frac2a_44_, s_frac2a_43_, s_frac2a_42_, s_frac2a_41_, 
        s_frac2a_40_, s_frac2a_39_, s_frac2a_38_, s_frac2a_37_, s_frac2a_36_, 
        s_frac2a_35_, s_frac2a_34_, s_frac2a_33_, s_frac2a_32_, s_frac2a_31_, 
        s_frac2a_30_, s_frac2a_29_, s_frac2a_28_, s_frac2a_27_, s_frac2a_26_, 
        s_frac2a_25_, s_frac2a_24_, s_frac2a_23_}), .SUM({n____return7070_24_, 
        n7072_23_, n____return7070_22_, n____return7070_21_, 
        n____return7070_20_, n____return7070_19_, n____return7070_18_, 
        n____return7070_17_, n____return7070_16_, n____return7070_15_, 
        n____return7070_14_, n____return7070_13_, n____return7070_12_, 
        n____return7070_11_, n____return7070_10_, n____return7070_9_, 
        n____return7070_8_, n____return7070_7_, n____return7070_6_, 
        n____return7070_5_, n____return7070_4_, n____return7070_3_, 
        n____return7070_2_, n____return7070_1_, n____return7070_0_}) );
  post_norm_mul_DW01_dec_9_0 sub_192_minus_minus ( .A(s_expo1), .SUM({n6653_8_, 
        n____return6651_7_, n____return6651_6_, n____return6651_5_, 
        n____return6651_4_, n____return6651_3_, n____return6651_2_, 
        n____return6651_1_, n____return6651_0_}) );
  post_norm_mul_DW01_sub_7_0 r64 ( .A({1'b0, n12474, n12476, n12480, n12478, 
        n12472, n10296}), .B({U1086_U4_Z_6, n13444, n13475, n13458, n13455, 
        n13461, n13447}), .CI(1'b0), .DIFF({n____return6004_6_, 
        n____return5956_5_, n____return5956_4_, n____return5956_3_, 
        n____return5956_2_, n____return5956_1_, n____return5956_0_}) );
  post_norm_mul_DW01_sub_10_0 sub_141_minus_minus ( .A({n10407, n12774, n12808, 
        s_exp_10a_6_, n13444, n13475, n13459, n13456, n13462, n13446}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, s_zeros}), .CI(1'b0), .DIFF(s_exp_10b) );
  post_norm_mul_DW01_cmp2_6_0 gt_197_gt_gt ( .A({s_r_zeros_5_, s_r_zeros_4_, 
        s_r_zeros_3_, s_r_zeros_2_, s_r_zeros_1_, s_r_zeros_0_}), .B({
        n____return6722_5_, n12246, n____return6722_3_, n12365, 
        n____return6722_1_, n10403}), .LEQ(1'b0), .TC(1'b0), .LT_LE(
        n____return6760) );
endmodule


module pre_norm_div_DW01_sub_10_1 ( A, B, CI, DIFF, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] DIFF;
  input CI;
  output CO;
  wire   carry_9_, carry_8_, carry_7_, carry_5_, carry_4_, carry_3_, carry_2_,
         carry_1_, B_not_4_, B_not_3_, B_not_2_, B_not_1_, B_not_0_, n102, n6,
         n8, n10, n12, n14, n16, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101;

  buf02 U6 ( .Y(DIFF[4]), .A(n102) );
  xor2 U7 ( .Y(n6), .A0(B_not_0_), .A1(A[0]) );
  inv01 U8 ( .Y(DIFF[0]), .A(n6) );
  xor2 U9 ( .Y(n8), .A0(A[6]), .A1(n19) );
  inv01 U10 ( .Y(DIFF[6]), .A(n8) );
  xor2 U11 ( .Y(n10), .A0(A[8]), .A1(n21) );
  inv01 U12 ( .Y(DIFF[8]), .A(n10) );
  xor2 U13 ( .Y(n12), .A0(A[5]), .A1(n101) );
  inv01 U14 ( .Y(DIFF[5]), .A(n12) );
  xor2 U15 ( .Y(n14), .A0(A[7]), .A1(n20) );
  inv01 U16 ( .Y(DIFF[7]), .A(n14) );
  xor2 U17 ( .Y(n16), .A0(carry_9_), .A1(A[9]) );
  inv01 U18 ( .Y(DIFF[9]), .A(n16) );
  nor02 U19 ( .Y(n18), .A0(A[5]), .A1(n101) );
  inv02 U20 ( .Y(n19), .A(n18) );
  buf02 U21 ( .Y(n20), .A(carry_7_) );
  buf02 U22 ( .Y(n21), .A(carry_8_) );
  inv01 U23 ( .Y(DIFF[3]), .A(n22) );
  inv02 U24 ( .Y(carry_4_), .A(n23) );
  inv02 U25 ( .Y(n24), .A(B_not_3_) );
  inv02 U26 ( .Y(n25), .A(A[3]) );
  inv02 U27 ( .Y(n26), .A(carry_3_) );
  nor02 U28 ( .Y(n27), .A0(n24), .A1(n28) );
  nor02 U29 ( .Y(n29), .A0(n25), .A1(n30) );
  nor02 U30 ( .Y(n31), .A0(n26), .A1(n32) );
  nor02 U31 ( .Y(n33), .A0(n26), .A1(n34) );
  nor02 U32 ( .Y(n22), .A0(n35), .A1(n36) );
  nor02 U33 ( .Y(n37), .A0(n25), .A1(n26) );
  nor02 U34 ( .Y(n38), .A0(n24), .A1(n26) );
  nor02 U35 ( .Y(n39), .A0(n24), .A1(n25) );
  nor02 U36 ( .Y(n23), .A0(n39), .A1(n40) );
  nor02 U37 ( .Y(n41), .A0(A[3]), .A1(carry_3_) );
  inv01 U38 ( .Y(n28), .A(n41) );
  nor02 U39 ( .Y(n42), .A0(B_not_3_), .A1(carry_3_) );
  inv01 U40 ( .Y(n30), .A(n42) );
  nor02 U41 ( .Y(n43), .A0(B_not_3_), .A1(A[3]) );
  inv01 U42 ( .Y(n32), .A(n43) );
  nor02 U43 ( .Y(n44), .A0(n24), .A1(n25) );
  inv01 U44 ( .Y(n34), .A(n44) );
  nor02 U45 ( .Y(n45), .A0(n27), .A1(n29) );
  inv01 U46 ( .Y(n35), .A(n45) );
  nor02 U47 ( .Y(n46), .A0(n31), .A1(n33) );
  inv01 U48 ( .Y(n36), .A(n46) );
  nor02 U49 ( .Y(n47), .A0(n37), .A1(n38) );
  inv01 U50 ( .Y(n40), .A(n47) );
  inv02 U51 ( .Y(n48), .A(n79) );
  inv01 U52 ( .Y(DIFF[2]), .A(n49) );
  inv02 U53 ( .Y(carry_3_), .A(n50) );
  inv02 U54 ( .Y(n51), .A(B_not_2_) );
  inv02 U55 ( .Y(n52), .A(A[2]) );
  inv02 U56 ( .Y(n53), .A(carry_2_) );
  nor02 U57 ( .Y(n54), .A0(n51), .A1(n55) );
  nor02 U58 ( .Y(n56), .A0(n52), .A1(n57) );
  nor02 U59 ( .Y(n58), .A0(n53), .A1(n59) );
  nor02 U60 ( .Y(n60), .A0(n53), .A1(n61) );
  nor02 U61 ( .Y(n49), .A0(n62), .A1(n63) );
  nor02 U62 ( .Y(n64), .A0(n52), .A1(n53) );
  nor02 U63 ( .Y(n65), .A0(n51), .A1(n53) );
  nor02 U64 ( .Y(n66), .A0(n51), .A1(n52) );
  nor02 U65 ( .Y(n50), .A0(n66), .A1(n67) );
  nor02 U66 ( .Y(n68), .A0(A[2]), .A1(carry_2_) );
  inv01 U67 ( .Y(n55), .A(n68) );
  nor02 U68 ( .Y(n69), .A0(B_not_2_), .A1(carry_2_) );
  inv01 U69 ( .Y(n57), .A(n69) );
  nor02 U70 ( .Y(n70), .A0(B_not_2_), .A1(A[2]) );
  inv01 U71 ( .Y(n59), .A(n70) );
  nor02 U72 ( .Y(n71), .A0(n51), .A1(n52) );
  inv01 U73 ( .Y(n61), .A(n71) );
  nor02 U74 ( .Y(n72), .A0(n54), .A1(n56) );
  inv01 U75 ( .Y(n62), .A(n72) );
  nor02 U76 ( .Y(n73), .A0(n58), .A1(n60) );
  inv01 U77 ( .Y(n63), .A(n73) );
  nor02 U78 ( .Y(n74), .A0(n64), .A1(n65) );
  inv01 U79 ( .Y(n67), .A(n74) );
  inv01 U80 ( .Y(DIFF[1]), .A(n75) );
  inv02 U81 ( .Y(carry_2_), .A(n76) );
  inv02 U82 ( .Y(n77), .A(B_not_1_) );
  inv02 U83 ( .Y(n78), .A(A[1]) );
  inv02 U84 ( .Y(n79), .A(carry_1_) );
  nor02 U85 ( .Y(n80), .A0(n77), .A1(n81) );
  nor02 U86 ( .Y(n82), .A0(n78), .A1(n83) );
  nor02 U87 ( .Y(n84), .A0(n79), .A1(n85) );
  nor02 U88 ( .Y(n86), .A0(n79), .A1(n87) );
  nor02 U89 ( .Y(n75), .A0(n88), .A1(n89) );
  nor02 U90 ( .Y(n90), .A0(n78), .A1(n79) );
  nor02 U91 ( .Y(n91), .A0(n77), .A1(n79) );
  nor02 U92 ( .Y(n92), .A0(n77), .A1(n78) );
  nor02 U93 ( .Y(n76), .A0(n92), .A1(n93) );
  nor02 U94 ( .Y(n94), .A0(A[1]), .A1(carry_1_) );
  inv01 U95 ( .Y(n81), .A(n94) );
  nor02 U96 ( .Y(n95), .A0(B_not_1_), .A1(n48) );
  inv01 U97 ( .Y(n83), .A(n95) );
  nor02 U98 ( .Y(n96), .A0(B_not_1_), .A1(A[1]) );
  inv01 U99 ( .Y(n85), .A(n96) );
  nor02 U100 ( .Y(n97), .A0(n77), .A1(n78) );
  inv01 U101 ( .Y(n87), .A(n97) );
  nor02 U102 ( .Y(n98), .A0(n80), .A1(n82) );
  inv01 U103 ( .Y(n88), .A(n98) );
  nor02 U104 ( .Y(n99), .A0(n84), .A1(n86) );
  inv01 U105 ( .Y(n89), .A(n99) );
  nor02 U106 ( .Y(n100), .A0(n90), .A1(n91) );
  inv01 U107 ( .Y(n93), .A(n100) );
  buf02 U108 ( .Y(n101), .A(carry_5_) );
  inv02 U109 ( .Y(B_not_0_), .A(B[0]) );
  inv02 U110 ( .Y(B_not_3_), .A(B[3]) );
  inv02 U111 ( .Y(B_not_1_), .A(B[1]) );
  inv02 U112 ( .Y(B_not_2_), .A(B[2]) );
  inv02 U113 ( .Y(B_not_4_), .A(B[4]) );
  or02 U114 ( .Y(carry_9_), .A0(A[8]), .A1(n21) );
  or02 U115 ( .Y(carry_8_), .A0(A[7]), .A1(n20) );
  or02 U116 ( .Y(carry_7_), .A0(A[6]), .A1(n19) );
  or02 U117 ( .Y(carry_1_), .A0(B_not_0_), .A1(A[0]) );
  fadd1 U2_4 ( .S(n102), .CO(carry_5_), .A(A[4]), .B(B_not_4_), .CI(carry_4_)
         );
endmodule


module pre_norm_div_DW01_add_10_1 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   carry_9_, carry_8_, carry_7_, carry_6_, carry_5_, carry_4_, carry_3_,
         carry_2_, carry_1_, n212, n213, n2, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211;

  buf02 U4 ( .Y(SUM[9]), .A(n212) );
  and02 U5 ( .Y(n2), .A0(A[0]), .A1(B[0]) );
  buf02 U6 ( .Y(SUM[0]), .A(n213) );
  inv02 U7 ( .Y(SUM[7]), .A(n4) );
  inv02 U8 ( .Y(carry_8_), .A(n5) );
  inv02 U9 ( .Y(n6), .A(B[7]) );
  inv02 U10 ( .Y(n7), .A(A[7]) );
  inv02 U11 ( .Y(n8), .A(carry_7_) );
  nor02 U12 ( .Y(n9), .A0(n6), .A1(n10) );
  nor02 U13 ( .Y(n11), .A0(n7), .A1(n12) );
  nor02 U14 ( .Y(n13), .A0(n8), .A1(n14) );
  nor02 U15 ( .Y(n15), .A0(n8), .A1(n16) );
  nor02 U16 ( .Y(n4), .A0(n17), .A1(n18) );
  nor02 U17 ( .Y(n19), .A0(n7), .A1(n8) );
  nor02 U18 ( .Y(n20), .A0(n6), .A1(n8) );
  nor02 U19 ( .Y(n21), .A0(n6), .A1(n7) );
  nor02 U20 ( .Y(n5), .A0(n21), .A1(n22) );
  nor02 U21 ( .Y(n23), .A0(A[7]), .A1(carry_7_) );
  inv01 U22 ( .Y(n10), .A(n23) );
  nor02 U23 ( .Y(n24), .A0(B[7]), .A1(carry_7_) );
  inv01 U24 ( .Y(n12), .A(n24) );
  nor02 U25 ( .Y(n25), .A0(B[7]), .A1(A[7]) );
  inv01 U26 ( .Y(n14), .A(n25) );
  nor02 U27 ( .Y(n26), .A0(n6), .A1(n7) );
  inv01 U28 ( .Y(n16), .A(n26) );
  nor02 U29 ( .Y(n27), .A0(n9), .A1(n11) );
  inv01 U30 ( .Y(n17), .A(n27) );
  nor02 U31 ( .Y(n28), .A0(n13), .A1(n15) );
  inv01 U32 ( .Y(n18), .A(n28) );
  nor02 U33 ( .Y(n29), .A0(n19), .A1(n20) );
  inv01 U34 ( .Y(n22), .A(n29) );
  inv02 U35 ( .Y(SUM[8]), .A(n30) );
  inv02 U36 ( .Y(carry_9_), .A(n31) );
  inv02 U37 ( .Y(n32), .A(B[8]) );
  inv02 U38 ( .Y(n33), .A(A[8]) );
  inv02 U39 ( .Y(n34), .A(carry_8_) );
  nor02 U40 ( .Y(n35), .A0(n32), .A1(n36) );
  nor02 U41 ( .Y(n37), .A0(n33), .A1(n38) );
  nor02 U42 ( .Y(n39), .A0(n34), .A1(n40) );
  nor02 U43 ( .Y(n41), .A0(n34), .A1(n42) );
  nor02 U44 ( .Y(n30), .A0(n43), .A1(n44) );
  nor02 U45 ( .Y(n45), .A0(n33), .A1(n34) );
  nor02 U46 ( .Y(n46), .A0(n32), .A1(n34) );
  nor02 U47 ( .Y(n47), .A0(n32), .A1(n33) );
  nor02 U48 ( .Y(n31), .A0(n47), .A1(n48) );
  nor02 U49 ( .Y(n49), .A0(A[8]), .A1(carry_8_) );
  inv01 U50 ( .Y(n36), .A(n49) );
  nor02 U51 ( .Y(n50), .A0(B[8]), .A1(carry_8_) );
  inv01 U52 ( .Y(n38), .A(n50) );
  nor02 U53 ( .Y(n51), .A0(B[8]), .A1(A[8]) );
  inv01 U54 ( .Y(n40), .A(n51) );
  nor02 U55 ( .Y(n52), .A0(n32), .A1(n33) );
  inv01 U56 ( .Y(n42), .A(n52) );
  nor02 U57 ( .Y(n53), .A0(n35), .A1(n37) );
  inv01 U58 ( .Y(n43), .A(n53) );
  nor02 U59 ( .Y(n54), .A0(n39), .A1(n41) );
  inv01 U60 ( .Y(n44), .A(n54) );
  nor02 U61 ( .Y(n55), .A0(n45), .A1(n46) );
  inv01 U62 ( .Y(n48), .A(n55) );
  inv02 U63 ( .Y(SUM[5]), .A(n56) );
  inv02 U64 ( .Y(carry_6_), .A(n57) );
  inv02 U65 ( .Y(n58), .A(B[5]) );
  inv02 U66 ( .Y(n59), .A(A[5]) );
  inv02 U67 ( .Y(n60), .A(carry_5_) );
  nor02 U68 ( .Y(n61), .A0(n58), .A1(n62) );
  nor02 U69 ( .Y(n63), .A0(n59), .A1(n64) );
  nor02 U70 ( .Y(n65), .A0(n60), .A1(n66) );
  nor02 U71 ( .Y(n67), .A0(n60), .A1(n68) );
  nor02 U72 ( .Y(n56), .A0(n69), .A1(n70) );
  nor02 U73 ( .Y(n71), .A0(n59), .A1(n60) );
  nor02 U74 ( .Y(n72), .A0(n58), .A1(n60) );
  nor02 U75 ( .Y(n73), .A0(n58), .A1(n59) );
  nor02 U76 ( .Y(n57), .A0(n73), .A1(n74) );
  nor02 U77 ( .Y(n75), .A0(A[5]), .A1(carry_5_) );
  inv01 U78 ( .Y(n62), .A(n75) );
  nor02 U79 ( .Y(n76), .A0(B[5]), .A1(carry_5_) );
  inv01 U80 ( .Y(n64), .A(n76) );
  nor02 U81 ( .Y(n77), .A0(B[5]), .A1(A[5]) );
  inv01 U82 ( .Y(n66), .A(n77) );
  nor02 U83 ( .Y(n78), .A0(n58), .A1(n59) );
  inv01 U84 ( .Y(n68), .A(n78) );
  nor02 U85 ( .Y(n79), .A0(n61), .A1(n63) );
  inv01 U86 ( .Y(n69), .A(n79) );
  nor02 U87 ( .Y(n80), .A0(n65), .A1(n67) );
  inv01 U88 ( .Y(n70), .A(n80) );
  nor02 U89 ( .Y(n81), .A0(n71), .A1(n72) );
  inv01 U90 ( .Y(n74), .A(n81) );
  inv02 U91 ( .Y(SUM[6]), .A(n82) );
  inv02 U92 ( .Y(carry_7_), .A(n83) );
  inv02 U93 ( .Y(n84), .A(B[6]) );
  inv02 U94 ( .Y(n85), .A(A[6]) );
  inv02 U95 ( .Y(n86), .A(carry_6_) );
  nor02 U96 ( .Y(n87), .A0(n84), .A1(n88) );
  nor02 U97 ( .Y(n89), .A0(n85), .A1(n90) );
  nor02 U98 ( .Y(n91), .A0(n86), .A1(n92) );
  nor02 U99 ( .Y(n93), .A0(n86), .A1(n94) );
  nor02 U100 ( .Y(n82), .A0(n95), .A1(n96) );
  nor02 U101 ( .Y(n97), .A0(n85), .A1(n86) );
  nor02 U102 ( .Y(n98), .A0(n84), .A1(n86) );
  nor02 U103 ( .Y(n99), .A0(n84), .A1(n85) );
  nor02 U104 ( .Y(n83), .A0(n99), .A1(n100) );
  nor02 U105 ( .Y(n101), .A0(A[6]), .A1(carry_6_) );
  inv01 U106 ( .Y(n88), .A(n101) );
  nor02 U107 ( .Y(n102), .A0(B[6]), .A1(carry_6_) );
  inv01 U108 ( .Y(n90), .A(n102) );
  nor02 U109 ( .Y(n103), .A0(B[6]), .A1(A[6]) );
  inv01 U110 ( .Y(n92), .A(n103) );
  nor02 U111 ( .Y(n104), .A0(n84), .A1(n85) );
  inv01 U112 ( .Y(n94), .A(n104) );
  nor02 U113 ( .Y(n105), .A0(n87), .A1(n89) );
  inv01 U114 ( .Y(n95), .A(n105) );
  nor02 U115 ( .Y(n106), .A0(n91), .A1(n93) );
  inv01 U116 ( .Y(n96), .A(n106) );
  nor02 U117 ( .Y(n107), .A0(n97), .A1(n98) );
  inv01 U118 ( .Y(n100), .A(n107) );
  inv02 U119 ( .Y(SUM[4]), .A(n108) );
  inv02 U120 ( .Y(carry_5_), .A(n109) );
  inv02 U121 ( .Y(n110), .A(B[4]) );
  inv02 U122 ( .Y(n111), .A(A[4]) );
  inv02 U123 ( .Y(n112), .A(carry_4_) );
  nor02 U124 ( .Y(n113), .A0(n110), .A1(n114) );
  nor02 U125 ( .Y(n115), .A0(n111), .A1(n116) );
  nor02 U126 ( .Y(n117), .A0(n112), .A1(n118) );
  nor02 U127 ( .Y(n119), .A0(n112), .A1(n120) );
  nor02 U128 ( .Y(n108), .A0(n121), .A1(n122) );
  nor02 U129 ( .Y(n123), .A0(n111), .A1(n112) );
  nor02 U130 ( .Y(n124), .A0(n110), .A1(n112) );
  nor02 U131 ( .Y(n125), .A0(n110), .A1(n111) );
  nor02 U132 ( .Y(n109), .A0(n125), .A1(n126) );
  nor02 U133 ( .Y(n127), .A0(A[4]), .A1(carry_4_) );
  inv01 U134 ( .Y(n114), .A(n127) );
  nor02 U135 ( .Y(n128), .A0(B[4]), .A1(carry_4_) );
  inv01 U136 ( .Y(n116), .A(n128) );
  nor02 U137 ( .Y(n129), .A0(B[4]), .A1(A[4]) );
  inv01 U138 ( .Y(n118), .A(n129) );
  nor02 U139 ( .Y(n130), .A0(n110), .A1(n111) );
  inv01 U140 ( .Y(n120), .A(n130) );
  nor02 U141 ( .Y(n131), .A0(n113), .A1(n115) );
  inv01 U142 ( .Y(n121), .A(n131) );
  nor02 U143 ( .Y(n132), .A0(n117), .A1(n119) );
  inv01 U144 ( .Y(n122), .A(n132) );
  nor02 U145 ( .Y(n133), .A0(n123), .A1(n124) );
  inv01 U146 ( .Y(n126), .A(n133) );
  inv02 U147 ( .Y(SUM[3]), .A(n134) );
  inv02 U148 ( .Y(carry_4_), .A(n135) );
  inv02 U149 ( .Y(n136), .A(B[3]) );
  inv02 U150 ( .Y(n137), .A(A[3]) );
  inv02 U151 ( .Y(n138), .A(carry_3_) );
  nor02 U152 ( .Y(n139), .A0(n136), .A1(n140) );
  nor02 U153 ( .Y(n141), .A0(n137), .A1(n142) );
  nor02 U154 ( .Y(n143), .A0(n138), .A1(n144) );
  nor02 U155 ( .Y(n145), .A0(n138), .A1(n146) );
  nor02 U156 ( .Y(n134), .A0(n147), .A1(n148) );
  nor02 U157 ( .Y(n149), .A0(n137), .A1(n138) );
  nor02 U158 ( .Y(n150), .A0(n136), .A1(n138) );
  nor02 U159 ( .Y(n151), .A0(n136), .A1(n137) );
  nor02 U160 ( .Y(n135), .A0(n151), .A1(n152) );
  nor02 U161 ( .Y(n153), .A0(A[3]), .A1(carry_3_) );
  inv01 U162 ( .Y(n140), .A(n153) );
  nor02 U163 ( .Y(n154), .A0(B[3]), .A1(carry_3_) );
  inv01 U164 ( .Y(n142), .A(n154) );
  nor02 U165 ( .Y(n155), .A0(B[3]), .A1(A[3]) );
  inv01 U166 ( .Y(n144), .A(n155) );
  nor02 U167 ( .Y(n156), .A0(n136), .A1(n137) );
  inv01 U168 ( .Y(n146), .A(n156) );
  nor02 U169 ( .Y(n157), .A0(n139), .A1(n141) );
  inv01 U170 ( .Y(n147), .A(n157) );
  nor02 U171 ( .Y(n158), .A0(n143), .A1(n145) );
  inv01 U172 ( .Y(n148), .A(n158) );
  nor02 U173 ( .Y(n159), .A0(n149), .A1(n150) );
  inv01 U174 ( .Y(n152), .A(n159) );
  inv02 U175 ( .Y(SUM[2]), .A(n160) );
  inv02 U176 ( .Y(carry_3_), .A(n161) );
  inv02 U177 ( .Y(n162), .A(B[2]) );
  inv02 U178 ( .Y(n163), .A(A[2]) );
  inv02 U179 ( .Y(n164), .A(carry_2_) );
  nor02 U180 ( .Y(n165), .A0(n162), .A1(n166) );
  nor02 U181 ( .Y(n167), .A0(n163), .A1(n168) );
  nor02 U182 ( .Y(n169), .A0(n164), .A1(n170) );
  nor02 U183 ( .Y(n171), .A0(n164), .A1(n172) );
  nor02 U184 ( .Y(n160), .A0(n173), .A1(n174) );
  nor02 U185 ( .Y(n175), .A0(n163), .A1(n164) );
  nor02 U186 ( .Y(n176), .A0(n162), .A1(n164) );
  nor02 U187 ( .Y(n177), .A0(n162), .A1(n163) );
  nor02 U188 ( .Y(n161), .A0(n177), .A1(n178) );
  nor02 U189 ( .Y(n179), .A0(A[2]), .A1(carry_2_) );
  inv01 U190 ( .Y(n166), .A(n179) );
  nor02 U191 ( .Y(n180), .A0(B[2]), .A1(carry_2_) );
  inv01 U192 ( .Y(n168), .A(n180) );
  nor02 U193 ( .Y(n181), .A0(B[2]), .A1(A[2]) );
  inv01 U194 ( .Y(n170), .A(n181) );
  nor02 U195 ( .Y(n182), .A0(n162), .A1(n163) );
  inv01 U196 ( .Y(n172), .A(n182) );
  nor02 U197 ( .Y(n183), .A0(n165), .A1(n167) );
  inv01 U198 ( .Y(n173), .A(n183) );
  nor02 U199 ( .Y(n184), .A0(n169), .A1(n171) );
  inv01 U200 ( .Y(n174), .A(n184) );
  nor02 U201 ( .Y(n185), .A0(n175), .A1(n176) );
  inv01 U202 ( .Y(n178), .A(n185) );
  inv02 U203 ( .Y(SUM[1]), .A(n186) );
  inv02 U204 ( .Y(carry_2_), .A(n187) );
  inv02 U205 ( .Y(n188), .A(B[1]) );
  inv02 U206 ( .Y(n189), .A(A[1]) );
  inv02 U207 ( .Y(n190), .A(carry_1_) );
  nor02 U208 ( .Y(n191), .A0(n188), .A1(n192) );
  nor02 U209 ( .Y(n193), .A0(n189), .A1(n194) );
  nor02 U210 ( .Y(n195), .A0(n190), .A1(n196) );
  nor02 U211 ( .Y(n197), .A0(n190), .A1(n198) );
  nor02 U212 ( .Y(n186), .A0(n199), .A1(n200) );
  nor02 U213 ( .Y(n201), .A0(n189), .A1(n190) );
  nor02 U214 ( .Y(n202), .A0(n188), .A1(n190) );
  nor02 U215 ( .Y(n203), .A0(n188), .A1(n189) );
  nor02 U216 ( .Y(n187), .A0(n203), .A1(n204) );
  nor02 U217 ( .Y(n205), .A0(A[1]), .A1(n2) );
  inv01 U218 ( .Y(n192), .A(n205) );
  nor02 U219 ( .Y(n206), .A0(B[1]), .A1(n2) );
  inv01 U220 ( .Y(n194), .A(n206) );
  nor02 U221 ( .Y(n207), .A0(B[1]), .A1(A[1]) );
  inv01 U222 ( .Y(n196), .A(n207) );
  nor02 U223 ( .Y(n208), .A0(n188), .A1(n189) );
  inv01 U224 ( .Y(n198), .A(n208) );
  nor02 U225 ( .Y(n209), .A0(n191), .A1(n193) );
  inv01 U226 ( .Y(n199), .A(n209) );
  nor02 U227 ( .Y(n210), .A0(n195), .A1(n197) );
  inv01 U228 ( .Y(n200), .A(n210) );
  nor02 U229 ( .Y(n211), .A0(n201), .A1(n202) );
  inv01 U230 ( .Y(n204), .A(n211) );
  and02 U231 ( .Y(carry_1_), .A0(A[0]), .A1(B[0]) );
  xor2 U232 ( .Y(n213), .A0(B[0]), .A1(A[0]) );
  fadd1 U1_9 ( .S(n212), .A(A[9]), .B(B[9]), .CI(carry_9_) );
endmodule


module pre_norm_div_DW01_sub_10_0 ( A, B, CI, DIFF, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] DIFF;
  input CI;
  output CO;
  wire   carry_9_, carry_5_, carry_4_, carry_3_, carry_2_, n124, n125, n126,
         n127, n128, n5, n6, n7, n8, n9, n10, n15, n16, n18, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123;
  wire   [9:0] B_not;

  nand02 U6 ( .Y(n5), .A0(n8), .A1(B_not[7]) );
  inv02 U7 ( .Y(n6), .A(n5) );
  nand02 U8 ( .Y(n7), .A0(n10), .A1(B_not[6]) );
  inv02 U9 ( .Y(n8), .A(n7) );
  nand02 U10 ( .Y(n9), .A0(carry_5_), .A1(B_not[5]) );
  inv02 U11 ( .Y(n10), .A(n9) );
  buf02 U12 ( .Y(DIFF[5]), .A(n128) );
  buf02 U13 ( .Y(DIFF[7]), .A(n126) );
  buf02 U14 ( .Y(DIFF[8]), .A(n125) );
  buf02 U15 ( .Y(DIFF[6]), .A(n127) );
  nor02 U16 ( .Y(n15), .A0(B_not[0]), .A1(A[0]) );
  inv02 U17 ( .Y(n16), .A(n15) );
  buf02 U18 ( .Y(DIFF[9]), .A(n124) );
  xor2 U19 ( .Y(n18), .A0(B_not[0]), .A1(A[0]) );
  inv02 U20 ( .Y(DIFF[0]), .A(n18) );
  inv02 U21 ( .Y(DIFF[4]), .A(n20) );
  inv02 U22 ( .Y(carry_5_), .A(n21) );
  inv02 U23 ( .Y(n22), .A(B_not[4]) );
  inv02 U24 ( .Y(n23), .A(A[4]) );
  inv02 U25 ( .Y(n24), .A(carry_4_) );
  nor02 U26 ( .Y(n25), .A0(n22), .A1(n26) );
  nor02 U27 ( .Y(n27), .A0(n23), .A1(n28) );
  nor02 U28 ( .Y(n29), .A0(n24), .A1(n30) );
  nor02 U29 ( .Y(n31), .A0(n24), .A1(n32) );
  nor02 U30 ( .Y(n20), .A0(n33), .A1(n34) );
  nor02 U31 ( .Y(n35), .A0(n23), .A1(n24) );
  nor02 U32 ( .Y(n36), .A0(n22), .A1(n24) );
  nor02 U33 ( .Y(n37), .A0(n22), .A1(n23) );
  nor02 U34 ( .Y(n21), .A0(n37), .A1(n38) );
  nor02 U35 ( .Y(n39), .A0(A[4]), .A1(carry_4_) );
  inv01 U36 ( .Y(n26), .A(n39) );
  nor02 U37 ( .Y(n40), .A0(B_not[4]), .A1(carry_4_) );
  inv01 U38 ( .Y(n28), .A(n40) );
  nor02 U39 ( .Y(n41), .A0(B_not[4]), .A1(A[4]) );
  inv01 U40 ( .Y(n30), .A(n41) );
  nor02 U41 ( .Y(n42), .A0(n22), .A1(n23) );
  inv01 U42 ( .Y(n32), .A(n42) );
  nor02 U43 ( .Y(n43), .A0(n25), .A1(n27) );
  inv01 U44 ( .Y(n33), .A(n43) );
  nor02 U45 ( .Y(n44), .A0(n29), .A1(n31) );
  inv01 U46 ( .Y(n34), .A(n44) );
  nor02 U47 ( .Y(n45), .A0(n35), .A1(n36) );
  inv01 U48 ( .Y(n38), .A(n45) );
  inv02 U49 ( .Y(B_not[4]), .A(B[4]) );
  inv02 U50 ( .Y(DIFF[3]), .A(n46) );
  inv02 U51 ( .Y(carry_4_), .A(n47) );
  inv02 U52 ( .Y(n48), .A(B_not[3]) );
  inv02 U53 ( .Y(n49), .A(A[3]) );
  inv02 U54 ( .Y(n50), .A(carry_3_) );
  nor02 U55 ( .Y(n51), .A0(n48), .A1(n52) );
  nor02 U56 ( .Y(n53), .A0(n49), .A1(n54) );
  nor02 U57 ( .Y(n55), .A0(n50), .A1(n56) );
  nor02 U58 ( .Y(n57), .A0(n50), .A1(n58) );
  nor02 U59 ( .Y(n46), .A0(n59), .A1(n60) );
  nor02 U60 ( .Y(n61), .A0(n49), .A1(n50) );
  nor02 U61 ( .Y(n62), .A0(n48), .A1(n50) );
  nor02 U62 ( .Y(n63), .A0(n48), .A1(n49) );
  nor02 U63 ( .Y(n47), .A0(n63), .A1(n64) );
  nor02 U64 ( .Y(n65), .A0(A[3]), .A1(carry_3_) );
  inv01 U65 ( .Y(n52), .A(n65) );
  nor02 U66 ( .Y(n66), .A0(B_not[3]), .A1(carry_3_) );
  inv01 U67 ( .Y(n54), .A(n66) );
  nor02 U68 ( .Y(n67), .A0(B_not[3]), .A1(A[3]) );
  inv01 U69 ( .Y(n56), .A(n67) );
  nor02 U70 ( .Y(n68), .A0(n48), .A1(n49) );
  inv01 U71 ( .Y(n58), .A(n68) );
  nor02 U72 ( .Y(n69), .A0(n51), .A1(n53) );
  inv01 U73 ( .Y(n59), .A(n69) );
  nor02 U74 ( .Y(n70), .A0(n55), .A1(n57) );
  inv01 U75 ( .Y(n60), .A(n70) );
  nor02 U76 ( .Y(n71), .A0(n61), .A1(n62) );
  inv01 U77 ( .Y(n64), .A(n71) );
  inv02 U78 ( .Y(B_not[3]), .A(B[3]) );
  inv02 U79 ( .Y(DIFF[2]), .A(n72) );
  inv02 U80 ( .Y(carry_3_), .A(n73) );
  inv02 U81 ( .Y(n74), .A(B_not[2]) );
  inv02 U82 ( .Y(n75), .A(A[2]) );
  inv02 U83 ( .Y(n76), .A(carry_2_) );
  nor02 U84 ( .Y(n77), .A0(n74), .A1(n78) );
  nor02 U85 ( .Y(n79), .A0(n75), .A1(n80) );
  nor02 U86 ( .Y(n81), .A0(n76), .A1(n82) );
  nor02 U87 ( .Y(n83), .A0(n76), .A1(n84) );
  nor02 U88 ( .Y(n72), .A0(n85), .A1(n86) );
  nor02 U89 ( .Y(n87), .A0(n75), .A1(n76) );
  nor02 U90 ( .Y(n88), .A0(n74), .A1(n76) );
  nor02 U91 ( .Y(n89), .A0(n74), .A1(n75) );
  nor02 U92 ( .Y(n73), .A0(n89), .A1(n90) );
  nor02 U93 ( .Y(n91), .A0(A[2]), .A1(carry_2_) );
  inv01 U94 ( .Y(n78), .A(n91) );
  nor02 U95 ( .Y(n92), .A0(B_not[2]), .A1(carry_2_) );
  inv01 U96 ( .Y(n80), .A(n92) );
  nor02 U97 ( .Y(n93), .A0(B_not[2]), .A1(A[2]) );
  inv01 U98 ( .Y(n82), .A(n93) );
  nor02 U99 ( .Y(n94), .A0(n74), .A1(n75) );
  inv01 U100 ( .Y(n84), .A(n94) );
  nor02 U101 ( .Y(n95), .A0(n77), .A1(n79) );
  inv01 U102 ( .Y(n85), .A(n95) );
  nor02 U103 ( .Y(n96), .A0(n81), .A1(n83) );
  inv01 U104 ( .Y(n86), .A(n96) );
  nor02 U105 ( .Y(n97), .A0(n87), .A1(n88) );
  inv01 U106 ( .Y(n90), .A(n97) );
  inv02 U107 ( .Y(B_not[2]), .A(B[2]) );
  inv02 U108 ( .Y(DIFF[1]), .A(n98) );
  inv02 U109 ( .Y(carry_2_), .A(n99) );
  inv02 U110 ( .Y(n100), .A(B_not[1]) );
  inv02 U111 ( .Y(n101), .A(A[1]) );
  inv02 U112 ( .Y(n102), .A(n16) );
  nor02 U113 ( .Y(n103), .A0(n100), .A1(n104) );
  nor02 U114 ( .Y(n105), .A0(n101), .A1(n106) );
  nor02 U115 ( .Y(n107), .A0(n102), .A1(n108) );
  nor02 U116 ( .Y(n109), .A0(n102), .A1(n110) );
  nor02 U117 ( .Y(n98), .A0(n111), .A1(n112) );
  nor02 U118 ( .Y(n113), .A0(n101), .A1(n102) );
  nor02 U119 ( .Y(n114), .A0(n100), .A1(n102) );
  nor02 U120 ( .Y(n115), .A0(n100), .A1(n101) );
  nor02 U121 ( .Y(n99), .A0(n115), .A1(n116) );
  nor02 U122 ( .Y(n117), .A0(A[1]), .A1(n16) );
  inv01 U123 ( .Y(n104), .A(n117) );
  nor02 U124 ( .Y(n118), .A0(B_not[1]), .A1(n16) );
  inv01 U125 ( .Y(n106), .A(n118) );
  nor02 U126 ( .Y(n119), .A0(B_not[1]), .A1(A[1]) );
  inv01 U127 ( .Y(n108), .A(n119) );
  nor02 U128 ( .Y(n120), .A0(n100), .A1(n101) );
  inv01 U129 ( .Y(n110), .A(n120) );
  nor02 U130 ( .Y(n121), .A0(n103), .A1(n105) );
  inv01 U131 ( .Y(n111), .A(n121) );
  nor02 U132 ( .Y(n122), .A0(n107), .A1(n109) );
  inv01 U133 ( .Y(n112), .A(n122) );
  nor02 U134 ( .Y(n123), .A0(n113), .A1(n114) );
  inv01 U135 ( .Y(n116), .A(n123) );
  inv02 U136 ( .Y(B_not[1]), .A(B[1]) );
  xor2 U137 ( .Y(n124), .A0(B_not[9]), .A1(carry_9_) );
  and02 U138 ( .Y(carry_9_), .A0(n6), .A1(B_not[8]) );
  xor2 U139 ( .Y(n125), .A0(B_not[8]), .A1(n6) );
  xor2 U140 ( .Y(n126), .A0(B_not[7]), .A1(n8) );
  xor2 U141 ( .Y(n127), .A0(B_not[6]), .A1(n10) );
  xor2 U142 ( .Y(n128), .A0(B_not[5]), .A1(carry_5_) );
  inv04 U143 ( .Y(B_not[9]), .A(B[9]) );
  inv04 U144 ( .Y(B_not[8]), .A(B[8]) );
  inv04 U145 ( .Y(B_not[7]), .A(B[7]) );
  inv04 U146 ( .Y(B_not[6]), .A(B[6]) );
  inv04 U147 ( .Y(B_not[5]), .A(B[5]) );
  inv04 U148 ( .Y(B_not[0]), .A(B[0]) );
endmodule


module pre_norm_div ( clk_i, opa_i, opb_i, exp_10_o, dvdnd_50_o, dvsor_27_o );
  input [31:0] opa_i;
  input [31:0] opb_i;
  output [9:0] exp_10_o;
  output [49:0] dvdnd_50_o;
  output [26:0] dvsor_27_o;
  input clk_i;
  wire   n6466, n6467, n6468, n6469, n6470, n6471, s_dvd_zeros_4_,
         s_dvd_zeros_3_, s_dvd_zeros_2_, s_dvd_zeros_1_, s_dvd_zeros_0_,
         s_div_zeros_4_, s_div_zeros_3_, s_div_zeros_2_, s_div_zeros_1_,
         s_div_zeros_0_, n____return3431_0_, s_expa_in_8_, s_expa_in_7_,
         s_expa_in_6_, s_expa_in_5_, s_expa_in_4_, s_expa_in_3_, s_expa_in_2_,
         s_expa_in_1_, s_expa_in_0_, n____return3477_0_, s_expb_in_9_,
         s_expb_in_8_, s_expb_in_7_, s_expb_in_6_, s_expb_in_5_, s_expb_in_4_,
         s_expb_in_3_, s_expb_in_2_, s_expb_in_1_, s_expb_in_0_, n3654_8_,
         n____return3652_9_, n____return3652_7_, n____return3652_6_,
         n____return3652_5_, n____return3652_4_, n____return3652_3_,
         n____return3652_2_, n____return3652_1_, n____return3652_0_,
         n____return3612_9_, n____return3612_8_, n____return3612_7_,
         n____return3612_6_, n____return3612_5_, n____return3612_4_,
         n____return3612_3_, n____return3612_2_, n____return3612_1_,
         n____return3612_0_, n____return3578_9_, n____return3578_8_,
         n____return3578_7_, n____return3578_6_, n____return3578_5_,
         n____return3578_4_, n____return3578_3_, n____return3578_2_,
         n____return3578_1_, n____return3578_0_, n____return3540_6_,
         n____return3540_5_, n____return3540_4_, n____return3540_3_,
         n____return3540_2_, n____return3540_1_, n____return3540_0_, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4369, n4371, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4391,
         n4392, n4394, n4396, n4398, n4400, n4401, n4403, n4405, n4407, n4409,
         n4410, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5089, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465;
  wire   [9:0] s_exp_10_o;
  assign dvdnd_50_o[25] = 1'b0;
  assign dvdnd_50_o[24] = 1'b0;
  assign dvdnd_50_o[23] = 1'b0;
  assign dvdnd_50_o[22] = 1'b0;
  assign dvdnd_50_o[21] = 1'b0;
  assign dvdnd_50_o[20] = 1'b0;
  assign dvdnd_50_o[19] = 1'b0;
  assign dvdnd_50_o[18] = 1'b0;
  assign dvdnd_50_o[17] = 1'b0;
  assign dvdnd_50_o[16] = 1'b0;
  assign dvdnd_50_o[15] = 1'b0;
  assign dvdnd_50_o[14] = 1'b0;
  assign dvdnd_50_o[13] = 1'b0;
  assign dvdnd_50_o[12] = 1'b0;
  assign dvdnd_50_o[11] = 1'b0;
  assign dvdnd_50_o[10] = 1'b0;
  assign dvdnd_50_o[9] = 1'b0;
  assign dvdnd_50_o[8] = 1'b0;
  assign dvdnd_50_o[7] = 1'b0;
  assign dvdnd_50_o[6] = 1'b0;
  assign dvdnd_50_o[5] = 1'b0;
  assign dvdnd_50_o[4] = 1'b0;
  assign dvdnd_50_o[3] = 1'b0;
  assign dvdnd_50_o[2] = 1'b0;
  assign dvdnd_50_o[1] = 1'b0;
  assign dvdnd_50_o[0] = 1'b0;
  assign dvsor_27_o[26] = 1'b0;
  assign dvsor_27_o[25] = 1'b0;
  assign dvsor_27_o[24] = 1'b0;

  dff s_expa_in_reg_9_ ( .QB(n6465), .D(1'b0), .CLK(clk_i) );
  dff s_expb_in_reg_9_ ( .Q(s_expb_in_9_), .D(1'b0), .CLK(clk_i) );
  dff exp_10_o_reg_9_ ( .Q(exp_10_o[9]), .D(s_exp_10_o[9]), .CLK(clk_i) );
  dff exp_10_o_reg_8_ ( .Q(exp_10_o[8]), .D(s_exp_10_o[8]), .CLK(clk_i) );
  dff exp_10_o_reg_7_ ( .Q(exp_10_o[7]), .D(s_exp_10_o[7]), .CLK(clk_i) );
  dff exp_10_o_reg_6_ ( .Q(exp_10_o[6]), .D(s_exp_10_o[6]), .CLK(clk_i) );
  dff exp_10_o_reg_5_ ( .Q(exp_10_o[5]), .D(s_exp_10_o[5]), .CLK(clk_i) );
  dff exp_10_o_reg_4_ ( .Q(exp_10_o[4]), .D(s_exp_10_o[4]), .CLK(clk_i) );
  dff exp_10_o_reg_3_ ( .Q(exp_10_o[3]), .D(s_exp_10_o[3]), .CLK(clk_i) );
  dff exp_10_o_reg_2_ ( .Q(exp_10_o[2]), .D(s_exp_10_o[2]), .CLK(clk_i) );
  dff exp_10_o_reg_1_ ( .Q(exp_10_o[1]), .D(s_exp_10_o[1]), .CLK(clk_i) );
  dff exp_10_o_reg_0_ ( .Q(exp_10_o[0]), .D(s_exp_10_o[0]), .CLK(clk_i) );
  dff s_expa_in_reg_8_ ( .Q(s_expa_in_8_), .D(1'b0), .CLK(clk_i) );
  dff s_expa_in_reg_7_ ( .Q(s_expa_in_7_), .D(opa_i[30]), .CLK(clk_i) );
  dff s_expa_in_reg_6_ ( .Q(s_expa_in_6_), .D(opa_i[29]), .CLK(clk_i) );
  dff s_expa_in_reg_5_ ( .Q(s_expa_in_5_), .D(opa_i[28]), .CLK(clk_i) );
  dff s_expa_in_reg_4_ ( .Q(s_expa_in_4_), .D(opa_i[27]), .CLK(clk_i) );
  dff s_expa_in_reg_3_ ( .Q(s_expa_in_3_), .D(opa_i[26]), .CLK(clk_i) );
  dff s_expa_in_reg_2_ ( .Q(s_expa_in_2_), .D(opa_i[25]), .CLK(clk_i) );
  dff s_expa_in_reg_1_ ( .Q(s_expa_in_1_), .D(opa_i[24]), .CLK(clk_i) );
  dff s_expa_in_reg_0_ ( .Q(s_expa_in_0_), .D(n____return3431_0_), .CLK(clk_i)
         );
  dff s_expb_in_reg_8_ ( .Q(s_expb_in_8_), .D(1'b0), .CLK(clk_i) );
  dff s_expb_in_reg_7_ ( .Q(s_expb_in_7_), .D(opb_i[30]), .CLK(clk_i) );
  dff s_expb_in_reg_6_ ( .Q(s_expb_in_6_), .D(opb_i[29]), .CLK(clk_i) );
  dff s_expb_in_reg_5_ ( .Q(s_expb_in_5_), .D(opb_i[28]), .CLK(clk_i) );
  dff s_expb_in_reg_4_ ( .Q(s_expb_in_4_), .D(opb_i[27]), .CLK(clk_i) );
  dff s_expb_in_reg_3_ ( .Q(s_expb_in_3_), .D(opb_i[26]), .CLK(clk_i) );
  dff s_expb_in_reg_2_ ( .Q(s_expb_in_2_), .D(opb_i[25]), .CLK(clk_i) );
  dff s_expb_in_reg_1_ ( .Q(s_expb_in_1_), .D(opb_i[24]), .CLK(clk_i) );
  dff s_expb_in_reg_0_ ( .Q(s_expb_in_0_), .D(n____return3477_0_), .CLK(clk_i)
         );
  dff s_exp_10_o_reg_9_ ( .Q(s_exp_10_o[9]), .D(n____return3652_9_), .CLK(
        clk_i) );
  dff s_exp_10_o_reg_8_ ( .Q(s_exp_10_o[8]), .D(n3654_8_), .CLK(clk_i) );
  dff s_exp_10_o_reg_7_ ( .Q(s_exp_10_o[7]), .D(n____return3652_7_), .CLK(
        clk_i) );
  dff s_exp_10_o_reg_6_ ( .Q(s_exp_10_o[6]), .D(n____return3652_6_), .CLK(
        clk_i) );
  dff s_exp_10_o_reg_5_ ( .Q(s_exp_10_o[5]), .D(n____return3652_5_), .CLK(
        clk_i) );
  dff s_exp_10_o_reg_4_ ( .Q(s_exp_10_o[4]), .D(n____return3652_4_), .CLK(
        clk_i) );
  dff s_exp_10_o_reg_3_ ( .Q(s_exp_10_o[3]), .D(n____return3652_3_), .CLK(
        clk_i) );
  dff s_exp_10_o_reg_2_ ( .Q(s_exp_10_o[2]), .D(n____return3652_2_), .CLK(
        clk_i) );
  dff s_exp_10_o_reg_1_ ( .Q(s_exp_10_o[1]), .D(n____return3652_1_), .CLK(
        clk_i) );
  dff s_exp_10_o_reg_0_ ( .Q(s_exp_10_o[0]), .D(n____return3652_0_), .CLK(
        clk_i) );
  inv01 U1095 ( .Y(n4316), .A(n6455) );
  inv01 U1096 ( .Y(n4317), .A(n6453) );
  inv01 U1097 ( .Y(n4318), .A(n6451) );
  inv01 U1098 ( .Y(n4319), .A(n6449) );
  buf02 U1099 ( .Y(n4320), .A(n6269) );
  inv01 U1100 ( .Y(n6157), .A(n4321) );
  nor02 U1101 ( .Y(n4322), .A0(n6173), .A1(n4323) );
  nor02 U1102 ( .Y(n4324), .A0(n6173), .A1(n4325) );
  nor02 U1103 ( .Y(n4326), .A0(n6173), .A1(n4327) );
  nor02 U1104 ( .Y(n4328), .A0(n6173), .A1(n4329) );
  nor02 U1105 ( .Y(n4330), .A0(opb_i[2]), .A1(n4331) );
  nor02 U1106 ( .Y(n4332), .A0(opb_i[2]), .A1(n4333) );
  nor02 U1107 ( .Y(n4334), .A0(opb_i[2]), .A1(n4335) );
  nor02 U1108 ( .Y(n4336), .A0(opb_i[2]), .A1(n4337) );
  nor02 U1109 ( .Y(n4321), .A0(n4338), .A1(n4339) );
  nor02 U1110 ( .Y(n4340), .A0(n6140), .A1(n6141) );
  inv01 U1111 ( .Y(n4323), .A(n4340) );
  nor02 U1112 ( .Y(n4341), .A0(opb_i[0]), .A1(n6141) );
  inv01 U1113 ( .Y(n4325), .A(n4341) );
  nor02 U1114 ( .Y(n4342), .A0(n6140), .A1(opb_i[1]) );
  inv01 U1115 ( .Y(n4327), .A(n4342) );
  nor02 U1116 ( .Y(n4343), .A0(opb_i[0]), .A1(opb_i[1]) );
  inv01 U1117 ( .Y(n4329), .A(n4343) );
  nor02 U1118 ( .Y(n4344), .A0(n6140), .A1(n6141) );
  inv01 U1119 ( .Y(n4331), .A(n4344) );
  nor02 U1120 ( .Y(n4345), .A0(opb_i[0]), .A1(n6141) );
  inv01 U1121 ( .Y(n4333), .A(n4345) );
  nor02 U1122 ( .Y(n4346), .A0(n6140), .A1(opb_i[1]) );
  inv01 U1123 ( .Y(n4335), .A(n4346) );
  nor02 U1124 ( .Y(n4347), .A0(opb_i[0]), .A1(opb_i[1]) );
  inv01 U1125 ( .Y(n4337), .A(n4347) );
  nor02 U1126 ( .Y(n4348), .A0(n4322), .A1(n4324) );
  inv01 U1127 ( .Y(n4349), .A(n4348) );
  nor02 U1128 ( .Y(n4350), .A0(n4326), .A1(n4328) );
  inv01 U1129 ( .Y(n4351), .A(n4350) );
  nor02 U1130 ( .Y(n4352), .A0(n4349), .A1(n4351) );
  inv01 U1131 ( .Y(n4338), .A(n4352) );
  nor02 U1132 ( .Y(n4353), .A0(n4330), .A1(n4332) );
  inv01 U1133 ( .Y(n4354), .A(n4353) );
  nor02 U1134 ( .Y(n4355), .A0(n4334), .A1(n4336) );
  inv01 U1135 ( .Y(n4356), .A(n4355) );
  nor02 U1136 ( .Y(n4357), .A0(n4354), .A1(n4356) );
  inv01 U1137 ( .Y(n4339), .A(n4357) );
  buf08 U1138 ( .Y(n6140), .A(n6171) );
  buf08 U1139 ( .Y(n6141), .A(n6170) );
  inv04 U1140 ( .Y(n6173), .A(n6139) );
  nand02 U1141 ( .Y(n4358), .A0(opb_i[1]), .A1(n5161) );
  inv02 U1142 ( .Y(n4359), .A(n4358) );
  buf02 U1143 ( .Y(n4360), .A(opa_i[0]) );
  inv02 U1144 ( .Y(n4361), .A(n4360) );
  buf02 U1145 ( .Y(n4362), .A(n6440) );
  buf02 U1146 ( .Y(n4363), .A(opb_i[18]) );
  inv01 U1147 ( .Y(n4364), .A(n4363) );
  buf02 U1148 ( .Y(n4365), .A(opb_i[18]) );
  inv01 U1149 ( .Y(n4366), .A(n4365) );
  or02 U1150 ( .Y(n4367), .A0(n6367), .A1(n6122) );
  inv01 U1151 ( .Y(dvdnd_50_o[28]), .A(n4367) );
  or02 U1152 ( .Y(n4369), .A0(n5700), .A1(n6122) );
  inv01 U1153 ( .Y(dvdnd_50_o[26]), .A(n4369) );
  or02 U1154 ( .Y(n4371), .A0(n6369), .A1(n6120) );
  inv01 U1155 ( .Y(dvdnd_50_o[27]), .A(n4371) );
  ao22 U1156 ( .Y(n4373), .A0(n6298), .A1(n6304), .B0(n6086), .B1(n6332) );
  inv01 U1157 ( .Y(n4374), .A(n4373) );
  ao22 U1158 ( .Y(n4375), .A0(n6027), .A1(n6111), .B0(n6147), .B1(n6167) );
  inv01 U1159 ( .Y(n4376), .A(n4375) );
  ao22 U1160 ( .Y(n4377), .A0(n6156), .A1(n6111), .B0(n6166), .B1(n6167) );
  inv01 U1161 ( .Y(n4378), .A(n4377) );
  ao22 U1162 ( .Y(n4379), .A0(n6084), .A1(n6111), .B0(n6176), .B1(n6167) );
  inv01 U1163 ( .Y(n4380), .A(n4379) );
  or02 U1164 ( .Y(n4381), .A0(n6027), .A1(n6130) );
  inv01 U1165 ( .Y(dvsor_27_o[1]), .A(n4381) );
  ao22 U1166 ( .Y(n4383), .A0(n6088), .A1(n6198), .B0(n6159), .B1(n6165) );
  inv01 U1167 ( .Y(n4384), .A(n4383) );
  ao22 U1168 ( .Y(n4385), .A0(n6124), .A1(n6340), .B0(n6333), .B1(n6314) );
  inv01 U1169 ( .Y(n4386), .A(n4385) );
  ao22 U1170 ( .Y(n4387), .A0(n6124), .A1(n6346), .B0(n6333), .B1(n6320) );
  inv01 U1171 ( .Y(n4388), .A(n4387) );
  or02 U1172 ( .Y(n4389), .A0(n6156), .A1(n6130) );
  inv01 U1173 ( .Y(dvsor_27_o[3]), .A(n4389) );
  inv02 U1174 ( .Y(n4812), .A(opa_i[11]) );
  buf02 U1175 ( .Y(n4391), .A(s_div_zeros_2_) );
  or02 U1176 ( .Y(n4392), .A0(n6109), .A1(n6318) );
  inv01 U1177 ( .Y(dvdnd_50_o[31]), .A(n4392) );
  or02 U1178 ( .Y(n4394), .A0(n6128), .A1(n5163) );
  inv01 U1179 ( .Y(dvsor_27_o[0]), .A(n4394) );
  or02 U1180 ( .Y(n4396), .A0(n6084), .A1(n6128) );
  inv01 U1181 ( .Y(dvsor_27_o[2]), .A(n4396) );
  inv02 U1182 ( .Y(n4712), .A(opa_i[13]) );
  or02 U1183 ( .Y(n4398), .A0(n6357), .A1(n6120) );
  inv01 U1184 ( .Y(dvdnd_50_o[29]), .A(n4398) );
  buf02 U1185 ( .Y(n4400), .A(s_dvd_zeros_4_) );
  or02 U1186 ( .Y(n4401), .A0(n6118), .A1(n6154) );
  inv01 U1187 ( .Y(dvsor_27_o[6]), .A(n4401) );
  or02 U1188 ( .Y(n4403), .A0(n6118), .A1(n6153) );
  inv01 U1189 ( .Y(dvsor_27_o[7]), .A(n4403) );
  or02 U1190 ( .Y(n4405), .A0(n6118), .A1(n6155) );
  inv01 U1191 ( .Y(dvsor_27_o[5]), .A(n4405) );
  or02 U1192 ( .Y(n4407), .A0(n6110), .A1(n6312) );
  inv01 U1193 ( .Y(dvdnd_50_o[32]), .A(n4407) );
  buf02 U1194 ( .Y(n4409), .A(s_div_zeros_4_) );
  or02 U1195 ( .Y(n4410), .A0(n6305), .A1(n6109) );
  inv01 U1196 ( .Y(dvdnd_50_o[33]), .A(n4410) );
  ao22 U1197 ( .Y(n4412), .A0(n6123), .A1(n6211), .B0(n6088), .B1(n6183) );
  inv01 U1198 ( .Y(n4413), .A(n4412) );
  ao22 U1199 ( .Y(n4414), .A0(n6123), .A1(n6206), .B0(n6199), .B1(n6178) );
  inv01 U1200 ( .Y(n4415), .A(n4414) );
  nand02 U1201 ( .Y(n6376), .A0(n4416), .A1(n4417) );
  inv01 U1202 ( .Y(n4418), .A(n6354) );
  inv01 U1203 ( .Y(n4419), .A(n6089) );
  inv01 U1204 ( .Y(n4420), .A(n6367) );
  inv01 U1205 ( .Y(n4421), .A(n6360) );
  nand02 U1206 ( .Y(n4422), .A0(n4418), .A1(n4419) );
  nand02 U1207 ( .Y(n4423), .A0(n4418), .A1(n4420) );
  nand02 U1208 ( .Y(n4424), .A0(n4419), .A1(n4421) );
  nand02 U1209 ( .Y(n4425), .A0(n4420), .A1(n4421) );
  nand02 U1210 ( .Y(n4426), .A0(n4422), .A1(n4423) );
  inv01 U1211 ( .Y(n4416), .A(n4426) );
  nand02 U1212 ( .Y(n4427), .A0(n4424), .A1(n4425) );
  inv01 U1213 ( .Y(n4417), .A(n4427) );
  ao22 U1214 ( .Y(n4428), .A0(n6369), .A1(n6089), .B0(n6362), .B1(n6354) );
  inv01 U1215 ( .Y(n4429), .A(n4428) );
  ao22 U1216 ( .Y(n4430), .A0(n6357), .A1(n6089), .B0(n6365), .B1(n6354) );
  inv01 U1217 ( .Y(n4431), .A(n4430) );
  nor02 U1218 ( .Y(n4432), .A0(n5566), .A1(n6354) );
  inv02 U1219 ( .Y(n4433), .A(n4432) );
  nor02 U1220 ( .Y(n4434), .A0(n5678), .A1(n6167) );
  inv02 U1221 ( .Y(n4435), .A(n4434) );
  inv01 U1222 ( .Y(n6411), .A(n4436) );
  nand02 U1223 ( .Y(n4436), .A0(opa_i[9]), .A1(n4437) );
  nand02 U1224 ( .Y(n4438), .A0(n6430), .A1(n6070) );
  inv01 U1225 ( .Y(n4437), .A(n4438) );
  nand02 U1226 ( .Y(n4439), .A0(s_expa_in_7_), .A1(n6447) );
  inv02 U1227 ( .Y(n4908), .A(opa_i[22]) );
  inv02 U1228 ( .Y(n4801), .A(opa_i[6]) );
  buf02 U1229 ( .Y(dvsor_27_o[22]), .A(n6469) );
  inv02 U1230 ( .Y(n6030), .A(opa_i[19]) );
  inv02 U1231 ( .Y(n5077), .A(opa_i[19]) );
  buf02 U1232 ( .Y(dvdnd_50_o[48]), .A(n6466) );
  buf02 U1233 ( .Y(dvdnd_50_o[47]), .A(n6467) );
  buf02 U1234 ( .Y(dvsor_27_o[21]), .A(n6470) );
  buf02 U1235 ( .Y(dvdnd_50_o[46]), .A(n6468) );
  buf02 U1236 ( .Y(dvsor_27_o[20]), .A(n6471) );
  buf02 U1237 ( .Y(n4446), .A(opb_i[21]) );
  inv01 U1238 ( .Y(n4447), .A(n4446) );
  inv01 U1239 ( .Y(dvsor_27_o[23]), .A(n4448) );
  inv01 U1240 ( .Y(n4449), .A(n5506) );
  inv01 U1241 ( .Y(n4450), .A(n4735) );
  inv01 U1242 ( .Y(n4451), .A(n4447) );
  inv01 U1243 ( .Y(n4452), .A(n6158) );
  nor02 U1244 ( .Y(n4448), .A0(n4453), .A1(n4454) );
  nor02 U1245 ( .Y(n4455), .A0(n4449), .A1(n4450) );
  inv01 U1246 ( .Y(n4453), .A(n4455) );
  nor02 U1247 ( .Y(n4456), .A0(n4451), .A1(n4452) );
  inv01 U1248 ( .Y(n4454), .A(n4456) );
  inv02 U1249 ( .Y(n5014), .A(opa_i[21]) );
  inv01 U1250 ( .Y(dvdnd_50_o[49]), .A(n4457) );
  inv01 U1251 ( .Y(n4458), .A(n5504) );
  inv01 U1252 ( .Y(n4459), .A(n4737) );
  inv01 U1253 ( .Y(n4460), .A(n5014) );
  inv01 U1254 ( .Y(n4461), .A(n5086) );
  nor02 U1255 ( .Y(n4457), .A0(n4462), .A1(n4463) );
  nor02 U1256 ( .Y(n4464), .A0(n4458), .A1(n4459) );
  inv01 U1257 ( .Y(n4462), .A(n4464) );
  nor02 U1258 ( .Y(n4465), .A0(n4460), .A1(n4461) );
  inv01 U1259 ( .Y(n4463), .A(n4465) );
  nand02 U1260 ( .Y(n6222), .A0(n4466), .A1(n4467) );
  inv01 U1261 ( .Y(n4468), .A(opb_i[12]) );
  inv01 U1262 ( .Y(n4469), .A(opb_i[13]) );
  inv01 U1263 ( .Y(n4470), .A(n6141) );
  inv01 U1264 ( .Y(n4471), .A(n6140) );
  nand02 U1265 ( .Y(n4472), .A0(n4468), .A1(n4469) );
  nand02 U1266 ( .Y(n4473), .A0(n4468), .A1(n4470) );
  nand02 U1267 ( .Y(n4474), .A0(n4469), .A1(n4471) );
  nand02 U1268 ( .Y(n4475), .A0(n4470), .A1(n4471) );
  nand02 U1269 ( .Y(n4476), .A0(n4472), .A1(n4473) );
  inv01 U1270 ( .Y(n4466), .A(n4476) );
  nand02 U1271 ( .Y(n4477), .A0(n4474), .A1(n4475) );
  inv01 U1272 ( .Y(n4467), .A(n4477) );
  nand02 U1273 ( .Y(n6237), .A0(n4478), .A1(n4479) );
  inv01 U1274 ( .Y(n4480), .A(opb_i[8]) );
  inv01 U1275 ( .Y(n4481), .A(opb_i[9]) );
  inv01 U1276 ( .Y(n4482), .A(n6141) );
  inv01 U1277 ( .Y(n4483), .A(n6140) );
  nand02 U1278 ( .Y(n4484), .A0(n4480), .A1(n4481) );
  nand02 U1279 ( .Y(n4485), .A0(n4480), .A1(n4482) );
  nand02 U1280 ( .Y(n4486), .A0(n4481), .A1(n4483) );
  nand02 U1281 ( .Y(n4487), .A0(n4482), .A1(n4483) );
  nand02 U1282 ( .Y(n4488), .A0(n4484), .A1(n4485) );
  inv01 U1283 ( .Y(n4478), .A(n4488) );
  nand02 U1284 ( .Y(n4489), .A0(n4486), .A1(n4487) );
  inv01 U1285 ( .Y(n4479), .A(n4489) );
  inv02 U1286 ( .Y(n5928), .A(n5927) );
  nand02 U1287 ( .Y(n6225), .A0(n4490), .A1(n4491) );
  inv01 U1288 ( .Y(n4492), .A(opb_i[11]) );
  inv01 U1289 ( .Y(n4493), .A(opb_i[12]) );
  inv01 U1290 ( .Y(n4494), .A(n6141) );
  inv01 U1291 ( .Y(n4495), .A(n6140) );
  nand02 U1292 ( .Y(n4496), .A0(n4492), .A1(n4493) );
  nand02 U1293 ( .Y(n4497), .A0(n4492), .A1(n4494) );
  nand02 U1294 ( .Y(n4498), .A0(n4493), .A1(n4495) );
  nand02 U1295 ( .Y(n4499), .A0(n4494), .A1(n4495) );
  nand02 U1296 ( .Y(n4500), .A0(n4496), .A1(n4497) );
  inv01 U1297 ( .Y(n4490), .A(n4500) );
  nand02 U1298 ( .Y(n4501), .A0(n4498), .A1(n4499) );
  inv01 U1299 ( .Y(n4491), .A(n4501) );
  nand02 U1300 ( .Y(n6231), .A0(n4502), .A1(n4503) );
  inv01 U1301 ( .Y(n4504), .A(opb_i[10]) );
  inv01 U1302 ( .Y(n4505), .A(opb_i[11]) );
  inv01 U1303 ( .Y(n4506), .A(n6141) );
  inv01 U1304 ( .Y(n4507), .A(n6140) );
  nand02 U1305 ( .Y(n4508), .A0(n4504), .A1(n4505) );
  nand02 U1306 ( .Y(n4509), .A0(n4504), .A1(n4506) );
  nand02 U1307 ( .Y(n4510), .A0(n4505), .A1(n4507) );
  nand02 U1308 ( .Y(n4511), .A0(n4506), .A1(n4507) );
  nand02 U1309 ( .Y(n4512), .A0(n4508), .A1(n4509) );
  inv01 U1310 ( .Y(n4502), .A(n4512) );
  nand02 U1311 ( .Y(n4513), .A0(n4510), .A1(n4511) );
  inv01 U1312 ( .Y(n4503), .A(n4513) );
  nand02 U1313 ( .Y(n6230), .A0(n4514), .A1(n4515) );
  inv01 U1314 ( .Y(n4516), .A(opb_i[2]) );
  inv01 U1315 ( .Y(n4517), .A(opb_i[3]) );
  inv01 U1316 ( .Y(n4518), .A(n6141) );
  inv01 U1317 ( .Y(n4519), .A(n6140) );
  nand02 U1318 ( .Y(n4520), .A0(n4516), .A1(n4517) );
  nand02 U1319 ( .Y(n4521), .A0(n4516), .A1(n4518) );
  nand02 U1320 ( .Y(n4522), .A0(n4517), .A1(n4519) );
  nand02 U1321 ( .Y(n4523), .A0(n4518), .A1(n4519) );
  nand02 U1322 ( .Y(n4524), .A0(n4520), .A1(n4521) );
  inv01 U1323 ( .Y(n4514), .A(n4524) );
  nand02 U1324 ( .Y(n4525), .A0(n4522), .A1(n4523) );
  inv01 U1325 ( .Y(n4515), .A(n4525) );
  nand02 U1326 ( .Y(n6236), .A0(n4526), .A1(n4527) );
  inv01 U1327 ( .Y(n4528), .A(opb_i[4]) );
  inv01 U1328 ( .Y(n4529), .A(opb_i[5]) );
  inv01 U1329 ( .Y(n4530), .A(n6141) );
  inv01 U1330 ( .Y(n4531), .A(n6140) );
  nand02 U1331 ( .Y(n4532), .A0(n4528), .A1(n4529) );
  nand02 U1332 ( .Y(n4533), .A0(n4528), .A1(n4530) );
  nand02 U1333 ( .Y(n4534), .A0(n4529), .A1(n4531) );
  nand02 U1334 ( .Y(n4535), .A0(n4530), .A1(n4531) );
  nand02 U1335 ( .Y(n4536), .A0(n4532), .A1(n4533) );
  inv01 U1336 ( .Y(n4526), .A(n4536) );
  nand02 U1337 ( .Y(n4537), .A0(n4534), .A1(n4535) );
  inv01 U1338 ( .Y(n4527), .A(n4537) );
  nand02 U1339 ( .Y(n6227), .A0(n4538), .A1(n4539) );
  inv01 U1340 ( .Y(n4540), .A(opb_i[7]) );
  inv01 U1341 ( .Y(n4541), .A(opb_i[8]) );
  inv01 U1342 ( .Y(n4542), .A(n6141) );
  inv01 U1343 ( .Y(n4543), .A(n6140) );
  nand02 U1344 ( .Y(n4544), .A0(n4540), .A1(n4541) );
  nand02 U1345 ( .Y(n4545), .A0(n4540), .A1(n4542) );
  nand02 U1346 ( .Y(n4546), .A0(n4541), .A1(n4543) );
  nand02 U1347 ( .Y(n4547), .A0(n4542), .A1(n4543) );
  nand02 U1348 ( .Y(n4548), .A0(n4544), .A1(n4545) );
  inv01 U1349 ( .Y(n4538), .A(n4548) );
  nand02 U1350 ( .Y(n4549), .A0(n4546), .A1(n4547) );
  inv01 U1351 ( .Y(n4539), .A(n4549) );
  nand02 U1352 ( .Y(n6224), .A0(n4550), .A1(n4551) );
  inv01 U1353 ( .Y(n4552), .A(opb_i[3]) );
  inv01 U1354 ( .Y(n4553), .A(opb_i[4]) );
  inv01 U1355 ( .Y(n4554), .A(n6141) );
  inv01 U1356 ( .Y(n4555), .A(n6140) );
  nand02 U1357 ( .Y(n4556), .A0(n4552), .A1(n4553) );
  nand02 U1358 ( .Y(n4557), .A0(n4552), .A1(n4554) );
  nand02 U1359 ( .Y(n4558), .A0(n4553), .A1(n4555) );
  nand02 U1360 ( .Y(n4559), .A0(n4554), .A1(n4555) );
  nand02 U1361 ( .Y(n4560), .A0(n4556), .A1(n4557) );
  inv01 U1362 ( .Y(n4550), .A(n4560) );
  nand02 U1363 ( .Y(n4561), .A0(n4558), .A1(n4559) );
  inv01 U1364 ( .Y(n4551), .A(n4561) );
  nand02 U1365 ( .Y(n6228), .A0(n4562), .A1(n4563) );
  inv01 U1366 ( .Y(n4564), .A(opb_i[6]) );
  inv01 U1367 ( .Y(n4565), .A(opb_i[7]) );
  inv01 U1368 ( .Y(n4566), .A(n6141) );
  inv01 U1369 ( .Y(n4567), .A(n6140) );
  nand02 U1370 ( .Y(n4568), .A0(n4564), .A1(n4565) );
  nand02 U1371 ( .Y(n4569), .A0(n4564), .A1(n4566) );
  nand02 U1372 ( .Y(n4570), .A0(n4565), .A1(n4567) );
  nand02 U1373 ( .Y(n4571), .A0(n4566), .A1(n4567) );
  nand02 U1374 ( .Y(n4572), .A0(n4568), .A1(n4569) );
  inv01 U1375 ( .Y(n4562), .A(n4572) );
  nand02 U1376 ( .Y(n4573), .A0(n4570), .A1(n4571) );
  inv01 U1377 ( .Y(n4563), .A(n4573) );
  nand02 U1378 ( .Y(n6234), .A0(n4574), .A1(n4575) );
  inv01 U1379 ( .Y(n4576), .A(opb_i[1]) );
  inv01 U1380 ( .Y(n4577), .A(opb_i[2]) );
  inv01 U1381 ( .Y(n4578), .A(n6141) );
  inv01 U1382 ( .Y(n4579), .A(n6140) );
  nand02 U1383 ( .Y(n4580), .A0(n4576), .A1(n4577) );
  nand02 U1384 ( .Y(n4581), .A0(n4576), .A1(n4578) );
  nand02 U1385 ( .Y(n4582), .A0(n4577), .A1(n4579) );
  nand02 U1386 ( .Y(n4583), .A0(n4578), .A1(n4579) );
  nand02 U1387 ( .Y(n4584), .A0(n4580), .A1(n4581) );
  inv01 U1388 ( .Y(n4574), .A(n4584) );
  nand02 U1389 ( .Y(n4585), .A0(n4582), .A1(n4583) );
  inv01 U1390 ( .Y(n4575), .A(n4585) );
  nand02 U1391 ( .Y(n6232), .A0(n4586), .A1(n4587) );
  inv01 U1392 ( .Y(n4588), .A(opb_i[9]) );
  inv01 U1393 ( .Y(n4589), .A(opb_i[10]) );
  inv01 U1394 ( .Y(n4590), .A(n6141) );
  inv01 U1395 ( .Y(n4591), .A(n6140) );
  nand02 U1396 ( .Y(n4592), .A0(n4588), .A1(n4589) );
  nand02 U1397 ( .Y(n4593), .A0(n4588), .A1(n4590) );
  nand02 U1398 ( .Y(n4594), .A0(n4589), .A1(n4591) );
  nand02 U1399 ( .Y(n4595), .A0(n4590), .A1(n4591) );
  nand02 U1400 ( .Y(n4596), .A0(n4592), .A1(n4593) );
  inv01 U1401 ( .Y(n4586), .A(n4596) );
  nand02 U1402 ( .Y(n4597), .A0(n4594), .A1(n4595) );
  inv01 U1403 ( .Y(n4587), .A(n4597) );
  inv04 U1404 ( .Y(n6158), .A(opb_i[20]) );
  nand02 U1405 ( .Y(n6235), .A0(n4598), .A1(n4599) );
  inv01 U1406 ( .Y(n4600), .A(opb_i[5]) );
  inv01 U1407 ( .Y(n4601), .A(opb_i[6]) );
  inv01 U1408 ( .Y(n4602), .A(n6141) );
  inv01 U1409 ( .Y(n4603), .A(n6140) );
  nand02 U1410 ( .Y(n4604), .A0(n4600), .A1(n4601) );
  nand02 U1411 ( .Y(n4605), .A0(n4600), .A1(n4602) );
  nand02 U1412 ( .Y(n4606), .A0(n4601), .A1(n4603) );
  nand02 U1413 ( .Y(n4607), .A0(n4602), .A1(n4603) );
  nand02 U1414 ( .Y(n4608), .A0(n4604), .A1(n4605) );
  inv01 U1415 ( .Y(n4598), .A(n4608) );
  nand02 U1416 ( .Y(n4609), .A0(n4606), .A1(n4607) );
  inv01 U1417 ( .Y(n4599), .A(n4609) );
  nand02 U1418 ( .Y(n6208), .A0(n4610), .A1(n4611) );
  inv01 U1419 ( .Y(n4612), .A(opb_i[16]) );
  inv01 U1420 ( .Y(n4613), .A(opb_i[17]) );
  inv01 U1421 ( .Y(n4614), .A(n6141) );
  inv01 U1422 ( .Y(n4615), .A(n6140) );
  nand02 U1423 ( .Y(n4616), .A0(n4612), .A1(n4613) );
  nand02 U1424 ( .Y(n4617), .A0(n4612), .A1(n4614) );
  nand02 U1425 ( .Y(n4618), .A0(n4613), .A1(n4615) );
  nand02 U1426 ( .Y(n4619), .A0(n4614), .A1(n4615) );
  nand02 U1427 ( .Y(n4620), .A0(n4616), .A1(n4617) );
  inv01 U1428 ( .Y(n4610), .A(n4620) );
  nand02 U1429 ( .Y(n4621), .A0(n4618), .A1(n4619) );
  inv01 U1430 ( .Y(n4611), .A(n4621) );
  or03 U1431 ( .Y(n4622), .A0(n6261), .A1(n6254), .A2(n6262) );
  inv01 U1432 ( .Y(n4623), .A(n4622) );
  or03 U1433 ( .Y(n4624), .A0(n6257), .A1(n6260), .A2(n6258) );
  inv01 U1434 ( .Y(n4625), .A(n4624) );
  nand02 U1435 ( .Y(n6214), .A0(n4626), .A1(n4627) );
  inv01 U1436 ( .Y(n4628), .A(opb_i[15]) );
  inv01 U1437 ( .Y(n4629), .A(opb_i[16]) );
  inv01 U1438 ( .Y(n4630), .A(n6141) );
  inv01 U1439 ( .Y(n4631), .A(n6140) );
  nand02 U1440 ( .Y(n4632), .A0(n4628), .A1(n4629) );
  nand02 U1441 ( .Y(n4633), .A0(n4628), .A1(n4630) );
  nand02 U1442 ( .Y(n4634), .A0(n4629), .A1(n4631) );
  nand02 U1443 ( .Y(n4635), .A0(n4630), .A1(n4631) );
  nand02 U1444 ( .Y(n4636), .A0(n4632), .A1(n4633) );
  inv01 U1445 ( .Y(n4626), .A(n4636) );
  nand02 U1446 ( .Y(n4637), .A0(n4634), .A1(n4635) );
  inv01 U1447 ( .Y(n4627), .A(n4637) );
  nand02 U1448 ( .Y(n6219), .A0(n4638), .A1(n4639) );
  inv01 U1449 ( .Y(n4640), .A(opb_i[14]) );
  inv01 U1450 ( .Y(n4641), .A(opb_i[15]) );
  inv01 U1451 ( .Y(n4642), .A(n6141) );
  inv01 U1452 ( .Y(n4643), .A(n6140) );
  nand02 U1453 ( .Y(n4644), .A0(n4640), .A1(n4641) );
  nand02 U1454 ( .Y(n4645), .A0(n4640), .A1(n4642) );
  nand02 U1455 ( .Y(n4646), .A0(n4641), .A1(n4643) );
  nand02 U1456 ( .Y(n4647), .A0(n4642), .A1(n4643) );
  nand02 U1457 ( .Y(n4648), .A0(n4644), .A1(n4645) );
  inv01 U1458 ( .Y(n4638), .A(n4648) );
  nand02 U1459 ( .Y(n4649), .A0(n4646), .A1(n4647) );
  inv01 U1460 ( .Y(n4639), .A(n4649) );
  nand02 U1461 ( .Y(n6221), .A0(n4650), .A1(n4651) );
  inv01 U1462 ( .Y(n4652), .A(opb_i[13]) );
  inv01 U1463 ( .Y(n4653), .A(opb_i[14]) );
  inv01 U1464 ( .Y(n4654), .A(n6141) );
  inv01 U1465 ( .Y(n4655), .A(n6140) );
  nand02 U1466 ( .Y(n4656), .A0(n4652), .A1(n4653) );
  nand02 U1467 ( .Y(n4657), .A0(n4652), .A1(n4654) );
  nand02 U1468 ( .Y(n4658), .A0(n4653), .A1(n4655) );
  nand02 U1469 ( .Y(n4659), .A0(n4654), .A1(n4655) );
  nand02 U1470 ( .Y(n4660), .A0(n4656), .A1(n4657) );
  inv01 U1471 ( .Y(n4650), .A(n4660) );
  nand02 U1472 ( .Y(n4661), .A0(n4658), .A1(n4659) );
  inv01 U1473 ( .Y(n4651), .A(n4661) );
  nand02 U1474 ( .Y(n6202), .A0(n4662), .A1(n4663) );
  inv01 U1475 ( .Y(n4664), .A(opb_i[17]) );
  inv01 U1476 ( .Y(n4665), .A(opb_i[18]) );
  inv01 U1477 ( .Y(n4666), .A(n6141) );
  inv01 U1478 ( .Y(n4667), .A(n6140) );
  nand02 U1479 ( .Y(n4668), .A0(n4664), .A1(n4665) );
  nand02 U1480 ( .Y(n4669), .A0(n4664), .A1(n4666) );
  nand02 U1481 ( .Y(n4670), .A0(n4665), .A1(n4667) );
  nand02 U1482 ( .Y(n4671), .A0(n4666), .A1(n4667) );
  nand02 U1483 ( .Y(n4672), .A0(n4668), .A1(n4669) );
  inv01 U1484 ( .Y(n4662), .A(n4672) );
  nand02 U1485 ( .Y(n4673), .A0(n4670), .A1(n4671) );
  inv01 U1486 ( .Y(n4663), .A(n4673) );
  inv02 U1487 ( .Y(n6149), .A(n6152) );
  or03 U1488 ( .Y(n4674), .A0(n6391), .A1(n6392), .A2(n6384) );
  inv01 U1489 ( .Y(n4675), .A(n4674) );
  or03 U1490 ( .Y(n4676), .A0(n5680), .A1(n6389), .A2(n6388) );
  inv01 U1491 ( .Y(n4677), .A(n4676) );
  inv01 U1492 ( .Y(n6438), .A(n4678) );
  inv01 U1493 ( .Y(n4679), .A(n6386) );
  inv01 U1494 ( .Y(n4680), .A(n6387) );
  inv01 U1495 ( .Y(n4681), .A(n6385) );
  nand02 U1496 ( .Y(n4678), .A0(n4681), .A1(n4682) );
  nand02 U1497 ( .Y(n4683), .A0(n4679), .A1(n4680) );
  inv01 U1498 ( .Y(n4682), .A(n4683) );
  nand03 U1499 ( .Y(n4684), .A0(n5155), .A1(n6049), .A2(n6293) );
  inv02 U1500 ( .Y(n4685), .A(n4684) );
  nand03 U1501 ( .Y(n4686), .A0(n5157), .A1(n6055), .A2(n6295) );
  inv02 U1502 ( .Y(n4687), .A(n4686) );
  or03 U1503 ( .Y(n4688), .A0(n6395), .A1(n6393), .A2(n6394) );
  inv01 U1504 ( .Y(n4689), .A(n4688) );
  ao22 U1505 ( .Y(n4690), .A0(n6298), .A1(n6325), .B0(n6086), .B1(n6326) );
  inv01 U1506 ( .Y(n4691), .A(n4690) );
  ao22 U1507 ( .Y(n4692), .A0(n6159), .A1(n6184), .B0(n6088), .B1(n6185) );
  inv01 U1508 ( .Y(n4693), .A(n4692) );
  ao22 U1509 ( .Y(n4694), .A0(n6298), .A1(n6319), .B0(n6086), .B1(n6320) );
  inv01 U1510 ( .Y(n4695), .A(n4694) );
  ao22 U1511 ( .Y(n4696), .A0(n6298), .A1(n6313), .B0(n6086), .B1(n6314) );
  inv01 U1512 ( .Y(n4697), .A(n4696) );
  ao22 U1513 ( .Y(n4698), .A0(n6159), .A1(n6191), .B0(n6088), .B1(n6192) );
  inv01 U1514 ( .Y(n4699), .A(n4698) );
  ao22 U1515 ( .Y(n4700), .A0(n6159), .A1(n6177), .B0(n6088), .B1(n6178) );
  inv01 U1516 ( .Y(n4701), .A(n4700) );
  nand02 U1517 ( .Y(n6270), .A0(n4702), .A1(n4703) );
  inv01 U1518 ( .Y(n4704), .A(opb_i[22]) );
  inv01 U1519 ( .Y(n4705), .A(n4447) );
  nand02 U1520 ( .Y(n4702), .A0(n4704), .A1(n4705) );
  nand02 U1521 ( .Y(n4703), .A0(n4704), .A1(n6158) );
  ao22 U1522 ( .Y(n4706), .A0(n6163), .A1(n6181), .B0(n6123), .B1(n6182) );
  inv01 U1523 ( .Y(n4707), .A(n4706) );
  ao22 U1524 ( .Y(n4708), .A0(n6163), .A1(n6174), .B0(n6123), .B1(n6175) );
  inv01 U1525 ( .Y(n4709), .A(n4708) );
  nand02 U1526 ( .Y(n6359), .A0(n4710), .A1(n4711) );
  inv01 U1527 ( .Y(n4713), .A(opa_i[12]) );
  inv01 U1528 ( .Y(n4714), .A(n6137) );
  inv01 U1529 ( .Y(n4715), .A(n6309) );
  nand02 U1530 ( .Y(n4716), .A0(n4712), .A1(n4713) );
  nand02 U1531 ( .Y(n4717), .A0(n4712), .A1(n4714) );
  nand02 U1532 ( .Y(n4718), .A0(n4713), .A1(n4715) );
  nand02 U1533 ( .Y(n4719), .A0(n4714), .A1(n4715) );
  nand02 U1534 ( .Y(n4720), .A0(n4716), .A1(n4717) );
  inv01 U1535 ( .Y(n4710), .A(n4720) );
  nand02 U1536 ( .Y(n4721), .A0(n4718), .A1(n4719) );
  inv01 U1537 ( .Y(n4711), .A(n4721) );
  nand02 U1538 ( .Y(n6368), .A0(n4722), .A1(n4723) );
  inv01 U1539 ( .Y(n4724), .A(opa_i[8]) );
  inv01 U1540 ( .Y(n4725), .A(opa_i[7]) );
  inv01 U1541 ( .Y(n4726), .A(n6137) );
  inv01 U1542 ( .Y(n4727), .A(n6309) );
  nand02 U1543 ( .Y(n4728), .A0(n4724), .A1(n4725) );
  nand02 U1544 ( .Y(n4729), .A0(n4724), .A1(n4726) );
  nand02 U1545 ( .Y(n4730), .A0(n4725), .A1(n4727) );
  nand02 U1546 ( .Y(n4731), .A0(n4726), .A1(n4727) );
  nand02 U1547 ( .Y(n4732), .A0(n4728), .A1(n4729) );
  inv01 U1548 ( .Y(n4722), .A(n4732) );
  nand02 U1549 ( .Y(n4733), .A0(n4730), .A1(n4731) );
  inv01 U1550 ( .Y(n4723), .A(n4733) );
  ao22 U1551 ( .Y(n4734), .A0(n6163), .A1(n6164), .B0(n6123), .B1(n6165) );
  inv01 U1552 ( .Y(n4735), .A(n4734) );
  ao22 U1553 ( .Y(n4736), .A0(n6302), .A1(n6303), .B0(n6124), .B1(n6304) );
  inv01 U1554 ( .Y(n4737), .A(n4736) );
  ao22 U1555 ( .Y(n4738), .A0(n6316), .A1(n6302), .B0(n6124), .B1(n6317) );
  inv01 U1556 ( .Y(n4739), .A(n4738) );
  ao22 U1557 ( .Y(n4740), .A0(n6310), .A1(n6302), .B0(n6124), .B1(n6311) );
  inv01 U1558 ( .Y(n4741), .A(n4740) );
  nand02 U1559 ( .Y(n6379), .A0(n4742), .A1(n4743) );
  inv01 U1560 ( .Y(n4744), .A(opa_i[2]) );
  inv01 U1561 ( .Y(n4745), .A(n6137) );
  inv01 U1562 ( .Y(n4746), .A(n6309) );
  nand02 U1563 ( .Y(n4747), .A0(n4744), .A1(n6044) );
  nand02 U1564 ( .Y(n4748), .A0(n4744), .A1(n4745) );
  nand02 U1565 ( .Y(n4749), .A0(n6044), .A1(n4746) );
  nand02 U1566 ( .Y(n4750), .A0(n4745), .A1(n4746) );
  nand02 U1567 ( .Y(n4751), .A0(n4747), .A1(n4748) );
  inv01 U1568 ( .Y(n4742), .A(n4751) );
  nand02 U1569 ( .Y(n4752), .A0(n4749), .A1(n4750) );
  inv01 U1570 ( .Y(n4743), .A(n4752) );
  nand02 U1571 ( .Y(n6361), .A0(n4753), .A1(n4754) );
  inv01 U1572 ( .Y(n4755), .A(opa_i[12]) );
  inv01 U1573 ( .Y(n4756), .A(n6137) );
  inv01 U1574 ( .Y(n4757), .A(n6309) );
  nand02 U1575 ( .Y(n4758), .A0(n4755), .A1(n4812) );
  nand02 U1576 ( .Y(n4759), .A0(n4755), .A1(n4756) );
  nand02 U1577 ( .Y(n4760), .A0(n4812), .A1(n4757) );
  nand02 U1578 ( .Y(n4761), .A0(n4756), .A1(n4757) );
  nand02 U1579 ( .Y(n4762), .A0(n4758), .A1(n4759) );
  inv01 U1580 ( .Y(n4753), .A(n4762) );
  nand02 U1581 ( .Y(n4763), .A0(n4760), .A1(n4761) );
  inv01 U1582 ( .Y(n4754), .A(n4763) );
  nand02 U1583 ( .Y(n6375), .A0(n4764), .A1(n4765) );
  inv01 U1584 ( .Y(n4766), .A(opa_i[5]) );
  inv01 U1585 ( .Y(n4767), .A(n6137) );
  inv01 U1586 ( .Y(n4768), .A(n6309) );
  nand02 U1587 ( .Y(n4769), .A0(n4766), .A1(n5682) );
  nand02 U1588 ( .Y(n4770), .A0(n4766), .A1(n4767) );
  nand02 U1589 ( .Y(n4771), .A0(n5682), .A1(n4768) );
  nand02 U1590 ( .Y(n4772), .A0(n4767), .A1(n4768) );
  nand02 U1591 ( .Y(n4773), .A0(n4769), .A1(n4770) );
  inv01 U1592 ( .Y(n4764), .A(n4773) );
  nand02 U1593 ( .Y(n4774), .A0(n4771), .A1(n4772) );
  inv01 U1594 ( .Y(n4765), .A(n4774) );
  nand02 U1595 ( .Y(n6378), .A0(n4775), .A1(n4776) );
  inv01 U1596 ( .Y(n4777), .A(opa_i[3]) );
  inv01 U1597 ( .Y(n4778), .A(opa_i[2]) );
  inv01 U1598 ( .Y(n4779), .A(n6137) );
  inv01 U1599 ( .Y(n4780), .A(n6309) );
  nand02 U1600 ( .Y(n4781), .A0(n4777), .A1(n4778) );
  nand02 U1601 ( .Y(n4782), .A0(n4777), .A1(n4779) );
  nand02 U1602 ( .Y(n4783), .A0(n4778), .A1(n4780) );
  nand02 U1603 ( .Y(n4784), .A0(n4779), .A1(n4780) );
  nand02 U1604 ( .Y(n4785), .A0(n4781), .A1(n4782) );
  inv01 U1605 ( .Y(n4775), .A(n4785) );
  nand02 U1606 ( .Y(n4786), .A0(n4783), .A1(n4784) );
  inv01 U1607 ( .Y(n4776), .A(n4786) );
  nand02 U1608 ( .Y(n6364), .A0(n4787), .A1(n4788) );
  inv01 U1609 ( .Y(n4789), .A(opa_i[10]) );
  inv01 U1610 ( .Y(n4790), .A(opa_i[9]) );
  inv01 U1611 ( .Y(n4791), .A(n6137) );
  inv01 U1612 ( .Y(n4792), .A(n6309) );
  nand02 U1613 ( .Y(n4793), .A0(n4789), .A1(n4790) );
  nand02 U1614 ( .Y(n4794), .A0(n4789), .A1(n4791) );
  nand02 U1615 ( .Y(n4795), .A0(n4790), .A1(n4792) );
  nand02 U1616 ( .Y(n4796), .A0(n4791), .A1(n4792) );
  nand02 U1617 ( .Y(n4797), .A0(n4793), .A1(n4794) );
  inv01 U1618 ( .Y(n4787), .A(n4797) );
  nand02 U1619 ( .Y(n4798), .A0(n4795), .A1(n4796) );
  inv01 U1620 ( .Y(n4788), .A(n4798) );
  nand02 U1621 ( .Y(n6374), .A0(n4799), .A1(n4800) );
  inv01 U1622 ( .Y(n4802), .A(n6137) );
  inv01 U1623 ( .Y(n4803), .A(n6309) );
  nand02 U1624 ( .Y(n4804), .A0(n4801), .A1(n6076) );
  nand02 U1625 ( .Y(n4805), .A0(n4801), .A1(n4802) );
  nand02 U1626 ( .Y(n4806), .A0(n6076), .A1(n4803) );
  nand02 U1627 ( .Y(n4807), .A0(n4802), .A1(n4803) );
  nand02 U1628 ( .Y(n4808), .A0(n4804), .A1(n4805) );
  inv01 U1629 ( .Y(n4799), .A(n4808) );
  nand02 U1630 ( .Y(n4809), .A0(n4806), .A1(n4807) );
  inv01 U1631 ( .Y(n4800), .A(n4809) );
  nand02 U1632 ( .Y(n6363), .A0(n4810), .A1(n4811) );
  inv01 U1633 ( .Y(n4813), .A(n6137) );
  inv01 U1634 ( .Y(n4814), .A(n6309) );
  nand02 U1635 ( .Y(n4815), .A0(n4812), .A1(n6070) );
  nand02 U1636 ( .Y(n4816), .A0(n4812), .A1(n4813) );
  nand02 U1637 ( .Y(n4817), .A0(n6070), .A1(n4814) );
  nand02 U1638 ( .Y(n4818), .A0(n4813), .A1(n4814) );
  nand02 U1639 ( .Y(n4819), .A0(n4815), .A1(n4816) );
  inv01 U1640 ( .Y(n4810), .A(n4819) );
  nand02 U1641 ( .Y(n4820), .A0(n4817), .A1(n4818) );
  inv01 U1642 ( .Y(n4811), .A(n4820) );
  nand02 U1643 ( .Y(n6377), .A0(n4821), .A1(n4822) );
  inv01 U1644 ( .Y(n4823), .A(opa_i[4]) );
  inv01 U1645 ( .Y(n4824), .A(n6137) );
  inv01 U1646 ( .Y(n4825), .A(n6309) );
  nand02 U1647 ( .Y(n4826), .A0(n4823), .A1(n6078) );
  nand02 U1648 ( .Y(n4827), .A0(n4823), .A1(n4824) );
  nand02 U1649 ( .Y(n4828), .A0(n6078), .A1(n4825) );
  nand02 U1650 ( .Y(n4829), .A0(n4824), .A1(n4825) );
  nand02 U1651 ( .Y(n4830), .A0(n4826), .A1(n4827) );
  inv01 U1652 ( .Y(n4821), .A(n4830) );
  nand02 U1653 ( .Y(n4831), .A0(n4828), .A1(n4829) );
  inv01 U1654 ( .Y(n4822), .A(n4831) );
  nand02 U1655 ( .Y(n6356), .A0(n4832), .A1(n4833) );
  inv01 U1656 ( .Y(n4834), .A(opa_i[14]) );
  inv01 U1657 ( .Y(n4835), .A(n6137) );
  inv01 U1658 ( .Y(n4836), .A(n6309) );
  nand02 U1659 ( .Y(n4837), .A0(n4834), .A1(n4712) );
  nand02 U1660 ( .Y(n4838), .A0(n4834), .A1(n4835) );
  nand02 U1661 ( .Y(n4839), .A0(n4712), .A1(n4836) );
  nand02 U1662 ( .Y(n4840), .A0(n4835), .A1(n4836) );
  nand02 U1663 ( .Y(n4841), .A0(n4837), .A1(n4838) );
  inv01 U1664 ( .Y(n4832), .A(n4841) );
  nand02 U1665 ( .Y(n4842), .A0(n4839), .A1(n4840) );
  inv01 U1666 ( .Y(n4833), .A(n4842) );
  nand02 U1667 ( .Y(n6366), .A0(n4843), .A1(n4844) );
  inv01 U1668 ( .Y(n4845), .A(opa_i[9]) );
  inv01 U1669 ( .Y(n4846), .A(n6137) );
  inv01 U1670 ( .Y(n4847), .A(n6309) );
  nand02 U1671 ( .Y(n4848), .A0(n4845), .A1(n6370) );
  nand02 U1672 ( .Y(n4849), .A0(n4845), .A1(n4846) );
  nand02 U1673 ( .Y(n4850), .A0(n6370), .A1(n4847) );
  nand02 U1674 ( .Y(n4851), .A0(n4846), .A1(n4847) );
  nand02 U1675 ( .Y(n4852), .A0(n4848), .A1(n4849) );
  inv01 U1676 ( .Y(n4843), .A(n4852) );
  nand02 U1677 ( .Y(n4853), .A0(n4850), .A1(n4851) );
  inv01 U1678 ( .Y(n4844), .A(n4853) );
  or02 U1679 ( .Y(n4854), .A0(n4439), .A1(n6446) );
  inv01 U1680 ( .Y(n4855), .A(n4854) );
  inv02 U1681 ( .Y(n6392), .A(n4856) );
  nand02 U1682 ( .Y(n4856), .A0(opa_i[16]), .A1(n4857) );
  nand02 U1683 ( .Y(n4858), .A0(n6441), .A1(n6005) );
  inv01 U1684 ( .Y(n4857), .A(n4858) );
  nand02 U1685 ( .Y(n6380), .A0(n4859), .A1(n4860) );
  inv01 U1686 ( .Y(n4861), .A(opa_i[1]) );
  inv01 U1687 ( .Y(n4862), .A(n6137) );
  inv01 U1688 ( .Y(n4863), .A(n6309) );
  nand02 U1689 ( .Y(n4864), .A0(n4861), .A1(n4361) );
  nand02 U1690 ( .Y(n4865), .A0(n4861), .A1(n4862) );
  nand02 U1691 ( .Y(n4866), .A0(n4361), .A1(n4863) );
  nand02 U1692 ( .Y(n4867), .A0(n4862), .A1(n4863) );
  nand02 U1693 ( .Y(n4868), .A0(n4864), .A1(n4865) );
  inv01 U1694 ( .Y(n4859), .A(n4868) );
  nand02 U1695 ( .Y(n4869), .A0(n4866), .A1(n4867) );
  inv01 U1696 ( .Y(n4860), .A(n4869) );
  nand02 U1697 ( .Y(n6348), .A0(n4870), .A1(n4871) );
  inv01 U1698 ( .Y(n4872), .A(opa_i[15]) );
  inv01 U1699 ( .Y(n4873), .A(n6137) );
  inv01 U1700 ( .Y(n4874), .A(n6309) );
  nand02 U1701 ( .Y(n4875), .A0(n4872), .A1(n6080) );
  nand02 U1702 ( .Y(n4876), .A0(n4872), .A1(n4873) );
  nand02 U1703 ( .Y(n4877), .A0(n6080), .A1(n4874) );
  nand02 U1704 ( .Y(n4878), .A0(n4873), .A1(n4874) );
  nand02 U1705 ( .Y(n4879), .A0(n4875), .A1(n4876) );
  inv01 U1706 ( .Y(n4870), .A(n4879) );
  nand02 U1707 ( .Y(n4880), .A0(n4877), .A1(n4878) );
  inv01 U1708 ( .Y(n4871), .A(n4880) );
  inv02 U1709 ( .Y(n6389), .A(n4881) );
  nand02 U1710 ( .Y(n4881), .A0(opa_i[2]), .A1(n4882) );
  nand02 U1711 ( .Y(n4883), .A0(n6437), .A1(n6078) );
  inv01 U1712 ( .Y(n4882), .A(n4883) );
  nand02 U1713 ( .Y(n6371), .A0(n4884), .A1(n4885) );
  inv01 U1714 ( .Y(n4886), .A(opa_i[7]) );
  inv01 U1715 ( .Y(n4887), .A(n6137) );
  inv01 U1716 ( .Y(n4888), .A(n6309) );
  nand02 U1717 ( .Y(n4889), .A0(n4886), .A1(n4801) );
  nand02 U1718 ( .Y(n4890), .A0(n4886), .A1(n4887) );
  nand02 U1719 ( .Y(n4891), .A0(n4801), .A1(n4888) );
  nand02 U1720 ( .Y(n4892), .A0(n4887), .A1(n4888) );
  nand02 U1721 ( .Y(n4893), .A0(n4889), .A1(n4890) );
  inv01 U1722 ( .Y(n4884), .A(n4893) );
  nand02 U1723 ( .Y(n4894), .A0(n4891), .A1(n4892) );
  inv01 U1724 ( .Y(n4885), .A(n4894) );
  nand02 U1725 ( .Y(n6336), .A0(n4895), .A1(n4896) );
  inv01 U1726 ( .Y(n4897), .A(opa_i[17]) );
  inv01 U1727 ( .Y(n4898), .A(n6137) );
  inv01 U1728 ( .Y(n4899), .A(n6309) );
  nand02 U1729 ( .Y(n4900), .A0(n4897), .A1(n5991) );
  nand02 U1730 ( .Y(n4901), .A0(n4897), .A1(n4898) );
  nand02 U1731 ( .Y(n4902), .A0(n5991), .A1(n4899) );
  nand02 U1732 ( .Y(n4903), .A0(n4898), .A1(n4899) );
  nand02 U1733 ( .Y(n4904), .A0(n4900), .A1(n4901) );
  inv01 U1734 ( .Y(n4895), .A(n4904) );
  nand02 U1735 ( .Y(n4905), .A0(n4902), .A1(n4903) );
  inv01 U1736 ( .Y(n4896), .A(n4905) );
  nand02 U1737 ( .Y(n6442), .A0(n4906), .A1(n4907) );
  inv01 U1738 ( .Y(n4909), .A(n5014) );
  inv01 U1739 ( .Y(n4910), .A(opa_i[20]) );
  nand02 U1740 ( .Y(n4906), .A0(n4908), .A1(n4909) );
  nand02 U1741 ( .Y(n4907), .A0(n4908), .A1(n4910) );
  nand02 U1742 ( .Y(n6342), .A0(n4911), .A1(n4912) );
  inv01 U1743 ( .Y(n4913), .A(opa_i[16]) );
  inv01 U1744 ( .Y(n4914), .A(n6137) );
  inv01 U1745 ( .Y(n4915), .A(n6309) );
  nand02 U1746 ( .Y(n4916), .A0(n4913), .A1(n5928) );
  nand02 U1747 ( .Y(n4917), .A0(n4913), .A1(n4914) );
  nand02 U1748 ( .Y(n4918), .A0(n5928), .A1(n4915) );
  nand02 U1749 ( .Y(n4919), .A0(n4914), .A1(n4915) );
  nand02 U1750 ( .Y(n4920), .A0(n4916), .A1(n4917) );
  inv01 U1751 ( .Y(n4911), .A(n4920) );
  nand02 U1752 ( .Y(n4921), .A0(n4918), .A1(n4919) );
  inv01 U1753 ( .Y(n4912), .A(n4921) );
  nand02 U1754 ( .Y(n6169), .A0(n4922), .A1(n4923) );
  inv01 U1755 ( .Y(n4924), .A(n6141) );
  inv01 U1756 ( .Y(n4925), .A(opb_i[21]) );
  inv01 U1757 ( .Y(n4926), .A(n6140) );
  nand02 U1758 ( .Y(n4927), .A0(n6158), .A1(n4924) );
  nand02 U1759 ( .Y(n4928), .A0(n6158), .A1(n4925) );
  nand02 U1760 ( .Y(n4929), .A0(n4924), .A1(n4926) );
  nand02 U1761 ( .Y(n4930), .A0(n4925), .A1(n4926) );
  nand02 U1762 ( .Y(n4931), .A0(n4927), .A1(n4928) );
  inv01 U1763 ( .Y(n4922), .A(n4931) );
  nand02 U1764 ( .Y(n4932), .A0(n4929), .A1(n4930) );
  inv01 U1765 ( .Y(n4923), .A(n4932) );
  buf02 U1766 ( .Y(n4933), .A(opb_i[12]) );
  inv01 U1767 ( .Y(n4934), .A(n4933) );
  buf02 U1768 ( .Y(n4935), .A(opb_i[8]) );
  inv01 U1769 ( .Y(n4936), .A(n4935) );
  or03 U1770 ( .Y(n4937), .A0(n6404), .A1(n6383), .A2(n6384) );
  inv01 U1771 ( .Y(n4938), .A(n4937) );
  inv02 U1772 ( .Y(n6388), .A(n4939) );
  nand02 U1773 ( .Y(n4939), .A0(opa_i[4]), .A1(n4940) );
  nand02 U1774 ( .Y(n4941), .A0(n6429), .A1(n6076) );
  inv01 U1775 ( .Y(n4940), .A(n4941) );
  inv02 U1776 ( .Y(n6258), .A(n4942) );
  nand02 U1777 ( .Y(n4942), .A0(opb_i[16]), .A1(n4943) );
  nand02 U1778 ( .Y(n4944), .A0(n6292), .A1(n5931) );
  inv01 U1779 ( .Y(n4943), .A(n4944) );
  nand02 U1780 ( .Y(n6168), .A0(n4945), .A1(n4946) );
  inv01 U1781 ( .Y(n4947), .A(n6173) );
  inv01 U1782 ( .Y(n4948), .A(opb_i[19]) );
  inv01 U1783 ( .Y(n4949), .A(n6172) );
  inv01 U1784 ( .Y(n4950), .A(opb_i[22]) );
  nand02 U1785 ( .Y(n4951), .A0(n4947), .A1(n4948) );
  nand02 U1786 ( .Y(n4952), .A0(n4947), .A1(n4949) );
  nand02 U1787 ( .Y(n4953), .A0(n4948), .A1(n4950) );
  nand02 U1788 ( .Y(n4954), .A0(n4949), .A1(n4950) );
  nand02 U1789 ( .Y(n4955), .A0(n4951), .A1(n4952) );
  inv01 U1790 ( .Y(n4945), .A(n4955) );
  nand02 U1791 ( .Y(n4956), .A0(n4953), .A1(n4954) );
  inv01 U1792 ( .Y(n4946), .A(n4956) );
  nand02 U1793 ( .Y(n6186), .A0(n4957), .A1(n4958) );
  inv01 U1794 ( .Y(n4959), .A(opb_i[17]) );
  inv01 U1795 ( .Y(n4960), .A(n6172) );
  inv01 U1796 ( .Y(n4961), .A(n6173) );
  nand02 U1797 ( .Y(n4962), .A0(n6158), .A1(n4959) );
  nand02 U1798 ( .Y(n4963), .A0(n6158), .A1(n4960) );
  nand02 U1799 ( .Y(n4964), .A0(n4959), .A1(n4961) );
  nand02 U1800 ( .Y(n4965), .A0(n4960), .A1(n4961) );
  nand02 U1801 ( .Y(n4966), .A0(n4962), .A1(n4963) );
  inv01 U1802 ( .Y(n4957), .A(n4966) );
  nand02 U1803 ( .Y(n4967), .A0(n4964), .A1(n4965) );
  inv01 U1804 ( .Y(n4958), .A(n4967) );
  nand02 U1805 ( .Y(n6179), .A0(n4968), .A1(n4969) );
  inv01 U1806 ( .Y(n4970), .A(n6173) );
  inv01 U1807 ( .Y(n4971), .A(opb_i[18]) );
  inv01 U1808 ( .Y(n4972), .A(n6172) );
  inv01 U1809 ( .Y(n4973), .A(opb_i[21]) );
  nand02 U1810 ( .Y(n4974), .A0(n4970), .A1(n4971) );
  nand02 U1811 ( .Y(n4975), .A0(n4970), .A1(n4972) );
  nand02 U1812 ( .Y(n4976), .A0(n4971), .A1(n4973) );
  nand02 U1813 ( .Y(n4977), .A0(n4972), .A1(n4973) );
  nand02 U1814 ( .Y(n4978), .A0(n4974), .A1(n4975) );
  inv01 U1815 ( .Y(n4968), .A(n4978) );
  nand02 U1816 ( .Y(n4979), .A0(n4976), .A1(n4977) );
  inv01 U1817 ( .Y(n4969), .A(n4979) );
  nand02 U1818 ( .Y(n6187), .A0(n4980), .A1(n4981) );
  inv01 U1819 ( .Y(n4982), .A(opb_i[19]) );
  inv01 U1820 ( .Y(n4983), .A(n6141) );
  inv01 U1821 ( .Y(n4984), .A(n6140) );
  nand02 U1822 ( .Y(n4985), .A0(n4364), .A1(n4982) );
  nand02 U1823 ( .Y(n4986), .A0(n4364), .A1(n4983) );
  nand02 U1824 ( .Y(n4987), .A0(n4982), .A1(n4984) );
  nand02 U1825 ( .Y(n4988), .A0(n4983), .A1(n4984) );
  nand02 U1826 ( .Y(n4989), .A0(n4985), .A1(n4986) );
  inv01 U1827 ( .Y(n4980), .A(n4989) );
  nand02 U1828 ( .Y(n4990), .A0(n4987), .A1(n4988) );
  inv01 U1829 ( .Y(n4981), .A(n4990) );
  buf02 U1830 ( .Y(n4991), .A(opb_i[4]) );
  inv01 U1831 ( .Y(n4992), .A(n4991) );
  inv02 U1832 ( .Y(n6261), .A(n4993) );
  nand02 U1833 ( .Y(n4993), .A0(opb_i[2]), .A1(n4994) );
  nand02 U1834 ( .Y(n4995), .A0(n6296), .A1(n6053) );
  inv01 U1835 ( .Y(n4994), .A(n4995) );
  inv02 U1836 ( .Y(n6260), .A(n4996) );
  nand02 U1837 ( .Y(n4996), .A0(opb_i[10]), .A1(n4997) );
  nand02 U1838 ( .Y(n4998), .A0(n6295), .A1(n6055) );
  inv01 U1839 ( .Y(n4997), .A(n4998) );
  nand02 U1840 ( .Y(n6180), .A0(n4999), .A1(n5000) );
  inv01 U1841 ( .Y(n5001), .A(opb_i[19]) );
  inv01 U1842 ( .Y(n5002), .A(n6141) );
  inv01 U1843 ( .Y(n5003), .A(n6140) );
  nand02 U1844 ( .Y(n5004), .A0(n5001), .A1(n6158) );
  nand02 U1845 ( .Y(n5005), .A0(n5001), .A1(n5002) );
  nand02 U1846 ( .Y(n5006), .A0(n6158), .A1(n5003) );
  nand02 U1847 ( .Y(n5007), .A0(n5002), .A1(n5003) );
  nand02 U1848 ( .Y(n5008), .A0(n5004), .A1(n5005) );
  inv01 U1849 ( .Y(n4999), .A(n5008) );
  nand02 U1850 ( .Y(n5009), .A0(n5006), .A1(n5007) );
  inv01 U1851 ( .Y(n5000), .A(n5009) );
  nand02 U1852 ( .Y(n6306), .A0(n5010), .A1(n5011) );
  inv01 U1853 ( .Y(n5012), .A(n6083) );
  inv01 U1854 ( .Y(n5013), .A(n5926) );
  nand02 U1855 ( .Y(n5015), .A0(n5012), .A1(n5013) );
  nand02 U1856 ( .Y(n5016), .A0(n5012), .A1(n5014) );
  nand02 U1857 ( .Y(n5017), .A0(n5013), .A1(n4908) );
  nand02 U1858 ( .Y(n5018), .A0(n5014), .A1(n4908) );
  nand02 U1859 ( .Y(n5019), .A0(n5015), .A1(n5016) );
  inv01 U1860 ( .Y(n5010), .A(n5019) );
  nand02 U1861 ( .Y(n5020), .A0(n5017), .A1(n5018) );
  inv01 U1862 ( .Y(n5011), .A(n5020) );
  inv02 U1863 ( .Y(n6257), .A(n5021) );
  nand02 U1864 ( .Y(n5021), .A0(opb_i[12]), .A1(n5022) );
  nand02 U1865 ( .Y(n5023), .A0(n5037), .A1(n6046) );
  inv01 U1866 ( .Y(n5022), .A(n5023) );
  buf02 U1867 ( .Y(n5024), .A(opb_i[16]) );
  inv01 U1868 ( .Y(n5025), .A(n5024) );
  buf02 U1869 ( .Y(n5026), .A(opa_i[13]) );
  inv01 U1870 ( .Y(n5027), .A(n5026) );
  buf02 U1871 ( .Y(n5028), .A(opa_i[6]) );
  inv01 U1872 ( .Y(n5029), .A(n5028) );
  inv02 U1873 ( .Y(n6435), .A(n5030) );
  nand02 U1874 ( .Y(n5030), .A0(n5091), .A1(n5031) );
  nand02 U1875 ( .Y(n5032), .A0(n5027), .A1(n6080) );
  inv02 U1876 ( .Y(n5031), .A(n5032) );
  inv02 U1877 ( .Y(n6429), .A(n5033) );
  nand02 U1878 ( .Y(n5033), .A0(n5093), .A1(n5034) );
  nand02 U1879 ( .Y(n5035), .A0(n5029), .A1(n6072) );
  inv02 U1880 ( .Y(n5034), .A(n5035) );
  nand03 U1881 ( .Y(n5036), .A0(n5162), .A1(n6059), .A2(n6294) );
  inv02 U1882 ( .Y(n5037), .A(n5036) );
  inv02 U1883 ( .Y(n6262), .A(n5038) );
  nand02 U1884 ( .Y(n5038), .A0(opb_i[4]), .A1(n5039) );
  nand02 U1885 ( .Y(n5040), .A0(n4685), .A1(n6057) );
  inv01 U1886 ( .Y(n5039), .A(n5040) );
  or03 U1887 ( .Y(n5041), .A0(n6275), .A1(n6263), .A2(n6266) );
  inv02 U1888 ( .Y(n5042), .A(n5041) );
  nand02 U1889 ( .Y(n6322), .A0(n5043), .A1(n5044) );
  inv01 U1890 ( .Y(n5045), .A(n6137) );
  inv01 U1891 ( .Y(n5046), .A(n6309) );
  nand02 U1892 ( .Y(n5047), .A0(n6007), .A1(n6010) );
  nand02 U1893 ( .Y(n5048), .A0(n6007), .A1(n5045) );
  nand02 U1894 ( .Y(n5049), .A0(n6011), .A1(n5046) );
  nand02 U1895 ( .Y(n5050), .A0(n5045), .A1(n5046) );
  nand02 U1896 ( .Y(n5051), .A0(n5047), .A1(n5048) );
  inv01 U1897 ( .Y(n5043), .A(n5051) );
  nand02 U1898 ( .Y(n5052), .A0(n5049), .A1(n5050) );
  inv01 U1899 ( .Y(n5044), .A(n5052) );
  nand02 U1900 ( .Y(n6321), .A0(n5053), .A1(n5054) );
  inv01 U1901 ( .Y(n5055), .A(n5926) );
  inv01 U1902 ( .Y(n5056), .A(n6083) );
  nand02 U1903 ( .Y(n5057), .A0(n5086), .A1(n5077) );
  nand02 U1904 ( .Y(n5058), .A0(n5086), .A1(n5055) );
  nand02 U1905 ( .Y(n5059), .A0(n6030), .A1(n5056) );
  nand02 U1906 ( .Y(n5060), .A0(n5055), .A1(n5056) );
  nand02 U1907 ( .Y(n5061), .A0(n5057), .A1(n5058) );
  inv01 U1908 ( .Y(n5053), .A(n5061) );
  nand02 U1909 ( .Y(n5062), .A0(n5059), .A1(n5060) );
  inv01 U1910 ( .Y(n5054), .A(n5062) );
  inv02 U1911 ( .Y(n____return3540_0_), .A(s_expa_in_0_) );
  ao22 U1912 ( .Y(n5063), .A0(n5926), .A1(opa_i[20]), .B0(opa_i[21]), .B1(
        n6083) );
  inv01 U1913 ( .Y(n5064), .A(n5063) );
  nand02 U1914 ( .Y(n6307), .A0(n5065), .A1(n5066) );
  inv01 U1915 ( .Y(n5067), .A(n6137) );
  inv01 U1916 ( .Y(n5068), .A(n6309) );
  nand02 U1917 ( .Y(n5069), .A0(n5086), .A1(n6030) );
  nand02 U1918 ( .Y(n5070), .A0(n6297), .A1(n5067) );
  nand02 U1919 ( .Y(n5071), .A0(n5077), .A1(n5068) );
  nand02 U1920 ( .Y(n5072), .A0(n5067), .A1(n5068) );
  nand02 U1921 ( .Y(n5073), .A0(n5069), .A1(n5070) );
  inv01 U1922 ( .Y(n5065), .A(n5073) );
  nand02 U1923 ( .Y(n5074), .A0(n5071), .A1(n5072) );
  inv01 U1924 ( .Y(n5066), .A(n5074) );
  nand02 U1925 ( .Y(n6315), .A0(n5075), .A1(n5076) );
  inv01 U1926 ( .Y(n5078), .A(n6137) );
  inv01 U1927 ( .Y(n5079), .A(n6309) );
  nand02 U1928 ( .Y(n5080), .A0(n5077), .A1(n6007) );
  nand02 U1929 ( .Y(n5081), .A0(n5077), .A1(n5078) );
  nand02 U1930 ( .Y(n5082), .A0(n6007), .A1(n5079) );
  nand02 U1931 ( .Y(n5083), .A0(n5078), .A1(n5079) );
  nand02 U1932 ( .Y(n5084), .A0(n5080), .A1(n5081) );
  inv01 U1933 ( .Y(n5075), .A(n5084) );
  nand02 U1934 ( .Y(n5085), .A0(n5082), .A1(n5083) );
  inv01 U1935 ( .Y(n5076), .A(n5085) );
  buf02 U1936 ( .Y(n5086), .A(n6297) );
  or03 U1937 ( .Y(n5087), .A0(n6109), .A1(s_dvd_zeros_3_), .A2(n5918) );
  inv01 U1938 ( .Y(dvdnd_50_o[30]), .A(n5087) );
  or03 U1939 ( .Y(n5089), .A0(n6118), .A1(n6081), .A2(n5914) );
  inv01 U1940 ( .Y(dvsor_27_o[4]), .A(n5089) );
  buf02 U1941 ( .Y(n5091), .A(n6434) );
  buf02 U1942 ( .Y(n5092), .A(n6434) );
  buf02 U1943 ( .Y(n5093), .A(n6436) );
  buf02 U1944 ( .Y(n5094), .A(n6436) );
  inv01 U1945 ( .Y(dvdnd_50_o[38]), .A(n5095) );
  nor02 U1946 ( .Y(n5096), .A0(n6350), .A1(n6136) );
  nor02 U1947 ( .Y(n5097), .A0(n6349), .A1(n6121) );
  nor02 U1948 ( .Y(n5098), .A0(n5918), .A1(n5566) );
  nor02 U1949 ( .Y(n5095), .A0(n5098), .A1(n5099) );
  nor02 U1950 ( .Y(n5100), .A0(n5096), .A1(n5097) );
  inv01 U1951 ( .Y(n5099), .A(n5100) );
  inv01 U1952 ( .Y(dvdnd_50_o[37]), .A(n5101) );
  nor02 U1953 ( .Y(n5102), .A0(n6365), .A1(n6136) );
  nor02 U1954 ( .Y(n5103), .A0(n6328), .A1(n6121) );
  nor02 U1955 ( .Y(n5104), .A0(n6357), .A1(n6132) );
  nor02 U1956 ( .Y(n5101), .A0(n5104), .A1(n5105) );
  nor02 U1957 ( .Y(n5106), .A0(n5102), .A1(n5103) );
  inv01 U1958 ( .Y(n5105), .A(n5106) );
  inv01 U1959 ( .Y(dvdnd_50_o[35]), .A(n5107) );
  nor02 U1960 ( .Y(n5108), .A0(n6362), .A1(n6136) );
  nor02 U1961 ( .Y(n5109), .A0(n6344), .A1(n6120) );
  nor02 U1962 ( .Y(n5110), .A0(n6369), .A1(n6132) );
  nor02 U1963 ( .Y(n5107), .A0(n5110), .A1(n5111) );
  nor02 U1964 ( .Y(n5112), .A0(n5108), .A1(n5109) );
  inv01 U1965 ( .Y(n5111), .A(n5112) );
  inv01 U1966 ( .Y(dvdnd_50_o[36]), .A(n5113) );
  nor02 U1967 ( .Y(n5114), .A0(n6360), .A1(n6136) );
  nor02 U1968 ( .Y(n5115), .A0(n6338), .A1(n6121) );
  nor02 U1969 ( .Y(n5116), .A0(n6367), .A1(n6132) );
  nor02 U1970 ( .Y(n5113), .A0(n5116), .A1(n5117) );
  nor02 U1971 ( .Y(n5118), .A0(n5114), .A1(n5115) );
  inv01 U1972 ( .Y(n5117), .A(n5118) );
  inv01 U1973 ( .Y(n6362), .A(n6347) );
  inv01 U1974 ( .Y(dvsor_27_o[12]), .A(n5119) );
  nor02 U1975 ( .Y(n5120), .A0(n6151), .A1(n6134) );
  nor02 U1976 ( .Y(n5121), .A0(n5914), .A1(n5678) );
  nor02 U1977 ( .Y(n5122), .A0(n6215), .A1(n6130) );
  nor02 U1978 ( .Y(n5119), .A0(n5122), .A1(n5123) );
  nor02 U1979 ( .Y(n5124), .A0(n5120), .A1(n5121) );
  inv01 U1980 ( .Y(n5123), .A(n5124) );
  inv01 U1981 ( .Y(dvsor_27_o[11]), .A(n5125) );
  nor02 U1982 ( .Y(n5126), .A0(n6194), .A1(n6129) );
  nor02 U1983 ( .Y(n5127), .A0(n6156), .A1(n6126) );
  nor02 U1984 ( .Y(n5128), .A0(n6166), .A1(n6134) );
  nor02 U1985 ( .Y(n5125), .A0(n5128), .A1(n5129) );
  nor02 U1986 ( .Y(n5130), .A0(n5126), .A1(n5127) );
  inv01 U1987 ( .Y(n5129), .A(n5130) );
  inv01 U1988 ( .Y(dvsor_27_o[10]), .A(n5131) );
  nor02 U1989 ( .Y(n5132), .A0(n6176), .A1(n6134) );
  nor02 U1990 ( .Y(n5133), .A0(n6084), .A1(n6126) );
  nor02 U1991 ( .Y(n5134), .A0(n6204), .A1(n6128) );
  nor02 U1992 ( .Y(n5131), .A0(n5134), .A1(n5135) );
  nor02 U1993 ( .Y(n5136), .A0(n5132), .A1(n5133) );
  inv01 U1994 ( .Y(n5135), .A(n5136) );
  inv01 U1995 ( .Y(dvsor_27_o[9]), .A(n5137) );
  nor02 U1996 ( .Y(n5138), .A0(n6148), .A1(n6129) );
  nor02 U1997 ( .Y(n5139), .A0(n6026), .A1(n6126) );
  nor02 U1998 ( .Y(n5140), .A0(n6147), .A1(n6134) );
  nor02 U1999 ( .Y(n5137), .A0(n5140), .A1(n5141) );
  nor02 U2000 ( .Y(n5142), .A0(n5138), .A1(n5139) );
  inv01 U2001 ( .Y(n5141), .A(n5142) );
  inv01 U2002 ( .Y(dvsor_27_o[8]), .A(n5143) );
  nor02 U2003 ( .Y(n5144), .A0(n6151), .A1(n6129) );
  nor02 U2004 ( .Y(n5145), .A0(n6126), .A1(n5163) );
  nor02 U2005 ( .Y(n5146), .A0(n6149), .A1(n6134) );
  nor02 U2006 ( .Y(n5143), .A0(n5146), .A1(n5147) );
  nor02 U2007 ( .Y(n5148), .A0(n5144), .A1(n5145) );
  inv01 U2008 ( .Y(n5147), .A(n5148) );
  buf02 U2009 ( .Y(n5163), .A(n6150) );
  inv01 U2010 ( .Y(dvdnd_50_o[34]), .A(n5149) );
  nor02 U2011 ( .Y(n5150), .A0(n6373), .A1(n6136) );
  nor02 U2012 ( .Y(n5151), .A0(n6132), .A1(n5699) );
  nor02 U2013 ( .Y(n5152), .A0(n6350), .A1(n6120) );
  nor02 U2014 ( .Y(n5149), .A0(n5152), .A1(n5153) );
  nor02 U2015 ( .Y(n5154), .A0(n5150), .A1(n5151) );
  inv01 U2016 ( .Y(n5153), .A(n5154) );
  inv02 U2017 ( .Y(n6120), .A(n6119) );
  inv04 U2018 ( .Y(n6136), .A(n6135) );
  inv01 U2019 ( .Y(n5155), .A(n5850) );
  buf02 U2020 ( .Y(n5156), .A(opb_i[10]) );
  inv02 U2021 ( .Y(n5157), .A(n5156) );
  nand03 U2022 ( .Y(n5158), .A0(n5673), .A1(n6078), .A2(n6437) );
  inv02 U2023 ( .Y(n5159), .A(n5158) );
  nand03 U2024 ( .Y(n5160), .A0(n6223), .A1(n6053), .A2(n6296) );
  inv02 U2025 ( .Y(n5161), .A(n5160) );
  inv01 U2026 ( .Y(n5162), .A(n5788) );
  ao32 U2027 ( .Y(n5164), .A0(n6189), .A1(n6098), .A2(n6163), .B0(n6123), .B1(
        n6190) );
  inv01 U2028 ( .Y(n5165), .A(n5164) );
  nand02 U2029 ( .Y(n6205), .A0(n5166), .A1(n5167) );
  inv02 U2030 ( .Y(n5168), .A(n6177) );
  inv02 U2031 ( .Y(n5169), .A(n6207) );
  inv02 U2032 ( .Y(n5170), .A(n6206) );
  inv02 U2033 ( .Y(n5171), .A(n5912) );
  inv02 U2034 ( .Y(n5172), .A(n6123) );
  inv02 U2035 ( .Y(n5173), .A(n6199) );
  nand02 U2036 ( .Y(n5174), .A0(n5170), .A1(n5175) );
  nand02 U2037 ( .Y(n5176), .A0(n5171), .A1(n5177) );
  nand02 U2038 ( .Y(n5178), .A0(n5172), .A1(n5179) );
  nand02 U2039 ( .Y(n5180), .A0(n5172), .A1(n5181) );
  nand02 U2040 ( .Y(n5182), .A0(n5173), .A1(n5183) );
  nand02 U2041 ( .Y(n5184), .A0(n5173), .A1(n5185) );
  nand02 U2042 ( .Y(n5186), .A0(n5173), .A1(n5187) );
  nand02 U2043 ( .Y(n5188), .A0(n5173), .A1(n5189) );
  nand02 U2044 ( .Y(n5190), .A0(n5168), .A1(n5169) );
  inv01 U2045 ( .Y(n5175), .A(n5190) );
  nand02 U2046 ( .Y(n5191), .A0(n5168), .A1(n5169) );
  inv01 U2047 ( .Y(n5177), .A(n5191) );
  nand02 U2048 ( .Y(n5192), .A0(n5168), .A1(n5170) );
  inv01 U2049 ( .Y(n5179), .A(n5192) );
  nand02 U2050 ( .Y(n5193), .A0(n5168), .A1(n5171) );
  inv01 U2051 ( .Y(n5181), .A(n5193) );
  nand02 U2052 ( .Y(n5194), .A0(n5169), .A1(n5170) );
  inv01 U2053 ( .Y(n5183), .A(n5194) );
  nand02 U2054 ( .Y(n5195), .A0(n5169), .A1(n5171) );
  inv01 U2055 ( .Y(n5185), .A(n5195) );
  nand02 U2056 ( .Y(n5196), .A0(n5170), .A1(n5172) );
  inv01 U2057 ( .Y(n5187), .A(n5196) );
  nand02 U2058 ( .Y(n5197), .A0(n5171), .A1(n5172) );
  inv01 U2059 ( .Y(n5189), .A(n5197) );
  nand02 U2060 ( .Y(n5198), .A0(n5174), .A1(n5176) );
  inv01 U2061 ( .Y(n5199), .A(n5198) );
  nand02 U2062 ( .Y(n5200), .A0(n5178), .A1(n5180) );
  inv01 U2063 ( .Y(n5201), .A(n5200) );
  nand02 U2064 ( .Y(n5202), .A0(n5199), .A1(n5201) );
  inv01 U2065 ( .Y(n5166), .A(n5202) );
  nand02 U2066 ( .Y(n5203), .A0(n5182), .A1(n5184) );
  inv01 U2067 ( .Y(n5204), .A(n5203) );
  nand02 U2068 ( .Y(n5205), .A0(n5186), .A1(n5188) );
  inv01 U2069 ( .Y(n5206), .A(n5205) );
  nand02 U2070 ( .Y(n5207), .A0(n5204), .A1(n5206) );
  inv01 U2071 ( .Y(n5167), .A(n5207) );
  nand02 U2072 ( .Y(n6195), .A0(n5208), .A1(n5209) );
  inv02 U2073 ( .Y(n5210), .A(n6160) );
  inv02 U2074 ( .Y(n5211), .A(n6198) );
  inv02 U2075 ( .Y(n5212), .A(n6197) );
  inv02 U2076 ( .Y(n5213), .A(n5912) );
  inv02 U2077 ( .Y(n5214), .A(n6123) );
  inv02 U2078 ( .Y(n5215), .A(n6199) );
  nand02 U2079 ( .Y(n5216), .A0(n5212), .A1(n5217) );
  nand02 U2080 ( .Y(n5218), .A0(n5213), .A1(n5219) );
  nand02 U2081 ( .Y(n5220), .A0(n5214), .A1(n5221) );
  nand02 U2082 ( .Y(n5222), .A0(n5214), .A1(n5223) );
  nand02 U2083 ( .Y(n5224), .A0(n5215), .A1(n5225) );
  nand02 U2084 ( .Y(n5226), .A0(n5215), .A1(n5227) );
  nand02 U2085 ( .Y(n5228), .A0(n5215), .A1(n5229) );
  nand02 U2086 ( .Y(n5230), .A0(n5215), .A1(n5231) );
  nand02 U2087 ( .Y(n5232), .A0(n5210), .A1(n5211) );
  inv01 U2088 ( .Y(n5217), .A(n5232) );
  nand02 U2089 ( .Y(n5233), .A0(n5210), .A1(n5211) );
  inv01 U2090 ( .Y(n5219), .A(n5233) );
  nand02 U2091 ( .Y(n5234), .A0(n5210), .A1(n5212) );
  inv01 U2092 ( .Y(n5221), .A(n5234) );
  nand02 U2093 ( .Y(n5235), .A0(n5210), .A1(n5213) );
  inv01 U2094 ( .Y(n5223), .A(n5235) );
  nand02 U2095 ( .Y(n5236), .A0(n5211), .A1(n5212) );
  inv01 U2096 ( .Y(n5225), .A(n5236) );
  nand02 U2097 ( .Y(n5237), .A0(n5211), .A1(n5213) );
  inv01 U2098 ( .Y(n5227), .A(n5237) );
  nand02 U2099 ( .Y(n5238), .A0(n5212), .A1(n5214) );
  inv01 U2100 ( .Y(n5229), .A(n5238) );
  nand02 U2101 ( .Y(n5239), .A0(n5213), .A1(n5214) );
  inv01 U2102 ( .Y(n5231), .A(n5239) );
  nand02 U2103 ( .Y(n5240), .A0(n5216), .A1(n5218) );
  inv01 U2104 ( .Y(n5241), .A(n5240) );
  nand02 U2105 ( .Y(n5242), .A0(n5220), .A1(n5222) );
  inv01 U2106 ( .Y(n5243), .A(n5242) );
  nand02 U2107 ( .Y(n5244), .A0(n5241), .A1(n5243) );
  inv01 U2108 ( .Y(n5208), .A(n5244) );
  nand02 U2109 ( .Y(n5245), .A0(n5224), .A1(n5226) );
  inv01 U2110 ( .Y(n5246), .A(n5245) );
  nand02 U2111 ( .Y(n5247), .A0(n5228), .A1(n5230) );
  inv01 U2112 ( .Y(n5248), .A(n5247) );
  nand02 U2113 ( .Y(n5249), .A0(n5246), .A1(n5248) );
  inv01 U2114 ( .Y(n5209), .A(n5249) );
  inv04 U2115 ( .Y(n6199), .A(n6102) );
  nand02 U2116 ( .Y(n6339), .A0(n5250), .A1(n5251) );
  inv02 U2117 ( .Y(n5252), .A(n6313) );
  inv02 U2118 ( .Y(n5253), .A(n6341) );
  inv02 U2119 ( .Y(n5254), .A(n6340) );
  inv02 U2120 ( .Y(n5255), .A(n6330) );
  inv02 U2121 ( .Y(n5256), .A(n6124) );
  inv02 U2122 ( .Y(n5257), .A(n6333) );
  nand02 U2123 ( .Y(n5258), .A0(n5254), .A1(n5259) );
  nand02 U2124 ( .Y(n5260), .A0(n5255), .A1(n5261) );
  nand02 U2125 ( .Y(n5262), .A0(n5256), .A1(n5263) );
  nand02 U2126 ( .Y(n5264), .A0(n5256), .A1(n5265) );
  nand02 U2127 ( .Y(n5266), .A0(n5257), .A1(n5267) );
  nand02 U2128 ( .Y(n5268), .A0(n5257), .A1(n5269) );
  nand02 U2129 ( .Y(n5270), .A0(n5257), .A1(n5271) );
  nand02 U2130 ( .Y(n5272), .A0(n5257), .A1(n5273) );
  nand02 U2131 ( .Y(n5274), .A0(n5252), .A1(n5253) );
  inv01 U2132 ( .Y(n5259), .A(n5274) );
  nand02 U2133 ( .Y(n5275), .A0(n5252), .A1(n5253) );
  inv01 U2134 ( .Y(n5261), .A(n5275) );
  nand02 U2135 ( .Y(n5276), .A0(n5252), .A1(n5254) );
  inv01 U2136 ( .Y(n5263), .A(n5276) );
  nand02 U2137 ( .Y(n5277), .A0(n5252), .A1(n5255) );
  inv01 U2138 ( .Y(n5265), .A(n5277) );
  nand02 U2139 ( .Y(n5278), .A0(n5253), .A1(n5254) );
  inv01 U2140 ( .Y(n5267), .A(n5278) );
  nand02 U2141 ( .Y(n5279), .A0(n5253), .A1(n5255) );
  inv01 U2142 ( .Y(n5269), .A(n5279) );
  nand02 U2143 ( .Y(n5280), .A0(n5254), .A1(n5256) );
  inv01 U2144 ( .Y(n5271), .A(n5280) );
  nand02 U2145 ( .Y(n5281), .A0(n5255), .A1(n5256) );
  inv01 U2146 ( .Y(n5273), .A(n5281) );
  nand02 U2147 ( .Y(n5282), .A0(n5258), .A1(n5260) );
  inv01 U2148 ( .Y(n5283), .A(n5282) );
  nand02 U2149 ( .Y(n5284), .A0(n5262), .A1(n5264) );
  inv01 U2150 ( .Y(n5285), .A(n5284) );
  nand02 U2151 ( .Y(n5286), .A0(n5283), .A1(n5285) );
  inv01 U2152 ( .Y(n5250), .A(n5286) );
  nand02 U2153 ( .Y(n5287), .A0(n5266), .A1(n5268) );
  inv01 U2154 ( .Y(n5288), .A(n5287) );
  nand02 U2155 ( .Y(n5289), .A0(n5270), .A1(n5272) );
  inv01 U2156 ( .Y(n5290), .A(n5289) );
  nand02 U2157 ( .Y(n5291), .A0(n5288), .A1(n5290) );
  inv01 U2158 ( .Y(n5251), .A(n5291) );
  nand02 U2159 ( .Y(n6345), .A0(n5292), .A1(n5293) );
  inv02 U2160 ( .Y(n5294), .A(n6319) );
  inv02 U2161 ( .Y(n5295), .A(n6347) );
  inv02 U2162 ( .Y(n5296), .A(n6346) );
  inv02 U2163 ( .Y(n5297), .A(n6330) );
  inv02 U2164 ( .Y(n5298), .A(n6124) );
  inv02 U2165 ( .Y(n5299), .A(n6333) );
  nand02 U2166 ( .Y(n5300), .A0(n5296), .A1(n5301) );
  nand02 U2167 ( .Y(n5302), .A0(n5297), .A1(n5303) );
  nand02 U2168 ( .Y(n5304), .A0(n5298), .A1(n5305) );
  nand02 U2169 ( .Y(n5306), .A0(n5298), .A1(n5307) );
  nand02 U2170 ( .Y(n5308), .A0(n5299), .A1(n5309) );
  nand02 U2171 ( .Y(n5310), .A0(n5299), .A1(n5311) );
  nand02 U2172 ( .Y(n5312), .A0(n5299), .A1(n5313) );
  nand02 U2173 ( .Y(n5314), .A0(n5299), .A1(n5315) );
  nand02 U2174 ( .Y(n5316), .A0(n5294), .A1(n5295) );
  inv01 U2175 ( .Y(n5301), .A(n5316) );
  nand02 U2176 ( .Y(n5317), .A0(n5294), .A1(n5295) );
  inv01 U2177 ( .Y(n5303), .A(n5317) );
  nand02 U2178 ( .Y(n5318), .A0(n5294), .A1(n5296) );
  inv01 U2179 ( .Y(n5305), .A(n5318) );
  nand02 U2180 ( .Y(n5319), .A0(n5294), .A1(n5297) );
  inv01 U2181 ( .Y(n5307), .A(n5319) );
  nand02 U2182 ( .Y(n5320), .A0(n5295), .A1(n5296) );
  inv01 U2183 ( .Y(n5309), .A(n5320) );
  nand02 U2184 ( .Y(n5321), .A0(n5295), .A1(n5297) );
  inv01 U2185 ( .Y(n5311), .A(n5321) );
  nand02 U2186 ( .Y(n5322), .A0(n5296), .A1(n5298) );
  inv01 U2187 ( .Y(n5313), .A(n5322) );
  nand02 U2188 ( .Y(n5323), .A0(n5297), .A1(n5298) );
  inv01 U2189 ( .Y(n5315), .A(n5323) );
  nand02 U2190 ( .Y(n5324), .A0(n5300), .A1(n5302) );
  inv01 U2191 ( .Y(n5325), .A(n5324) );
  nand02 U2192 ( .Y(n5326), .A0(n5304), .A1(n5306) );
  inv01 U2193 ( .Y(n5327), .A(n5326) );
  nand02 U2194 ( .Y(n5328), .A0(n5325), .A1(n5327) );
  inv01 U2195 ( .Y(n5292), .A(n5328) );
  nand02 U2196 ( .Y(n5329), .A0(n5308), .A1(n5310) );
  inv01 U2197 ( .Y(n5330), .A(n5329) );
  nand02 U2198 ( .Y(n5331), .A0(n5312), .A1(n5314) );
  inv01 U2199 ( .Y(n5332), .A(n5331) );
  nand02 U2200 ( .Y(n5333), .A0(n5330), .A1(n5332) );
  inv01 U2201 ( .Y(n5293), .A(n5333) );
  nand02 U2202 ( .Y(n6210), .A0(n5334), .A1(n5335) );
  inv02 U2203 ( .Y(n5336), .A(n6184) );
  inv02 U2204 ( .Y(n5337), .A(n6183) );
  inv02 U2205 ( .Y(n5338), .A(n6211) );
  inv02 U2206 ( .Y(n5339), .A(n5912) );
  inv02 U2207 ( .Y(n5340), .A(n6123) );
  inv02 U2208 ( .Y(n5341), .A(n6199) );
  nand02 U2209 ( .Y(n5342), .A0(n5338), .A1(n5343) );
  nand02 U2210 ( .Y(n5344), .A0(n5339), .A1(n5345) );
  nand02 U2211 ( .Y(n5346), .A0(n5340), .A1(n5347) );
  nand02 U2212 ( .Y(n5348), .A0(n5340), .A1(n5349) );
  nand02 U2213 ( .Y(n5350), .A0(n5341), .A1(n5351) );
  nand02 U2214 ( .Y(n5352), .A0(n5341), .A1(n5353) );
  nand02 U2215 ( .Y(n5354), .A0(n5341), .A1(n5355) );
  nand02 U2216 ( .Y(n5356), .A0(n5341), .A1(n5357) );
  nand02 U2217 ( .Y(n5358), .A0(n5336), .A1(n5337) );
  inv01 U2218 ( .Y(n5343), .A(n5358) );
  nand02 U2219 ( .Y(n5359), .A0(n5336), .A1(n5337) );
  inv01 U2220 ( .Y(n5345), .A(n5359) );
  nand02 U2221 ( .Y(n5360), .A0(n5336), .A1(n5338) );
  inv01 U2222 ( .Y(n5347), .A(n5360) );
  nand02 U2223 ( .Y(n5361), .A0(n5336), .A1(n5339) );
  inv01 U2224 ( .Y(n5349), .A(n5361) );
  nand02 U2225 ( .Y(n5362), .A0(n5337), .A1(n5338) );
  inv01 U2226 ( .Y(n5351), .A(n5362) );
  nand02 U2227 ( .Y(n5363), .A0(n5337), .A1(n5339) );
  inv01 U2228 ( .Y(n5353), .A(n5363) );
  nand02 U2229 ( .Y(n5364), .A0(n5338), .A1(n5340) );
  inv01 U2230 ( .Y(n5355), .A(n5364) );
  nand02 U2231 ( .Y(n5365), .A0(n5339), .A1(n5340) );
  inv01 U2232 ( .Y(n5357), .A(n5365) );
  nand02 U2233 ( .Y(n5366), .A0(n5342), .A1(n5344) );
  inv01 U2234 ( .Y(n5367), .A(n5366) );
  nand02 U2235 ( .Y(n5368), .A0(n5346), .A1(n5348) );
  inv01 U2236 ( .Y(n5369), .A(n5368) );
  nand02 U2237 ( .Y(n5370), .A0(n5367), .A1(n5369) );
  inv01 U2238 ( .Y(n5334), .A(n5370) );
  nand02 U2239 ( .Y(n5371), .A0(n5350), .A1(n5352) );
  inv01 U2240 ( .Y(n5372), .A(n5371) );
  nand02 U2241 ( .Y(n5373), .A0(n5354), .A1(n5356) );
  inv01 U2242 ( .Y(n5374), .A(n5373) );
  nand02 U2243 ( .Y(n5375), .A0(n5372), .A1(n5374) );
  inv01 U2244 ( .Y(n5335), .A(n5375) );
  inv04 U2245 ( .Y(n6333), .A(n6112) );
  nand02 U2246 ( .Y(n6329), .A0(n5376), .A1(n5377) );
  inv02 U2247 ( .Y(n5378), .A(n6299) );
  inv02 U2248 ( .Y(n5379), .A(n6332) );
  inv02 U2249 ( .Y(n5380), .A(n6331) );
  inv02 U2250 ( .Y(n5381), .A(n6330) );
  inv02 U2251 ( .Y(n5382), .A(n6124) );
  inv02 U2252 ( .Y(n5383), .A(n6333) );
  nand02 U2253 ( .Y(n5384), .A0(n5380), .A1(n5385) );
  nand02 U2254 ( .Y(n5386), .A0(n5381), .A1(n5387) );
  nand02 U2255 ( .Y(n5388), .A0(n5382), .A1(n5389) );
  nand02 U2256 ( .Y(n5390), .A0(n5382), .A1(n5391) );
  nand02 U2257 ( .Y(n5392), .A0(n5383), .A1(n5393) );
  nand02 U2258 ( .Y(n5394), .A0(n5383), .A1(n5395) );
  nand02 U2259 ( .Y(n5396), .A0(n5383), .A1(n5397) );
  nand02 U2260 ( .Y(n5398), .A0(n5383), .A1(n5399) );
  nand02 U2261 ( .Y(n5400), .A0(n5378), .A1(n5379) );
  inv01 U2262 ( .Y(n5385), .A(n5400) );
  nand02 U2263 ( .Y(n5401), .A0(n5378), .A1(n5379) );
  inv01 U2264 ( .Y(n5387), .A(n5401) );
  nand02 U2265 ( .Y(n5402), .A0(n5378), .A1(n5380) );
  inv01 U2266 ( .Y(n5389), .A(n5402) );
  nand02 U2267 ( .Y(n5403), .A0(n5378), .A1(n5381) );
  inv01 U2268 ( .Y(n5391), .A(n5403) );
  nand02 U2269 ( .Y(n5404), .A0(n5379), .A1(n5380) );
  inv01 U2270 ( .Y(n5393), .A(n5404) );
  nand02 U2271 ( .Y(n5405), .A0(n5379), .A1(n5381) );
  inv01 U2272 ( .Y(n5395), .A(n5405) );
  nand02 U2273 ( .Y(n5406), .A0(n5380), .A1(n5382) );
  inv01 U2274 ( .Y(n5397), .A(n5406) );
  nand02 U2275 ( .Y(n5407), .A0(n5381), .A1(n5382) );
  inv01 U2276 ( .Y(n5399), .A(n5407) );
  nand02 U2277 ( .Y(n5408), .A0(n5384), .A1(n5386) );
  inv01 U2278 ( .Y(n5409), .A(n5408) );
  nand02 U2279 ( .Y(n5410), .A0(n5388), .A1(n5390) );
  inv01 U2280 ( .Y(n5411), .A(n5410) );
  nand02 U2281 ( .Y(n5412), .A0(n5409), .A1(n5411) );
  inv01 U2282 ( .Y(n5376), .A(n5412) );
  nand02 U2283 ( .Y(n5413), .A0(n5392), .A1(n5394) );
  inv01 U2284 ( .Y(n5414), .A(n5413) );
  nand02 U2285 ( .Y(n5415), .A0(n5396), .A1(n5398) );
  inv01 U2286 ( .Y(n5416), .A(n5415) );
  nand02 U2287 ( .Y(n5417), .A0(n5414), .A1(n5416) );
  inv01 U2288 ( .Y(n5377), .A(n5417) );
  ao32 U2289 ( .Y(n5418), .A0(n6323), .A1(n6092), .A2(n6302), .B0(n6124), .B1(
        n6324) );
  inv01 U2290 ( .Y(n5419), .A(n5418) );
  nand02 U2291 ( .Y(n6216), .A0(n5420), .A1(n5421) );
  inv02 U2292 ( .Y(n5422), .A(n6217) );
  inv02 U2293 ( .Y(n5423), .A(n6191) );
  inv02 U2294 ( .Y(n5424), .A(n6199) );
  inv02 U2295 ( .Y(n5425), .A(n5912) );
  inv02 U2296 ( .Y(n5426), .A(n6123) );
  nand02 U2297 ( .Y(n5427), .A0(n5423), .A1(n5428) );
  nand02 U2298 ( .Y(n5429), .A0(n5424), .A1(n5430) );
  nand02 U2299 ( .Y(n5431), .A0(n5425), .A1(n5432) );
  nand02 U2300 ( .Y(n5433), .A0(n5425), .A1(n5434) );
  nand02 U2301 ( .Y(n5435), .A0(n5426), .A1(n5436) );
  nand02 U2302 ( .Y(n5437), .A0(n5426), .A1(n5438) );
  nand02 U2303 ( .Y(n5439), .A0(n5426), .A1(n5440) );
  nand02 U2304 ( .Y(n5441), .A0(n5426), .A1(n5442) );
  nand02 U2305 ( .Y(n5443), .A0(n6149), .A1(n5422) );
  inv01 U2306 ( .Y(n5428), .A(n5443) );
  nand02 U2307 ( .Y(n5444), .A0(n6149), .A1(n5422) );
  inv01 U2308 ( .Y(n5430), .A(n5444) );
  nand02 U2309 ( .Y(n5445), .A0(n6149), .A1(n5423) );
  inv01 U2310 ( .Y(n5432), .A(n5445) );
  nand02 U2311 ( .Y(n5446), .A0(n6149), .A1(n5424) );
  inv01 U2312 ( .Y(n5434), .A(n5446) );
  nand02 U2313 ( .Y(n5447), .A0(n5422), .A1(n5423) );
  inv01 U2314 ( .Y(n5436), .A(n5447) );
  nand02 U2315 ( .Y(n5448), .A0(n5422), .A1(n5424) );
  inv01 U2316 ( .Y(n5438), .A(n5448) );
  nand02 U2317 ( .Y(n5449), .A0(n5423), .A1(n5425) );
  inv01 U2318 ( .Y(n5440), .A(n5449) );
  nand02 U2319 ( .Y(n5450), .A0(n5424), .A1(n5425) );
  inv01 U2320 ( .Y(n5442), .A(n5450) );
  nand02 U2321 ( .Y(n5451), .A0(n5427), .A1(n5429) );
  inv01 U2322 ( .Y(n5452), .A(n5451) );
  nand02 U2323 ( .Y(n5453), .A0(n5431), .A1(n5433) );
  inv01 U2324 ( .Y(n5454), .A(n5453) );
  nand02 U2325 ( .Y(n5455), .A0(n5452), .A1(n5454) );
  inv01 U2326 ( .Y(n5420), .A(n5455) );
  nand02 U2327 ( .Y(n5456), .A0(n5435), .A1(n5437) );
  inv01 U2328 ( .Y(n5457), .A(n5456) );
  nand02 U2329 ( .Y(n5458), .A0(n5439), .A1(n5441) );
  inv01 U2330 ( .Y(n5459), .A(n5458) );
  nand02 U2331 ( .Y(n5460), .A0(n5457), .A1(n5459) );
  inv01 U2332 ( .Y(n5421), .A(n5460) );
  nand02 U2333 ( .Y(n6351), .A0(n5461), .A1(n5462) );
  inv02 U2334 ( .Y(n5463), .A(n6353) );
  inv02 U2335 ( .Y(n5464), .A(n6352) );
  inv02 U2336 ( .Y(n5465), .A(n6325) );
  inv02 U2337 ( .Y(n5466), .A(n6333) );
  inv02 U2338 ( .Y(n5467), .A(n6330) );
  inv02 U2339 ( .Y(n5468), .A(n6124) );
  nand02 U2340 ( .Y(n5469), .A0(n5465), .A1(n5470) );
  nand02 U2341 ( .Y(n5471), .A0(n5466), .A1(n5472) );
  nand02 U2342 ( .Y(n5473), .A0(n5467), .A1(n5474) );
  nand02 U2343 ( .Y(n5475), .A0(n5467), .A1(n5476) );
  nand02 U2344 ( .Y(n5477), .A0(n5468), .A1(n5478) );
  nand02 U2345 ( .Y(n5479), .A0(n5468), .A1(n5480) );
  nand02 U2346 ( .Y(n5481), .A0(n5468), .A1(n5482) );
  nand02 U2347 ( .Y(n5483), .A0(n5468), .A1(n5484) );
  nand02 U2348 ( .Y(n5485), .A0(n5463), .A1(n5464) );
  inv01 U2349 ( .Y(n5470), .A(n5485) );
  nand02 U2350 ( .Y(n5486), .A0(n5463), .A1(n5464) );
  inv01 U2351 ( .Y(n5472), .A(n5486) );
  nand02 U2352 ( .Y(n5487), .A0(n5463), .A1(n5465) );
  inv01 U2353 ( .Y(n5474), .A(n5487) );
  nand02 U2354 ( .Y(n5488), .A0(n5463), .A1(n5466) );
  inv01 U2355 ( .Y(n5476), .A(n5488) );
  nand02 U2356 ( .Y(n5489), .A0(n5464), .A1(n5465) );
  inv01 U2357 ( .Y(n5478), .A(n5489) );
  nand02 U2358 ( .Y(n5490), .A0(n5464), .A1(n5466) );
  inv01 U2359 ( .Y(n5480), .A(n5490) );
  nand02 U2360 ( .Y(n5491), .A0(n5465), .A1(n5467) );
  inv01 U2361 ( .Y(n5482), .A(n5491) );
  nand02 U2362 ( .Y(n5492), .A0(n5466), .A1(n5467) );
  inv01 U2363 ( .Y(n5484), .A(n5492) );
  nand02 U2364 ( .Y(n5493), .A0(n5469), .A1(n5471) );
  inv01 U2365 ( .Y(n5494), .A(n5493) );
  nand02 U2366 ( .Y(n5495), .A0(n5473), .A1(n5475) );
  inv01 U2367 ( .Y(n5496), .A(n5495) );
  nand02 U2368 ( .Y(n5497), .A0(n5494), .A1(n5496) );
  inv01 U2369 ( .Y(n5461), .A(n5497) );
  nand02 U2370 ( .Y(n5498), .A0(n5477), .A1(n5479) );
  inv01 U2371 ( .Y(n5499), .A(n5498) );
  nand02 U2372 ( .Y(n5500), .A0(n5481), .A1(n5483) );
  inv01 U2373 ( .Y(n5501), .A(n5500) );
  nand02 U2374 ( .Y(n5502), .A0(n5499), .A1(n5501) );
  inv01 U2375 ( .Y(n5462), .A(n5502) );
  ao221 U2376 ( .Y(n5503), .A0(n6298), .A1(n6299), .B0(n6086), .B1(n6300), 
        .C0(n6012) );
  inv01 U2377 ( .Y(n5504), .A(n5503) );
  ao221 U2378 ( .Y(n5505), .A0(n6159), .A1(n6160), .B0(n6088), .B1(n6161), 
        .C0(n6008) );
  inv01 U2379 ( .Y(n5506), .A(n5505) );
  inv01 U2380 ( .Y(n6268), .A(n5507) );
  inv01 U2381 ( .Y(n5508), .A(n6247) );
  inv01 U2382 ( .Y(n5509), .A(n6263) );
  inv01 U2383 ( .Y(n5510), .A(n6246) );
  inv01 U2384 ( .Y(n5511), .A(n4320) );
  nand02 U2385 ( .Y(n5507), .A0(n5512), .A1(n5513) );
  nand02 U2386 ( .Y(n5514), .A0(n5508), .A1(n5509) );
  inv01 U2387 ( .Y(n5512), .A(n5514) );
  nand02 U2388 ( .Y(n5515), .A0(n5510), .A1(n5511) );
  inv01 U2389 ( .Y(n5513), .A(n5515) );
  inv01 U2390 ( .Y(n6439), .A(n5516) );
  inv01 U2391 ( .Y(n5517), .A(n6392) );
  inv01 U2392 ( .Y(n5518), .A(n6390) );
  inv01 U2393 ( .Y(n5519), .A(n6391) );
  inv01 U2394 ( .Y(n5520), .A(n4362) );
  nand02 U2395 ( .Y(n5516), .A0(n5521), .A1(n5522) );
  nand02 U2396 ( .Y(n5523), .A0(n5517), .A1(n5518) );
  inv01 U2397 ( .Y(n5521), .A(n5523) );
  nand02 U2398 ( .Y(n5524), .A0(n5519), .A1(n5520) );
  inv01 U2399 ( .Y(n5522), .A(n5524) );
  inv01 U2400 ( .Y(dvdnd_50_o[41]), .A(n5525) );
  nor02 U2401 ( .Y(n5526), .A0(n6327), .A1(n6122) );
  nor02 U2402 ( .Y(n5527), .A0(n6357), .A1(n6358) );
  inv01 U2403 ( .Y(n5528), .A(n4374) );
  nor02 U2404 ( .Y(n5525), .A0(n5528), .A1(n5529) );
  nor02 U2405 ( .Y(n5530), .A0(n5526), .A1(n5527) );
  inv01 U2406 ( .Y(n5529), .A(n5530) );
  inv02 U2407 ( .Y(n6122), .A(n6119) );
  inv01 U2408 ( .Y(dvsor_27_o[13]), .A(n5531) );
  nor02 U2409 ( .Y(n5532), .A0(n6209), .A1(n6130) );
  nor02 U2410 ( .Y(n5533), .A0(n6148), .A1(n6134) );
  inv01 U2411 ( .Y(n5534), .A(n4413) );
  nor02 U2412 ( .Y(n5531), .A0(n5534), .A1(n5535) );
  nor02 U2413 ( .Y(n5536), .A0(n5532), .A1(n5533) );
  inv01 U2414 ( .Y(n5535), .A(n5536) );
  inv01 U2415 ( .Y(dvdnd_50_o[40]), .A(n5537) );
  nor02 U2416 ( .Y(n5538), .A0(n6360), .A1(n6132) );
  nor02 U2417 ( .Y(n5539), .A0(n6338), .A1(n6136) );
  inv01 U2418 ( .Y(n5540), .A(n4386) );
  nor02 U2419 ( .Y(n5537), .A0(n5540), .A1(n5541) );
  nor02 U2420 ( .Y(n5542), .A0(n5538), .A1(n5539) );
  inv01 U2421 ( .Y(n5541), .A(n5542) );
  inv01 U2422 ( .Y(dvdnd_50_o[39]), .A(n5543) );
  nor02 U2423 ( .Y(n5544), .A0(n6362), .A1(n6132) );
  nor02 U2424 ( .Y(n5545), .A0(n6344), .A1(n6136) );
  inv01 U2425 ( .Y(n5546), .A(n4388) );
  nor02 U2426 ( .Y(n5543), .A0(n5546), .A1(n5547) );
  nor02 U2427 ( .Y(n5548), .A0(n5544), .A1(n5545) );
  inv01 U2428 ( .Y(n5547), .A(n5548) );
  inv02 U2429 ( .Y(n6130), .A(n6127) );
  inv01 U2430 ( .Y(dvsor_27_o[14]), .A(n5549) );
  nor02 U2431 ( .Y(n5550), .A0(n6204), .A1(n6134) );
  nor02 U2432 ( .Y(n5551), .A0(n6176), .A1(n6126) );
  inv01 U2433 ( .Y(n5552), .A(n4415) );
  nor02 U2434 ( .Y(n5549), .A0(n5552), .A1(n5553) );
  nor02 U2435 ( .Y(n5554), .A0(n5550), .A1(n5551) );
  inv01 U2436 ( .Y(n5553), .A(n5554) );
  inv04 U2437 ( .Y(n6134), .A(n6133) );
  inv01 U2438 ( .Y(dvsor_27_o[15]), .A(n5555) );
  nor02 U2439 ( .Y(n5556), .A0(n6193), .A1(n6128) );
  nor02 U2440 ( .Y(n5557), .A0(n6156), .A1(n6220) );
  inv01 U2441 ( .Y(n5558), .A(n4384) );
  nor02 U2442 ( .Y(n5555), .A0(n5558), .A1(n5559) );
  nor02 U2443 ( .Y(n5560), .A0(n5556), .A1(n5557) );
  inv01 U2444 ( .Y(n5559), .A(n5560) );
  inv02 U2445 ( .Y(n6128), .A(n6127) );
  buf02 U2446 ( .Y(n5561), .A(n____return3540_1_) );
  buf02 U2447 ( .Y(n5562), .A(n____return3540_4_) );
  buf02 U2448 ( .Y(n5563), .A(n____return3540_3_) );
  buf02 U2449 ( .Y(n5564), .A(n____return3540_2_) );
  nor02 U2450 ( .Y(n5565), .A0(n6110), .A1(n6092) );
  inv02 U2451 ( .Y(n5566), .A(n5565) );
  buf02 U2452 ( .Y(n5567), .A(opa_i[11]) );
  inv01 U2453 ( .Y(n5568), .A(n5567) );
  inv01 U2454 ( .Y(dvdnd_50_o[43]), .A(n5569) );
  nor02 U2455 ( .Y(n5570), .A0(n6344), .A1(n6132) );
  nor02 U2456 ( .Y(n5571), .A0(n6343), .A1(n6136) );
  inv01 U2457 ( .Y(n5572), .A(n6345) );
  nor02 U2458 ( .Y(n5569), .A0(n5572), .A1(n5573) );
  nor02 U2459 ( .Y(n5574), .A0(n5570), .A1(n5571) );
  inv01 U2460 ( .Y(n5573), .A(n5574) );
  inv01 U2461 ( .Y(dvsor_27_o[19]), .A(n5575) );
  nor02 U2462 ( .Y(n5576), .A0(n6194), .A1(n6126) );
  nor02 U2463 ( .Y(n5577), .A0(n6193), .A1(n6134) );
  inv01 U2464 ( .Y(n5578), .A(n6195) );
  nor02 U2465 ( .Y(n5575), .A0(n5578), .A1(n5579) );
  nor02 U2466 ( .Y(n5580), .A0(n5576), .A1(n5577) );
  inv01 U2467 ( .Y(n5579), .A(n5580) );
  inv01 U2468 ( .Y(dvdnd_50_o[44]), .A(n5581) );
  nor02 U2469 ( .Y(n5582), .A0(n6338), .A1(n6132) );
  nor02 U2470 ( .Y(n5583), .A0(n6337), .A1(n6136) );
  inv01 U2471 ( .Y(n5584), .A(n6339) );
  nor02 U2472 ( .Y(n5581), .A0(n5584), .A1(n5585) );
  nor02 U2473 ( .Y(n5586), .A0(n5582), .A1(n5583) );
  inv01 U2474 ( .Y(n5585), .A(n5586) );
  inv04 U2475 ( .Y(n6132), .A(n6131) );
  inv01 U2476 ( .Y(dvsor_27_o[18]), .A(n5587) );
  nor02 U2477 ( .Y(n5588), .A0(n6204), .A1(n6126) );
  nor02 U2478 ( .Y(n5589), .A0(n6203), .A1(n6134) );
  inv01 U2479 ( .Y(n5590), .A(n6205) );
  nor02 U2480 ( .Y(n5587), .A0(n5590), .A1(n5591) );
  nor02 U2481 ( .Y(n5592), .A0(n5588), .A1(n5589) );
  inv01 U2482 ( .Y(n5591), .A(n5592) );
  inv01 U2483 ( .Y(dvsor_27_o[17]), .A(n5593) );
  nor02 U2484 ( .Y(n5594), .A0(n6209), .A1(n6134) );
  nor02 U2485 ( .Y(n5595), .A0(n6148), .A1(n6126) );
  inv01 U2486 ( .Y(n5596), .A(n6210) );
  nor02 U2487 ( .Y(n5593), .A0(n5596), .A1(n5597) );
  nor02 U2488 ( .Y(n5598), .A0(n5594), .A1(n5595) );
  inv01 U2489 ( .Y(n5597), .A(n5598) );
  inv01 U2490 ( .Y(dvdnd_50_o[45]), .A(n5599) );
  nor02 U2491 ( .Y(n5600), .A0(n6328), .A1(n6132) );
  nor02 U2492 ( .Y(n5601), .A0(n6327), .A1(n6136) );
  inv01 U2493 ( .Y(n5602), .A(n6329) );
  nor02 U2494 ( .Y(n5599), .A0(n5602), .A1(n5603) );
  nor02 U2495 ( .Y(n5604), .A0(n5600), .A1(n5601) );
  inv01 U2496 ( .Y(n5603), .A(n5604) );
  inv01 U2497 ( .Y(dvsor_27_o[16]), .A(n5605) );
  nor02 U2498 ( .Y(n5606), .A0(n6151), .A1(n6126) );
  nor02 U2499 ( .Y(n5607), .A0(n6215), .A1(n6134) );
  inv01 U2500 ( .Y(n5608), .A(n6216) );
  nor02 U2501 ( .Y(n5605), .A0(n5608), .A1(n5609) );
  nor02 U2502 ( .Y(n5610), .A0(n5606), .A1(n5607) );
  inv01 U2503 ( .Y(n5609), .A(n5610) );
  inv04 U2504 ( .Y(n6126), .A(n6125) );
  inv01 U2505 ( .Y(dvdnd_50_o[42]), .A(n5611) );
  nor02 U2506 ( .Y(n5612), .A0(n6350), .A1(n6132) );
  nor02 U2507 ( .Y(n5613), .A0(n6349), .A1(n6136) );
  inv01 U2508 ( .Y(n5614), .A(n6351) );
  nor02 U2509 ( .Y(n5611), .A0(n5614), .A1(n5615) );
  nor02 U2510 ( .Y(n5616), .A0(n5612), .A1(n5613) );
  inv01 U2511 ( .Y(n5615), .A(n5616) );
  nand02 U2512 ( .Y(n6431), .A0(n5617), .A1(n5618) );
  inv01 U2513 ( .Y(n5619), .A(n6421) );
  inv01 U2514 ( .Y(n5620), .A(opa_i[18]) );
  inv01 U2515 ( .Y(n5621), .A(n6011) );
  inv01 U2516 ( .Y(n5622), .A(n6012) );
  inv01 U2517 ( .Y(n5623), .A(n6432) );
  nand02 U2518 ( .Y(n5617), .A0(n5621), .A1(n5624) );
  nand02 U2519 ( .Y(n5618), .A0(n5622), .A1(n5623) );
  nand02 U2520 ( .Y(n5625), .A0(n5619), .A1(n5620) );
  inv01 U2521 ( .Y(n5624), .A(n5625) );
  inv01 U2522 ( .Y(n6460), .A(n5626) );
  inv01 U2523 ( .Y(n5627), .A(opb_i[23]) );
  inv01 U2524 ( .Y(n5628), .A(opb_i[24]) );
  inv01 U2525 ( .Y(n5629), .A(opb_i[25]) );
  inv01 U2526 ( .Y(n5630), .A(opb_i[26]) );
  nand02 U2527 ( .Y(n5626), .A0(n5631), .A1(n5632) );
  nand02 U2528 ( .Y(n5633), .A0(n5627), .A1(n5628) );
  inv01 U2529 ( .Y(n5631), .A(n5633) );
  nand02 U2530 ( .Y(n5634), .A0(n5629), .A1(n5630) );
  inv01 U2531 ( .Y(n5632), .A(n5634) );
  nand02 U2532 ( .Y(n6419), .A0(n5635), .A1(n5636) );
  inv01 U2533 ( .Y(n5637), .A(n6420) );
  inv01 U2534 ( .Y(n5638), .A(n6012) );
  inv01 U2535 ( .Y(n5639), .A(n6030) );
  inv01 U2536 ( .Y(n5640), .A(n6421) );
  inv01 U2537 ( .Y(n5641), .A(n6005) );
  nand02 U2538 ( .Y(n5635), .A0(n5639), .A1(n5642) );
  nand02 U2539 ( .Y(n5636), .A0(n5640), .A1(n5641) );
  nand02 U2540 ( .Y(n5643), .A0(n5637), .A1(n5638) );
  inv01 U2541 ( .Y(n5642), .A(n5643) );
  buf02 U2542 ( .Y(n6012), .A(n6301) );
  nand02 U2543 ( .Y(n6250), .A0(n5644), .A1(n5645) );
  inv01 U2544 ( .Y(n5646), .A(n6251) );
  inv01 U2545 ( .Y(n5647), .A(n6213) );
  inv01 U2546 ( .Y(n5648), .A(n6008) );
  inv01 U2547 ( .Y(n5649), .A(n6252) );
  nand02 U2548 ( .Y(n5644), .A0(n5647), .A1(n5650) );
  nand02 U2549 ( .Y(n5645), .A0(n5648), .A1(n5649) );
  nand02 U2550 ( .Y(n5651), .A0(n5646), .A1(n4366) );
  inv01 U2551 ( .Y(n5650), .A(n5651) );
  inv01 U2552 ( .Y(n6291), .A(n5652) );
  nor02 U2553 ( .Y(n5653), .A0(n6253), .A1(n5654) );
  nor02 U2554 ( .Y(n5655), .A0(n5931), .A1(n6251) );
  nor02 U2555 ( .Y(n5652), .A0(n5653), .A1(n5655) );
  nor02 U2556 ( .Y(n5656), .A0(n6200), .A1(n6008) );
  inv01 U2557 ( .Y(n5654), .A(n5656) );
  buf02 U2558 ( .Y(n6008), .A(n6162) );
  inv02 U2559 ( .Y(n6294), .A(n5657) );
  nand02 U2560 ( .Y(n5657), .A0(n6292), .A1(n5658) );
  nand02 U2561 ( .Y(n5659), .A0(n5931), .A1(n5025) );
  inv01 U2562 ( .Y(n5658), .A(n5659) );
  inv02 U2563 ( .Y(n6293), .A(n5660) );
  nand02 U2564 ( .Y(n5660), .A0(n4687), .A1(n5661) );
  nand02 U2565 ( .Y(n5662), .A0(n4936), .A1(n6051) );
  inv01 U2566 ( .Y(n5661), .A(n5662) );
  inv02 U2567 ( .Y(n6295), .A(n5663) );
  nand02 U2568 ( .Y(n5663), .A0(n5037), .A1(n5664) );
  nand02 U2569 ( .Y(n5665), .A0(n4934), .A1(n6046) );
  inv01 U2570 ( .Y(n5664), .A(n5665) );
  inv02 U2571 ( .Y(n6430), .A(n5666) );
  nand02 U2572 ( .Y(n5666), .A0(n6435), .A1(n5667) );
  nand02 U2573 ( .Y(n5668), .A0(n5568), .A1(n6074) );
  inv01 U2574 ( .Y(n5667), .A(n5668) );
  inv02 U2575 ( .Y(n6437), .A(n5669) );
  nand02 U2576 ( .Y(n5669), .A0(n6429), .A1(n5670) );
  nand02 U2577 ( .Y(n5671), .A0(n5682), .A1(n6076) );
  inv01 U2578 ( .Y(n5670), .A(n5671) );
  buf02 U2579 ( .Y(n5672), .A(opa_i[2]) );
  inv02 U2580 ( .Y(n5673), .A(n5672) );
  inv02 U2581 ( .Y(n6296), .A(n5674) );
  nand02 U2582 ( .Y(n5674), .A0(n4685), .A1(n5675) );
  nand02 U2583 ( .Y(n5676), .A0(n4992), .A1(n6057) );
  inv01 U2584 ( .Y(n5675), .A(n5676) );
  nor02 U2585 ( .Y(n5677), .A0(n6118), .A1(n6098) );
  inv02 U2586 ( .Y(n5678), .A(n5677) );
  nand02 U2587 ( .Y(n5679), .A0(opa_i[8]), .A1(n6444) );
  inv02 U2588 ( .Y(n5680), .A(n5679) );
  buf02 U2589 ( .Y(n5681), .A(opa_i[4]) );
  inv02 U2590 ( .Y(n5682), .A(n5681) );
  inv01 U2591 ( .Y(n6461), .A(n5683) );
  inv01 U2592 ( .Y(n5684), .A(opb_i[27]) );
  inv01 U2593 ( .Y(n5685), .A(opb_i[28]) );
  inv01 U2594 ( .Y(n5686), .A(opb_i[29]) );
  inv01 U2595 ( .Y(n5687), .A(opb_i[30]) );
  nand02 U2596 ( .Y(n5683), .A0(n5688), .A1(n5689) );
  nand02 U2597 ( .Y(n5690), .A0(n5684), .A1(n5685) );
  inv01 U2598 ( .Y(n5688), .A(n5690) );
  nand02 U2599 ( .Y(n5691), .A0(n5686), .A1(n5687) );
  inv01 U2600 ( .Y(n5689), .A(n5691) );
  buf02 U2601 ( .Y(n5692), .A(n____return3540_6_) );
  buf02 U2602 ( .Y(n5693), .A(n____return3540_5_) );
  xor2 U2603 ( .Y(n5694), .A0(s_expa_in_8_), .A1(n6445) );
  inv02 U2604 ( .Y(n5695), .A(n5694) );
  xor2 U2605 ( .Y(n5696), .A0(n5915), .A1(s_expa_in_7_) );
  inv02 U2606 ( .Y(n5697), .A(n5696) );
  inv01 U2607 ( .Y(n5698), .A(n6372) );
  inv01 U2608 ( .Y(n5699), .A(n5698) );
  inv01 U2609 ( .Y(n5700), .A(n5698) );
  inv01 U2610 ( .Y(n6464), .A(n5701) );
  inv01 U2611 ( .Y(n5702), .A(opa_i[27]) );
  inv01 U2612 ( .Y(n5703), .A(opa_i[28]) );
  inv01 U2613 ( .Y(n5704), .A(opa_i[29]) );
  inv01 U2614 ( .Y(n5705), .A(opa_i[30]) );
  nand02 U2615 ( .Y(n5701), .A0(n5706), .A1(n5707) );
  nand02 U2616 ( .Y(n5708), .A0(n5702), .A1(n5703) );
  inv01 U2617 ( .Y(n5706), .A(n5708) );
  nand02 U2618 ( .Y(n5709), .A0(n5704), .A1(n5705) );
  inv01 U2619 ( .Y(n5707), .A(n5709) );
  inv02 U2620 ( .Y(s_dvd_zeros_2_), .A(n5710) );
  inv01 U2621 ( .Y(n5711), .A(n6414) );
  inv01 U2622 ( .Y(n5712), .A(n6413) );
  inv01 U2623 ( .Y(n5713), .A(n6412) );
  inv01 U2624 ( .Y(n5714), .A(n4675) );
  nor02 U2625 ( .Y(n5710), .A0(n5715), .A1(n5716) );
  nor02 U2626 ( .Y(n5717), .A0(n5711), .A1(n5712) );
  inv01 U2627 ( .Y(n5715), .A(n5717) );
  nor02 U2628 ( .Y(n5718), .A0(n5713), .A1(n5714) );
  inv01 U2629 ( .Y(n5716), .A(n5718) );
  inv01 U2630 ( .Y(n6463), .A(n5719) );
  inv01 U2631 ( .Y(n5720), .A(opa_i[23]) );
  inv01 U2632 ( .Y(n5721), .A(opa_i[24]) );
  inv01 U2633 ( .Y(n5722), .A(opa_i[25]) );
  inv01 U2634 ( .Y(n5723), .A(opa_i[26]) );
  nand02 U2635 ( .Y(n5719), .A0(n5724), .A1(n5725) );
  nand02 U2636 ( .Y(n5726), .A0(n5720), .A1(n5721) );
  inv01 U2637 ( .Y(n5724), .A(n5726) );
  nand02 U2638 ( .Y(n5727), .A0(n5722), .A1(n5723) );
  inv01 U2639 ( .Y(n5725), .A(n5727) );
  xor2 U2640 ( .Y(n5728), .A0(n4855), .A1(n6465) );
  inv02 U2641 ( .Y(n5729), .A(n5728) );
  buf02 U2642 ( .Y(n6081), .A(s_div_zeros_3_) );
  buf02 U2643 ( .Y(n5730), .A(n6381) );
  nand02 U2644 ( .Y(n6185), .A0(n6225), .A1(n5731) );
  inv01 U2645 ( .Y(n5732), .A(n6139) );
  inv01 U2646 ( .Y(n5733), .A(n6046) );
  inv01 U2647 ( .Y(n5734), .A(n6138) );
  inv01 U2648 ( .Y(n5735), .A(n5157) );
  nand02 U2649 ( .Y(n5736), .A0(n5732), .A1(n5733) );
  nand02 U2650 ( .Y(n5737), .A0(n5734), .A1(n5735) );
  nand02 U2651 ( .Y(n5738), .A0(n5736), .A1(n5737) );
  inv01 U2652 ( .Y(n5731), .A(n5738) );
  nand02 U2653 ( .Y(n6192), .A0(n6231), .A1(n5739) );
  inv01 U2654 ( .Y(n5740), .A(n6139) );
  inv01 U2655 ( .Y(n5741), .A(n4934) );
  inv01 U2656 ( .Y(n5742), .A(n6138) );
  inv01 U2657 ( .Y(n5743), .A(n6051) );
  nand02 U2658 ( .Y(n5744), .A0(n5740), .A1(n5741) );
  nand02 U2659 ( .Y(n5745), .A0(n5742), .A1(n5743) );
  nand02 U2660 ( .Y(n5746), .A0(n5744), .A1(n5745) );
  inv01 U2661 ( .Y(n5739), .A(n5746) );
  inv02 U2662 ( .Y(n6209), .A(n6185) );
  inv02 U2663 ( .Y(n6215), .A(n6192) );
  inv02 U2664 ( .Y(n6326), .A(n5747) );
  nor02 U2665 ( .Y(n5748), .A0(n6074), .A1(n6143) );
  nor02 U2666 ( .Y(n5749), .A0(n5568), .A1(n6142) );
  inv01 U2667 ( .Y(n5750), .A(n6364) );
  nor02 U2668 ( .Y(n5747), .A0(n5750), .A1(n5751) );
  nor02 U2669 ( .Y(n5752), .A0(n5748), .A1(n5749) );
  inv01 U2670 ( .Y(n5751), .A(n5752) );
  inv02 U2671 ( .Y(n6349), .A(n6326) );
  inv02 U2672 ( .Y(n6161), .A(n5753) );
  nor02 U2673 ( .Y(n5754), .A0(n6059), .A1(n6139) );
  nor02 U2674 ( .Y(n5755), .A0(n4934), .A1(n6138) );
  inv01 U2675 ( .Y(n5756), .A(n6221) );
  nor02 U2676 ( .Y(n5753), .A0(n5756), .A1(n5757) );
  nor02 U2677 ( .Y(n5758), .A0(n5754), .A1(n5755) );
  inv01 U2678 ( .Y(n5757), .A(n5758) );
  inv02 U2679 ( .Y(n6193), .A(n6161) );
  inv02 U2680 ( .Y(n6300), .A(n5759) );
  nor02 U2681 ( .Y(n5760), .A0(n5928), .A1(n6143) );
  nor02 U2682 ( .Y(n5761), .A0(n6080), .A1(n6142) );
  inv01 U2683 ( .Y(n5762), .A(n6359) );
  nor02 U2684 ( .Y(n5759), .A0(n5762), .A1(n5763) );
  nor02 U2685 ( .Y(n5764), .A0(n5760), .A1(n5761) );
  inv01 U2686 ( .Y(n5763), .A(n5764) );
  inv02 U2687 ( .Y(n6346), .A(n5765) );
  nor02 U2688 ( .Y(n5766), .A0(n4361), .A1(n6142) );
  nor02 U2689 ( .Y(n5767), .A0(n6044), .A1(n6143) );
  nor02 U2690 ( .Y(n5765), .A0(n5766), .A1(n5767) );
  inv02 U2691 ( .Y(n6327), .A(n6300) );
  inv02 U2692 ( .Y(n6369), .A(n6346) );
  nand02 U2693 ( .Y(n6177), .A0(n6208), .A1(n5768) );
  inv01 U2694 ( .Y(n5769), .A(n6139) );
  inv01 U2695 ( .Y(n5770), .A(n4364) );
  inv01 U2696 ( .Y(n5771), .A(n6138) );
  inv01 U2697 ( .Y(n5772), .A(n6059) );
  nand02 U2698 ( .Y(n5773), .A0(n5769), .A1(n5770) );
  nand02 U2699 ( .Y(n5774), .A0(n5771), .A1(n5772) );
  nand02 U2700 ( .Y(n5775), .A0(n5773), .A1(n5774) );
  inv01 U2701 ( .Y(n5768), .A(n5775) );
  nand02 U2702 ( .Y(n6191), .A0(n6219), .A1(n5776) );
  inv01 U2703 ( .Y(n5777), .A(n6139) );
  inv01 U2704 ( .Y(n5778), .A(n5025) );
  inv01 U2705 ( .Y(n5779), .A(n6138) );
  inv01 U2706 ( .Y(n5780), .A(n6046) );
  nand02 U2707 ( .Y(n5781), .A0(n5777), .A1(n5778) );
  nand02 U2708 ( .Y(n5782), .A0(n5779), .A1(n5780) );
  nand02 U2709 ( .Y(n5783), .A0(n5781), .A1(n5782) );
  inv01 U2710 ( .Y(n5776), .A(n5783) );
  nand02 U2711 ( .Y(n6184), .A0(n6214), .A1(n5784) );
  inv01 U2712 ( .Y(n5785), .A(n6139) );
  inv01 U2713 ( .Y(n5786), .A(n6213) );
  inv01 U2714 ( .Y(n5787), .A(n6138) );
  inv01 U2715 ( .Y(n5788), .A(n6212) );
  nand02 U2716 ( .Y(n5789), .A0(n5785), .A1(n5786) );
  nand02 U2717 ( .Y(n5790), .A0(n5787), .A1(n5788) );
  nand02 U2718 ( .Y(n5791), .A0(n5789), .A1(n5790) );
  inv01 U2719 ( .Y(n5784), .A(n5791) );
  inv01 U2720 ( .Y(n6212), .A(opb_i[14]) );
  inv01 U2721 ( .Y(n6325), .A(n5792) );
  nor02 U2722 ( .Y(n5793), .A0(n5991), .A1(n6143) );
  nor02 U2723 ( .Y(n5794), .A0(n5929), .A1(n6142) );
  inv01 U2724 ( .Y(n5795), .A(n6356) );
  nor02 U2725 ( .Y(n5792), .A0(n5795), .A1(n5796) );
  nor02 U2726 ( .Y(n5797), .A0(n5793), .A1(n5794) );
  inv01 U2727 ( .Y(n5796), .A(n5797) );
  inv01 U2728 ( .Y(n6319), .A(n5798) );
  nor02 U2729 ( .Y(n5799), .A0(n6010), .A1(n6143) );
  nor02 U2730 ( .Y(n5800), .A0(n5991), .A1(n6142) );
  inv01 U2731 ( .Y(n5801), .A(n6348) );
  nor02 U2732 ( .Y(n5798), .A0(n5801), .A1(n5802) );
  nor02 U2733 ( .Y(n5803), .A0(n5799), .A1(n5800) );
  inv01 U2734 ( .Y(n5802), .A(n5803) );
  inv02 U2735 ( .Y(n6263), .A(n5804) );
  nand02 U2736 ( .Y(n5804), .A0(opb_i[0]), .A1(n5805) );
  nand02 U2737 ( .Y(n5806), .A0(n5161), .A1(n6229) );
  inv01 U2738 ( .Y(n5805), .A(n5806) );
  inv01 U2739 ( .Y(n6313), .A(n5807) );
  nor02 U2740 ( .Y(n5808), .A0(n6007), .A1(n6143) );
  nor02 U2741 ( .Y(n5809), .A0(n6011), .A1(n6142) );
  inv01 U2742 ( .Y(n5810), .A(n6342) );
  nor02 U2743 ( .Y(n5807), .A0(n5810), .A1(n5811) );
  nor02 U2744 ( .Y(n5812), .A0(n5808), .A1(n5809) );
  inv01 U2745 ( .Y(n5811), .A(n5812) );
  nand02 U2746 ( .Y(n6160), .A0(n6202), .A1(n5813) );
  inv01 U2747 ( .Y(n5814), .A(n6139) );
  inv01 U2748 ( .Y(n5815), .A(n6200) );
  inv01 U2749 ( .Y(n5816), .A(n6138) );
  inv01 U2750 ( .Y(n5817), .A(n5025) );
  nand02 U2751 ( .Y(n5818), .A0(n5814), .A1(n5815) );
  nand02 U2752 ( .Y(n5819), .A0(n5816), .A1(n5817) );
  nand02 U2753 ( .Y(n5820), .A0(n5818), .A1(n5819) );
  inv01 U2754 ( .Y(n5813), .A(n5820) );
  nand02 U2755 ( .Y(n6299), .A0(n6336), .A1(n5821) );
  inv01 U2756 ( .Y(n5822), .A(n6143) );
  inv01 U2757 ( .Y(n5823), .A(n5077) );
  inv01 U2758 ( .Y(n5824), .A(n6142) );
  inv01 U2759 ( .Y(n5825), .A(n6007) );
  nand02 U2760 ( .Y(n5826), .A0(n5822), .A1(n5823) );
  nand02 U2761 ( .Y(n5827), .A0(n5824), .A1(n5825) );
  nand02 U2762 ( .Y(n5828), .A0(n5826), .A1(n5827) );
  inv01 U2763 ( .Y(n5821), .A(n5828) );
  inv02 U2764 ( .Y(n6246), .A(n5829) );
  nand02 U2765 ( .Y(n5829), .A0(opb_i[8]), .A1(n5830) );
  nand02 U2766 ( .Y(n5831), .A0(n4687), .A1(n6051) );
  inv01 U2767 ( .Y(n5830), .A(n5831) );
  inv02 U2768 ( .Y(n6175), .A(n5832) );
  nor02 U2769 ( .Y(n5833), .A0(n5157), .A1(n6139) );
  nor02 U2770 ( .Y(n5834), .A0(n6049), .A1(n6138) );
  inv01 U2771 ( .Y(n5835), .A(n6237) );
  nor02 U2772 ( .Y(n5832), .A0(n5835), .A1(n5836) );
  nor02 U2773 ( .Y(n5837), .A0(n5833), .A1(n5834) );
  inv01 U2774 ( .Y(n5836), .A(n5837) );
  nand02 U2775 ( .Y(n6190), .A0(n6228), .A1(n5838) );
  inv01 U2776 ( .Y(n5839), .A(n6139) );
  inv01 U2777 ( .Y(n5840), .A(n4936) );
  inv01 U2778 ( .Y(n5841), .A(n6138) );
  inv01 U2779 ( .Y(n5842), .A(n6057) );
  nand02 U2780 ( .Y(n5843), .A0(n5839), .A1(n5840) );
  nand02 U2781 ( .Y(n5844), .A0(n5841), .A1(n5842) );
  nand02 U2782 ( .Y(n5845), .A0(n5843), .A1(n5844) );
  inv01 U2783 ( .Y(n5838), .A(n5845) );
  nand02 U2784 ( .Y(n6182), .A0(n6227), .A1(n5846) );
  inv01 U2785 ( .Y(n5847), .A(n6139) );
  inv01 U2786 ( .Y(n5848), .A(n6051) );
  inv01 U2787 ( .Y(n5849), .A(n6138) );
  inv01 U2788 ( .Y(n5850), .A(n6226) );
  nand02 U2789 ( .Y(n5851), .A0(n5847), .A1(n5848) );
  nand02 U2790 ( .Y(n5852), .A0(n5849), .A1(n5850) );
  nand02 U2791 ( .Y(n5853), .A0(n5851), .A1(n5852) );
  inv01 U2792 ( .Y(n5846), .A(n5853) );
  inv01 U2793 ( .Y(n6226), .A(opb_i[6]) );
  inv02 U2794 ( .Y(n6311), .A(n5854) );
  nor02 U2795 ( .Y(n5855), .A0(n6070), .A1(n6143) );
  nor02 U2796 ( .Y(n5856), .A0(n5959), .A1(n6142) );
  inv01 U2797 ( .Y(n5857), .A(n6368) );
  nor02 U2798 ( .Y(n5854), .A0(n5857), .A1(n5858) );
  nor02 U2799 ( .Y(n5859), .A0(n5855), .A1(n5856) );
  inv01 U2800 ( .Y(n5858), .A(n5859) );
  inv02 U2801 ( .Y(n6317), .A(n5860) );
  nor02 U2802 ( .Y(n5861), .A0(n5959), .A1(n6143) );
  nor02 U2803 ( .Y(n5862), .A0(n6370), .A1(n6142) );
  inv01 U2804 ( .Y(n5863), .A(n6371) );
  nor02 U2805 ( .Y(n5860), .A0(n5863), .A1(n5864) );
  nor02 U2806 ( .Y(n5865), .A0(n5861), .A1(n5862) );
  inv01 U2807 ( .Y(n5864), .A(n5865) );
  inv02 U2808 ( .Y(n6324), .A(n5866) );
  nor02 U2809 ( .Y(n5867), .A0(n6370), .A1(n6143) );
  nor02 U2810 ( .Y(n5868), .A0(n6072), .A1(n6142) );
  inv01 U2811 ( .Y(n5869), .A(n6374) );
  nor02 U2812 ( .Y(n5866), .A0(n5869), .A1(n5870) );
  nor02 U2813 ( .Y(n5871), .A0(n5867), .A1(n5868) );
  inv01 U2814 ( .Y(n5870), .A(n5871) );
  inv02 U2815 ( .Y(n6391), .A(n5872) );
  nand02 U2816 ( .Y(n5872), .A0(opa_i[0]), .A1(n5873) );
  nand02 U2817 ( .Y(n5874), .A0(n5159), .A1(n6044) );
  inv01 U2818 ( .Y(n5873), .A(n5874) );
  inv02 U2819 ( .Y(n6341), .A(n5875) );
  nor02 U2820 ( .Y(n5876), .A0(n5029), .A1(n6143) );
  nor02 U2821 ( .Y(n5877), .A0(n6076), .A1(n6142) );
  inv01 U2822 ( .Y(n5878), .A(n6377) );
  nor02 U2823 ( .Y(n5875), .A0(n5878), .A1(n5879) );
  nor02 U2824 ( .Y(n5880), .A0(n5876), .A1(n5877) );
  inv01 U2825 ( .Y(n5879), .A(n5880) );
  inv02 U2826 ( .Y(n6197), .A(n5881) );
  nor02 U2827 ( .Y(n5882), .A0(n6053), .A1(n6139) );
  nor02 U2828 ( .Y(n5883), .A0(n6233), .A1(n6138) );
  inv01 U2829 ( .Y(n5884), .A(n6234) );
  nor02 U2830 ( .Y(n5881), .A0(n5884), .A1(n5885) );
  nor02 U2831 ( .Y(n5886), .A0(n5882), .A1(n5883) );
  inv01 U2832 ( .Y(n5885), .A(n5886) );
  inv02 U2833 ( .Y(n6207), .A(n5887) );
  nor02 U2834 ( .Y(n5888), .A0(n6226), .A1(n6139) );
  nor02 U2835 ( .Y(n5889), .A0(n6053), .A1(n6138) );
  inv01 U2836 ( .Y(n5890), .A(n6236) );
  nor02 U2837 ( .Y(n5887), .A0(n5890), .A1(n5891) );
  nor02 U2838 ( .Y(n5892), .A0(n5888), .A1(n5889) );
  inv01 U2839 ( .Y(n5891), .A(n5892) );
  buf08 U2840 ( .Y(n6139), .A(n6201) );
  nand02 U2841 ( .Y(n6331), .A0(n6380), .A1(n5893) );
  inv01 U2842 ( .Y(n5894), .A(n6143) );
  inv01 U2843 ( .Y(n5895), .A(n6078) );
  inv01 U2844 ( .Y(n5896), .A(n6142) );
  inv01 U2845 ( .Y(n5897), .A(n5673) );
  nand02 U2846 ( .Y(n5898), .A0(n5894), .A1(n5895) );
  nand02 U2847 ( .Y(n5899), .A0(n5896), .A1(n5897) );
  nand02 U2848 ( .Y(n5900), .A0(n5898), .A1(n5899) );
  inv01 U2849 ( .Y(n5893), .A(n5900) );
  nand02 U2850 ( .Y(n6347), .A0(n6378), .A1(n5901) );
  inv01 U2851 ( .Y(n5902), .A(n6143) );
  inv01 U2852 ( .Y(n5903), .A(n6076) );
  inv01 U2853 ( .Y(n5904), .A(n6142) );
  inv01 U2854 ( .Y(n5905), .A(n5682) );
  nand02 U2855 ( .Y(n5906), .A0(n5902), .A1(n5903) );
  nand02 U2856 ( .Y(n5907), .A0(n5904), .A1(n5905) );
  nand02 U2857 ( .Y(n5908), .A0(n5906), .A1(n5907) );
  inv01 U2858 ( .Y(n5901), .A(n5908) );
  buf08 U2859 ( .Y(n6142), .A(n6334) );
  buf08 U2860 ( .Y(n6143), .A(n6335) );
  inv02 U2861 ( .Y(n6330), .A(n5909) );
  nand02 U2862 ( .Y(n5909), .A0(n6302), .A1(n5910) );
  nand02 U2863 ( .Y(n5911), .A0(n6354), .A1(n6113) );
  inv01 U2864 ( .Y(n5910), .A(n5911) );
  buf02 U2865 ( .Y(n5912), .A(n6196) );
  inv02 U2866 ( .Y(n6302), .A(n6355) );
  inv02 U2867 ( .Y(n6176), .A(n6207) );
  inv02 U2868 ( .Y(n6360), .A(n6341) );
  ao22 U2869 ( .Y(n5913), .A0(n6217), .A1(n6111), .B0(n6152), .B1(n6167) );
  inv02 U2870 ( .Y(n5914), .A(n5913) );
  buf02 U2871 ( .Y(n5915), .A(n6448) );
  buf02 U2872 ( .Y(n5916), .A(n6448) );
  inv02 U2873 ( .Y(n6370), .A(opa_i[8]) );
  ao22 U2874 ( .Y(n5917), .A0(n6352), .A1(s_dvd_zeros_2_), .B0(n6353), .B1(
        n6354) );
  inv02 U2875 ( .Y(n5918), .A(n5917) );
  inv02 U2876 ( .Y(s_dvd_zeros_0_), .A(n5919) );
  inv01 U2877 ( .Y(n5920), .A(n6439) );
  inv01 U2878 ( .Y(n5921), .A(n4677) );
  inv01 U2879 ( .Y(n5922), .A(n6438) );
  nor02 U2880 ( .Y(n5919), .A0(n5922), .A1(n5923) );
  nor02 U2881 ( .Y(n5924), .A0(n5920), .A1(n5921) );
  inv01 U2882 ( .Y(n5923), .A(n5924) );
  or02 U2883 ( .Y(n5925), .A0(n6382), .A1(s_dvd_zeros_1_) );
  inv02 U2884 ( .Y(n5926), .A(n5925) );
  buf02 U2885 ( .Y(n5927), .A(opa_i[15]) );
  inv02 U2886 ( .Y(n5929), .A(n5927) );
  or02 U2887 ( .Y(n5930), .A0(opb_i[18]), .A1(opb_i[17]) );
  inv02 U2888 ( .Y(n5931), .A(n5930) );
  nand02 U2889 ( .Y(n6152), .A0(n6230), .A1(n5932) );
  inv01 U2890 ( .Y(n5933), .A(n6139) );
  inv01 U2891 ( .Y(n5934), .A(n4992) );
  inv01 U2892 ( .Y(n5935), .A(n6138) );
  inv01 U2893 ( .Y(n5936), .A(n6229) );
  nand02 U2894 ( .Y(n5937), .A0(n5933), .A1(n5934) );
  nand02 U2895 ( .Y(n5938), .A0(n5935), .A1(n5936) );
  nand02 U2896 ( .Y(n5939), .A0(n5937), .A1(n5938) );
  inv01 U2897 ( .Y(n5932), .A(n5939) );
  inv02 U2898 ( .Y(n6229), .A(opb_i[1]) );
  inv02 U2899 ( .Y(n6178), .A(n5940) );
  nor02 U2900 ( .Y(n5941), .A0(n6212), .A1(n6139) );
  nor02 U2901 ( .Y(n5942), .A0(n6055), .A1(n6138) );
  inv01 U2902 ( .Y(n5943), .A(n6222) );
  nor02 U2903 ( .Y(n5940), .A0(n5943), .A1(n5944) );
  nor02 U2904 ( .Y(n5945), .A0(n5941), .A1(n5942) );
  inv01 U2905 ( .Y(n5944), .A(n5945) );
  inv02 U2906 ( .Y(n6165), .A(n5946) );
  nor02 U2907 ( .Y(n5947), .A0(n6055), .A1(n6139) );
  nor02 U2908 ( .Y(n5948), .A0(n4936), .A1(n6138) );
  inv01 U2909 ( .Y(n5949), .A(n6232) );
  nor02 U2910 ( .Y(n5946), .A0(n5949), .A1(n5950) );
  nor02 U2911 ( .Y(n5951), .A0(n5947), .A1(n5948) );
  inv01 U2912 ( .Y(n5950), .A(n5951) );
  inv02 U2913 ( .Y(n6194), .A(n6165) );
  buf08 U2914 ( .Y(n6138), .A(n6188) );
  inv02 U2915 ( .Y(n6304), .A(n5952) );
  nor02 U2916 ( .Y(n5953), .A0(n5568), .A1(n6143) );
  nor02 U2917 ( .Y(n5954), .A0(n6070), .A1(n6142) );
  inv01 U2918 ( .Y(n5955), .A(n6366) );
  nor02 U2919 ( .Y(n5952), .A0(n5955), .A1(n5956) );
  nor02 U2920 ( .Y(n5957), .A0(n5953), .A1(n5954) );
  inv01 U2921 ( .Y(n5956), .A(n5957) );
  buf02 U2922 ( .Y(n5958), .A(opa_i[9]) );
  inv02 U2923 ( .Y(n5959), .A(n5958) );
  inv02 U2924 ( .Y(n6353), .A(n5960) );
  nor02 U2925 ( .Y(n5961), .A0(n5682), .A1(n6143) );
  nor02 U2926 ( .Y(n5962), .A0(n6078), .A1(n6142) );
  inv01 U2927 ( .Y(n5963), .A(n6379) );
  nor02 U2928 ( .Y(n5960), .A0(n5963), .A1(n5964) );
  nor02 U2929 ( .Y(n5965), .A0(n5961), .A1(n5962) );
  inv01 U2930 ( .Y(n5964), .A(n5965) );
  inv02 U2931 ( .Y(n6328), .A(n6304) );
  inv02 U2932 ( .Y(n6320), .A(n5966) );
  nor02 U2933 ( .Y(n5967), .A0(n5027), .A1(n6143) );
  nor02 U2934 ( .Y(n5968), .A0(n6074), .A1(n6142) );
  inv01 U2935 ( .Y(n5969), .A(n6363) );
  nor02 U2936 ( .Y(n5966), .A0(n5969), .A1(n5970) );
  nor02 U2937 ( .Y(n5971), .A0(n5967), .A1(n5968) );
  inv01 U2938 ( .Y(n5970), .A(n5971) );
  inv02 U2939 ( .Y(n6340), .A(n5972) );
  nor02 U2940 ( .Y(n5973), .A0(n5673), .A1(n6143) );
  nor02 U2941 ( .Y(n5974), .A0(n4361), .A1(n5730) );
  nor02 U2942 ( .Y(n5975), .A0(n6044), .A1(n6142) );
  nor02 U2943 ( .Y(n5972), .A0(n5975), .A1(n5976) );
  nor02 U2944 ( .Y(n5977), .A0(n5973), .A1(n5974) );
  inv01 U2945 ( .Y(n5976), .A(n5977) );
  inv02 U2946 ( .Y(n6314), .A(n5978) );
  nor02 U2947 ( .Y(n5979), .A0(n6080), .A1(n6143) );
  nor02 U2948 ( .Y(n5980), .A0(n5027), .A1(n6142) );
  inv01 U2949 ( .Y(n5981), .A(n6361) );
  nor02 U2950 ( .Y(n5978), .A0(n5981), .A1(n5982) );
  nor02 U2951 ( .Y(n5983), .A0(n5979), .A1(n5980) );
  inv01 U2952 ( .Y(n5982), .A(n5983) );
  inv02 U2953 ( .Y(n6367), .A(n6340) );
  inv02 U2954 ( .Y(n6198), .A(n5984) );
  nor02 U2955 ( .Y(n5985), .A0(n6049), .A1(n6139) );
  nor02 U2956 ( .Y(n5986), .A0(n4992), .A1(n6138) );
  inv01 U2957 ( .Y(n5987), .A(n6235) );
  nor02 U2958 ( .Y(n5984), .A0(n5987), .A1(n5988) );
  nor02 U2959 ( .Y(n5989), .A0(n5985), .A1(n5986) );
  inv01 U2960 ( .Y(n5988), .A(n5989) );
  buf02 U2961 ( .Y(n5990), .A(opa_i[16]) );
  inv02 U2962 ( .Y(n5991), .A(n5990) );
  inv02 U2963 ( .Y(n6166), .A(n6198) );
  inv02 U2964 ( .Y(n6183), .A(n5992) );
  nor02 U2965 ( .Y(n5993), .A0(n6057), .A1(n6139) );
  nor02 U2966 ( .Y(n5994), .A0(n6223), .A1(n6138) );
  inv01 U2967 ( .Y(n5995), .A(n6224) );
  nor02 U2968 ( .Y(n5992), .A0(n5995), .A1(n5996) );
  nor02 U2969 ( .Y(n5997), .A0(n5993), .A1(n5994) );
  inv01 U2970 ( .Y(n5996), .A(n5997) );
  inv02 U2971 ( .Y(n6147), .A(n6183) );
  inv02 U2972 ( .Y(n6148), .A(n6182) );
  inv02 U2973 ( .Y(n6332), .A(n5998) );
  nor02 U2974 ( .Y(n5999), .A0(n6072), .A1(n6143) );
  nor02 U2975 ( .Y(n6000), .A0(n5029), .A1(n6142) );
  inv01 U2976 ( .Y(n6001), .A(n6375) );
  nor02 U2977 ( .Y(n5998), .A0(n6001), .A1(n6002) );
  nor02 U2978 ( .Y(n6003), .A0(n5999), .A1(n6000) );
  inv01 U2979 ( .Y(n6002), .A(n6003) );
  inv02 U2980 ( .Y(n6365), .A(n6332) );
  inv02 U2981 ( .Y(n6204), .A(n6175) );
  inv02 U2982 ( .Y(n6338), .A(n6311) );
  inv02 U2983 ( .Y(n6344), .A(n6317) );
  inv02 U2984 ( .Y(n6350), .A(n6324) );
  or02 U2985 ( .Y(n6004), .A0(opa_i[18]), .A1(opa_i[17]) );
  inv02 U2986 ( .Y(n6005), .A(n6004) );
  buf02 U2987 ( .Y(n6006), .A(opa_i[18]) );
  inv02 U2988 ( .Y(n6007), .A(n6006) );
  inv02 U2989 ( .Y(n6151), .A(n6190) );
  buf02 U2990 ( .Y(n6009), .A(opa_i[17]) );
  inv01 U2991 ( .Y(n6010), .A(n6009) );
  inv02 U2992 ( .Y(n6011), .A(n6009) );
  inv02 U2993 ( .Y(n6357), .A(n6331) );
  inv04 U2994 ( .Y(n6163), .A(n6218) );
  inv02 U2995 ( .Y(n6292), .A(n6013) );
  inv01 U2996 ( .Y(n6014), .A(n6253) );
  inv01 U2997 ( .Y(n6015), .A(opb_i[19]) );
  inv01 U2998 ( .Y(n6016), .A(n6008) );
  nand02 U2999 ( .Y(n6013), .A0(n6016), .A1(n6017) );
  nand02 U3000 ( .Y(n6018), .A0(n6014), .A1(n6015) );
  inv01 U3001 ( .Y(n6017), .A(n6018) );
  inv02 U3002 ( .Y(n6251), .A(n6292) );
  inv02 U3003 ( .Y(n6156), .A(n6197) );
  inv02 U3004 ( .Y(s_div_zeros_0_), .A(n6019) );
  inv01 U3005 ( .Y(n6020), .A(n6268) );
  inv01 U3006 ( .Y(n6021), .A(n4625) );
  inv01 U3007 ( .Y(n6022), .A(n4623) );
  nor02 U3008 ( .Y(n6019), .A0(n6022), .A1(n6023) );
  nor02 U3009 ( .Y(n6024), .A0(n6020), .A1(n6021) );
  inv01 U3010 ( .Y(n6023), .A(n6024) );
  ao22 U3011 ( .Y(n6025), .A0(opb_i[1]), .A1(n6173), .B0(opb_i[0]), .B1(n6141)
         );
  inv01 U3012 ( .Y(n6026), .A(n6025) );
  inv02 U3013 ( .Y(n6027), .A(n6025) );
  inv02 U3014 ( .Y(n6441), .A(n6028) );
  inv01 U3015 ( .Y(n6029), .A(n6420) );
  inv01 U3016 ( .Y(n6031), .A(n6012) );
  nand02 U3017 ( .Y(n6028), .A0(n6031), .A1(n6032) );
  nand02 U3018 ( .Y(n6033), .A0(n6029), .A1(n6030) );
  inv01 U3019 ( .Y(n6032), .A(n6033) );
  inv02 U3020 ( .Y(n6421), .A(n6441) );
  inv02 U3021 ( .Y(s_dvd_zeros_3_), .A(n6034) );
  inv01 U3022 ( .Y(n6035), .A(n6407) );
  inv01 U3023 ( .Y(n6036), .A(n6406) );
  inv01 U3024 ( .Y(n6037), .A(n4689) );
  inv01 U3025 ( .Y(n6038), .A(n6405) );
  nor02 U3026 ( .Y(n6034), .A0(n6039), .A1(n6040) );
  nor02 U3027 ( .Y(n6041), .A0(n6035), .A1(n6036) );
  inv01 U3028 ( .Y(n6039), .A(n6041) );
  nor02 U3029 ( .Y(n6042), .A0(n6037), .A1(n6038) );
  inv01 U3030 ( .Y(n6040), .A(n6042) );
  buf02 U3031 ( .Y(n6043), .A(opa_i[1]) );
  inv02 U3032 ( .Y(n6044), .A(n6043) );
  buf02 U3033 ( .Y(n6045), .A(opb_i[13]) );
  inv02 U3034 ( .Y(n6046), .A(n6045) );
  inv02 U3035 ( .Y(n6047), .A(n6238) );
  inv02 U3036 ( .Y(n6238), .A(s_div_zeros_1_) );
  buf02 U3037 ( .Y(n6048), .A(opb_i[7]) );
  inv02 U3038 ( .Y(n6049), .A(n6048) );
  buf02 U3039 ( .Y(n6050), .A(opb_i[9]) );
  inv02 U3040 ( .Y(n6051), .A(n6050) );
  buf02 U3041 ( .Y(n6052), .A(opb_i[3]) );
  inv02 U3042 ( .Y(n6053), .A(n6052) );
  buf02 U3043 ( .Y(n6054), .A(opb_i[11]) );
  inv02 U3044 ( .Y(n6055), .A(n6054) );
  buf02 U3045 ( .Y(n6056), .A(opb_i[5]) );
  inv02 U3046 ( .Y(n6057), .A(n6056) );
  buf02 U3047 ( .Y(n6058), .A(opb_i[15]) );
  inv02 U3048 ( .Y(n6059), .A(n6058) );
  inv02 U3049 ( .Y(s_dvd_zeros_1_), .A(n6060) );
  inv01 U3050 ( .Y(n6061), .A(n6425) );
  inv01 U3051 ( .Y(n6062), .A(n6424) );
  inv01 U3052 ( .Y(n6063), .A(n6423) );
  inv01 U3053 ( .Y(n6064), .A(n6422) );
  nor02 U3054 ( .Y(n6060), .A0(n6065), .A1(n6066) );
  nor02 U3055 ( .Y(n6067), .A0(n6061), .A1(n6062) );
  inv01 U3056 ( .Y(n6065), .A(n6067) );
  nor02 U3057 ( .Y(n6068), .A0(n6063), .A1(n6064) );
  inv01 U3058 ( .Y(n6066), .A(n6068) );
  buf02 U3059 ( .Y(n6069), .A(opa_i[10]) );
  inv02 U3060 ( .Y(n6070), .A(n6069) );
  buf02 U3061 ( .Y(n6071), .A(opa_i[7]) );
  inv02 U3062 ( .Y(n6072), .A(n6071) );
  buf02 U3063 ( .Y(n6073), .A(opa_i[12]) );
  inv02 U3064 ( .Y(n6074), .A(n6073) );
  buf02 U3065 ( .Y(n6075), .A(opa_i[5]) );
  inv02 U3066 ( .Y(n6076), .A(n6075) );
  buf02 U3067 ( .Y(n6077), .A(opa_i[3]) );
  inv02 U3068 ( .Y(n6078), .A(n6077) );
  buf02 U3069 ( .Y(n6079), .A(opa_i[14]) );
  inv02 U3070 ( .Y(n6080), .A(n6079) );
  or02 U3071 ( .Y(n6082), .A0(s_dvd_zeros_0_), .A1(s_dvd_zeros_1_) );
  inv02 U3072 ( .Y(n6083), .A(n6082) );
  buf02 U3073 ( .Y(n6084), .A(n6157) );
  inv02 U3074 ( .Y(n6092), .A(s_dvd_zeros_3_) );
  inv02 U3075 ( .Y(n6113), .A(s_dvd_zeros_3_) );
  or02 U3076 ( .Y(n6085), .A0(n5566), .A1(n6089) );
  inv02 U3077 ( .Y(n6086), .A(n6085) );
  inv02 U3078 ( .Y(n6098), .A(n6081) );
  inv02 U3079 ( .Y(n6103), .A(n6081) );
  or02 U3080 ( .Y(n6087), .A0(n5678), .A1(n6111) );
  inv02 U3081 ( .Y(n6088), .A(n6087) );
  inv02 U3082 ( .Y(n6089), .A(n6354) );
  inv02 U3083 ( .Y(n6298), .A(n6090) );
  inv01 U3084 ( .Y(n6091), .A(n6109) );
  inv01 U3085 ( .Y(n6093), .A(n6354) );
  nand02 U3086 ( .Y(n6090), .A0(n6093), .A1(n6094) );
  nand02 U3087 ( .Y(n6095), .A0(n6091), .A1(n6092) );
  inv01 U3088 ( .Y(n6094), .A(n6095) );
  inv04 U3089 ( .Y(n6354), .A(s_dvd_zeros_2_) );
  inv02 U3090 ( .Y(n6109), .A(n6108) );
  inv02 U3091 ( .Y(n6159), .A(n6096) );
  inv01 U3092 ( .Y(n6097), .A(n6118) );
  inv01 U3093 ( .Y(n6099), .A(n6167) );
  nand02 U3094 ( .Y(n6096), .A0(n6099), .A1(n6100) );
  nand02 U3095 ( .Y(n6101), .A0(n6097), .A1(n6098) );
  inv01 U3096 ( .Y(n6100), .A(n6101) );
  inv02 U3097 ( .Y(n6167), .A(n6111) );
  inv01 U3098 ( .Y(n6104), .A(n6111) );
  inv01 U3099 ( .Y(n6105), .A(n6118) );
  nand02 U3100 ( .Y(n6102), .A0(n6105), .A1(n6106) );
  nand02 U3101 ( .Y(n6107), .A0(n6103), .A1(n6104) );
  inv01 U3102 ( .Y(n6106), .A(n6107) );
  inv02 U3103 ( .Y(n6108), .A(n4400) );
  inv02 U3104 ( .Y(n6110), .A(n6108) );
  buf12 U3105 ( .Y(n6111), .A(n4391) );
  inv01 U3106 ( .Y(n6114), .A(n6089) );
  inv01 U3107 ( .Y(n6115), .A(n6110) );
  nand02 U3108 ( .Y(n6112), .A0(n6115), .A1(n6116) );
  nand02 U3109 ( .Y(n6117), .A0(n6113), .A1(n6114) );
  inv01 U3110 ( .Y(n6116), .A(n6117) );
  buf12 U3111 ( .Y(n6118), .A(n4409) );
  buf02 U3112 ( .Y(n6119), .A(n6333) );
  inv02 U3113 ( .Y(n6121), .A(n6119) );
  inv04 U3114 ( .Y(n6123), .A(n4435) );
  inv04 U3115 ( .Y(n6124), .A(n4433) );
  buf02 U3116 ( .Y(n6125), .A(n6088) );
  buf02 U3117 ( .Y(n6127), .A(n6199) );
  inv02 U3118 ( .Y(n6129), .A(n6127) );
  buf02 U3119 ( .Y(n6131), .A(n6086) );
  buf02 U3120 ( .Y(n6133), .A(n6159) );
  buf02 U3121 ( .Y(n6135), .A(n6298) );
  buf08 U3122 ( .Y(n6137), .A(n6308) );
  inv08 U3123 ( .Y(n6309), .A(n5730) );
  and03 U3124 ( .Y(n6425), .A0(n6427), .A1(n6428), .A2(n6426) );
  nor02 U3125 ( .Y(n6428), .A0(n6411), .A1(n6383) );
  nor02 U3126 ( .Y(n6427), .A0(n5680), .A1(n6386) );
  inv01 U3127 ( .Y(n6426), .A(n6388) );
  nor02 U3128 ( .Y(n6424), .A0(n6395), .A1(n6431) );
  inv01 U3129 ( .Y(n6423), .A(n6397) );
  nor02 U3130 ( .Y(n6422), .A0(n6392), .A1(n6391) );
  inv01 U3131 ( .Y(n6418), .A(n6411) );
  inv01 U3132 ( .Y(n6417), .A(n6390) );
  inv01 U3133 ( .Y(n6416), .A(n5680) );
  inv01 U3134 ( .Y(n6415), .A(n6389) );
  inv01 U3135 ( .Y(n6413), .A(n6419) );
  nor02 U3136 ( .Y(n6412), .A0(n6396), .A1(n6397) );
  and03 U3137 ( .Y(n6407), .A0(n6409), .A1(n6410), .A2(n6408) );
  inv01 U3138 ( .Y(n6410), .A(n6411) );
  nor02 U3139 ( .Y(n6409), .A0(n6385), .A1(n6386) );
  inv01 U3140 ( .Y(n6408), .A(n5680) );
  inv01 U3141 ( .Y(n6406), .A(n6390) );
  inv01 U3142 ( .Y(n6405), .A(n6396) );
  and03 U3143 ( .Y(n6401), .A0(n6403), .A1(n4938), .A2(n6402) );
  inv01 U3144 ( .Y(n6403), .A(n6387) );
  nor02 U3145 ( .Y(n6402), .A0(n6388), .A1(n6389) );
  inv01 U3146 ( .Y(n6400), .A(n6391) );
  inv01 U3147 ( .Y(n6399), .A(n6394) );
  inv01 U3148 ( .Y(n6398), .A(n6397) );
  nand03 U3150 ( .Y(s_div_zeros_1_), .A0(n6241), .A1(n6242), .A2(n6240) );
  and03 U3151 ( .Y(n6242), .A0(n6244), .A1(n6245), .A2(n6243) );
  nor02 U3152 ( .Y(n6245), .A0(n6246), .A1(n6248) );
  or02 U3153 ( .Y(n6248), .A0(n6250), .A1(n6249) );
  inv01 U3154 ( .Y(n6244), .A(n6255) );
  nor02 U3155 ( .Y(n6243), .A0(n6257), .A1(n6258) );
  nor02 U3156 ( .Y(n6241), .A0(n4359), .A1(n6262) );
  nor02 U3157 ( .Y(n6240), .A0(n6263), .A1(n6265) );
  and03 U3158 ( .Y(n6286), .A0(n6288), .A1(n6289), .A2(n6287) );
  nor02 U3159 ( .Y(n6289), .A0(n6246), .A1(n6290) );
  or02 U3160 ( .Y(n6290), .A0(n6291), .A1(n6249) );
  inv01 U3161 ( .Y(n6288), .A(n6258) );
  nor02 U3162 ( .Y(n6287), .A0(n6259), .A1(n6260) );
  nor02 U3163 ( .Y(n6285), .A0(n4359), .A1(n6261) );
  inv01 U3164 ( .Y(n6284), .A(n6263) );
  inv01 U3165 ( .Y(n6283), .A(n6267) );
  nand03 U3166 ( .Y(s_div_zeros_3_), .A0(n6277), .A1(n6278), .A2(n6276) );
  nor02 U3167 ( .Y(n6282), .A0(n6249), .A1(n6246) );
  nor02 U3168 ( .Y(n6281), .A0(n6255), .A1(n6257) );
  inv01 U3169 ( .Y(n6280), .A(n6256) );
  nor02 U3170 ( .Y(n6279), .A0(n6259), .A1(n6260) );
  inv01 U3171 ( .Y(n6277), .A(n6266) );
  inv01 U3172 ( .Y(n6276), .A(n6254) );
  inv01 U3173 ( .Y(n6274), .A(n6247) );
  or02 U3174 ( .Y(n6275), .A0(n6267), .A1(n6261) );
  nor02 U3175 ( .Y(n6273), .A0(n6262), .A1(n4359) );
  nor02 U3176 ( .Y(n6272), .A0(n6264), .A1(n6265) );
  inv01 U3178 ( .Y(n6164), .A(n6153) );
  nand02 U3179 ( .Y(n6153), .A0(n4378), .A1(n6103) );
  nand04 U3180 ( .Y(n6469), .A0(n4701), .A1(n4709), .A2(n6168), .A3(n6169) );
  inv01 U3181 ( .Y(n6174), .A(n6154) );
  nand02 U3182 ( .Y(n6154), .A0(n4380), .A1(n6098) );
  nand04 U3183 ( .Y(n6470), .A0(n4693), .A1(n4707), .A2(n6179), .A3(n6180) );
  inv01 U3184 ( .Y(n6181), .A(n6155) );
  nand02 U3185 ( .Y(n6155), .A0(n4376), .A1(n6103) );
  nand04 U3186 ( .Y(n6471), .A0(n4699), .A1(n5165), .A2(n6186), .A3(n6187) );
  inv01 U3187 ( .Y(n6172), .A(n6138) );
  inv01 U3188 ( .Y(n6189), .A(n5914) );
  inv01 U3189 ( .Y(n6203), .A(n6178) );
  and03 U3190 ( .Y(n6196), .A0(n6167), .A1(n6103), .A2(n6163) );
  inv01 U3191 ( .Y(n6218), .A(n6118) );
  inv01 U3192 ( .Y(n6220), .A(n6123) );
  inv01 U3193 ( .Y(n6206), .A(n6084) );
  inv01 U3194 ( .Y(n6211), .A(n6027) );
  inv01 U3195 ( .Y(n6217), .A(n5163) );
  nor02 U3196 ( .Y(n6171), .A0(n6238), .A1(s_div_zeros_0_) );
  nor02 U3197 ( .Y(n6170), .A0(n6239), .A1(s_div_zeros_1_) );
  nand02 U3198 ( .Y(n6188), .A0(n6047), .A1(s_div_zeros_0_) );
  nand02 U3199 ( .Y(n6150), .A0(n6173), .A1(opb_i[0]) );
  nand02 U3200 ( .Y(n6201), .A0(n6239), .A1(n6238) );
  inv01 U3201 ( .Y(n6252), .A(n6253) );
  inv01 U3202 ( .Y(n6213), .A(opb_i[17]) );
  inv01 U3203 ( .Y(n6239), .A(s_div_zeros_0_) );
  oai22 U3204 ( .Y(n6269), .A0(n6251), .A1(n4366), .B0(n6270), .B1(n6271) );
  nand04 U3205 ( .Y(s_div_zeros_4_), .A0(n6272), .A1(n6273), .A2(n5042), .A3(
        n6274) );
  and04 U3206 ( .Y(n6278), .A0(n6282), .A1(n6280), .A2(n6281), .A3(n6279) );
  nand04 U3207 ( .Y(s_div_zeros_2_), .A0(n6283), .A1(n6284), .A2(n6285), .A3(
        n6286) );
  inv01 U3208 ( .Y(n6200), .A(opb_i[19]) );
  and02 U3209 ( .Y(n6249), .A0(opb_i[9]), .A1(n4687) );
  and03 U3210 ( .Y(n6247), .A0(n6293), .A1(n6049), .A2(opb_i[6]) );
  and02 U3211 ( .Y(n6255), .A0(opb_i[13]), .A1(n5037) );
  and03 U3212 ( .Y(n6254), .A0(n6294), .A1(n6059), .A2(opb_i[14]) );
  and02 U3213 ( .Y(n6256), .A0(opb_i[15]), .A1(n6294) );
  and02 U3214 ( .Y(n6259), .A0(opb_i[11]), .A1(n6295) );
  and02 U3215 ( .Y(n6265), .A0(opb_i[5]), .A1(n4685) );
  and02 U3216 ( .Y(n6264), .A0(opb_i[7]), .A1(n6293) );
  and02 U3217 ( .Y(n6267), .A0(opb_i[3]), .A1(n6296) );
  and03 U3218 ( .Y(n6266), .A0(n6233), .A1(n6229), .A2(n5161) );
  nand02 U3219 ( .Y(n6253), .A0(n4447), .A1(n6158) );
  or02 U3220 ( .Y(n6162), .A0(n6271), .A1(opb_i[22]) );
  inv01 U3221 ( .Y(n6223), .A(opb_i[2]) );
  inv01 U3222 ( .Y(n6233), .A(opb_i[0]) );
  inv01 U3223 ( .Y(n6303), .A(n6305) );
  nand04 U3224 ( .Y(n6466), .A0(n4697), .A1(n4741), .A2(n6306), .A3(n6307) );
  inv01 U3225 ( .Y(n6310), .A(n6312) );
  nand04 U3226 ( .Y(n6467), .A0(n4695), .A1(n4739), .A2(n5064), .A3(n6315) );
  inv01 U3227 ( .Y(n6316), .A(n6318) );
  nand04 U3228 ( .Y(n6468), .A0(n4691), .A1(n5419), .A2(n6321), .A3(n6322) );
  inv01 U3229 ( .Y(n6323), .A(n5918) );
  inv01 U3230 ( .Y(n6337), .A(n6314) );
  inv01 U3231 ( .Y(n6343), .A(n6320) );
  inv01 U3232 ( .Y(n6355), .A(n6110) );
  inv01 U3233 ( .Y(n6358), .A(n6124) );
  inv01 U3234 ( .Y(n6373), .A(n6353) );
  nand02 U3235 ( .Y(n6305), .A0(n4431), .A1(n6092) );
  nand02 U3236 ( .Y(n6312), .A0(n6376), .A1(n6113) );
  nand02 U3237 ( .Y(n6318), .A0(n4429), .A1(n6113) );
  inv01 U3238 ( .Y(n6352), .A(n5699) );
  and02 U3239 ( .Y(n6308), .A0(s_dvd_zeros_1_), .A1(s_dvd_zeros_0_) );
  nand02 U3240 ( .Y(n6381), .A0(s_dvd_zeros_1_), .A1(n6382) );
  inv01 U3241 ( .Y(n6334), .A(n5926) );
  inv01 U3242 ( .Y(n6382), .A(s_dvd_zeros_0_) );
  inv01 U3243 ( .Y(n6335), .A(n6083) );
  nand04 U3244 ( .Y(s_dvd_zeros_4_), .A0(n6398), .A1(n6399), .A2(n6400), .A3(
        n6401) );
  and04 U3245 ( .Y(n6414), .A0(n6415), .A1(n6416), .A2(n6417), .A3(n6418) );
  nand02 U3246 ( .Y(n6372), .A0(n6083), .A1(opa_i[0]) );
  and02 U3247 ( .Y(n6383), .A0(opa_i[5]), .A1(n6429) );
  inv01 U3248 ( .Y(n6432), .A(n6420) );
  and03 U3249 ( .Y(n6394), .A0(n4361), .A1(n6044), .A2(n5159) );
  and02 U3250 ( .Y(n6393), .A0(opa_i[15]), .A1(n6433) );
  and03 U3251 ( .Y(n6395), .A0(n5092), .A1(n6080), .A2(opa_i[13]) );
  and02 U3252 ( .Y(n6397), .A0(opa_i[1]), .A1(n5159) );
  and03 U3253 ( .Y(n6396), .A0(n6435), .A1(n6074), .A2(opa_i[11]) );
  and02 U3254 ( .Y(n6404), .A0(opa_i[7]), .A1(n5093) );
  and02 U3255 ( .Y(n6384), .A0(opa_i[3]), .A1(n6437) );
  and02 U3256 ( .Y(n6390), .A0(opa_i[10]), .A1(n6430) );
  oai22 U3257 ( .Y(n6440), .A0(n6421), .A1(n6007), .B0(n6442), .B1(n6443) );
  and02 U3258 ( .Y(n6386), .A0(opa_i[12]), .A1(n6435) );
  and03 U3259 ( .Y(n6387), .A0(n5094), .A1(n6072), .A2(opa_i[6]) );
  and02 U3260 ( .Y(n6436), .A0(n6444), .A1(n6370) );
  and03 U3261 ( .Y(n6444), .A0(n6070), .A1(n5959), .A2(n6430) );
  and02 U3262 ( .Y(n6385), .A0(opa_i[14]), .A1(n5091) );
  and02 U3263 ( .Y(n6434), .A0(n6433), .A1(n5929) );
  and03 U3264 ( .Y(n6433), .A0(n6005), .A1(n5991), .A2(n6441) );
  nand02 U3265 ( .Y(n6420), .A0(n5014), .A1(n5086) );
  inv01 U3266 ( .Y(n6297), .A(opa_i[20]) );
  or02 U3267 ( .Y(n6301), .A0(n6443), .A1(opa_i[22]) );
  inv01 U3268 ( .Y(n6446), .A(s_expa_in_8_) );
  nand02 U3269 ( .Y(n6445), .A0(s_expa_in_7_), .A1(n6447) );
  inv01 U3270 ( .Y(n6447), .A(n5916) );
  ao21 U3271 ( .Y(n____return3540_6_), .A0(s_expa_in_6_), .A1(n6449), .B0(
        n5916) );
  nor02 U3272 ( .Y(n6448), .A0(n6449), .A1(s_expa_in_6_) );
  inv01 U3273 ( .Y(n6449), .A(n6450) );
  ao21 U3274 ( .Y(n____return3540_5_), .A0(s_expa_in_5_), .A1(n6451), .B0(
        n4319) );
  nor02 U3275 ( .Y(n6450), .A0(n6451), .A1(s_expa_in_5_) );
  inv01 U3276 ( .Y(n6451), .A(n6452) );
  ao21 U3277 ( .Y(n____return3540_4_), .A0(s_expa_in_4_), .A1(n6453), .B0(
        n4318) );
  nor02 U3278 ( .Y(n6452), .A0(n6453), .A1(s_expa_in_4_) );
  inv01 U3279 ( .Y(n6453), .A(n6454) );
  ao21 U3280 ( .Y(n____return3540_3_), .A0(s_expa_in_3_), .A1(n6455), .B0(
        n4317) );
  nor02 U3281 ( .Y(n6454), .A0(n6455), .A1(s_expa_in_3_) );
  inv01 U3282 ( .Y(n6455), .A(n6456) );
  ao21 U3283 ( .Y(n____return3540_2_), .A0(s_expa_in_2_), .A1(n6457), .B0(
        n4316) );
  nor02 U3284 ( .Y(n6456), .A0(n6457), .A1(s_expa_in_2_) );
  inv01 U3285 ( .Y(n6457), .A(n6458) );
  ao21 U3286 ( .Y(n____return3540_1_), .A0(s_expa_in_1_), .A1(s_expa_in_0_), 
        .B0(n6458) );
  nor02 U3287 ( .Y(n6458), .A0(s_expa_in_1_), .A1(s_expa_in_0_) );
  nand02 U3288 ( .Y(n____return3477_0_), .A0(n6271), .A1(n6459) );
  inv01 U3289 ( .Y(n6459), .A(opb_i[23]) );
  nand02 U3290 ( .Y(n6271), .A0(n6460), .A1(n6461) );
  nand02 U3291 ( .Y(n____return3431_0_), .A0(n6443), .A1(n6462) );
  inv01 U3292 ( .Y(n6462), .A(opa_i[23]) );
  nand02 U3293 ( .Y(n6443), .A0(n6463), .A1(n6464) );
  pre_norm_div_DW01_sub_10_1 sub_0_root_add_118_plus_plus_431 ( .A({
        n____return3612_9_, n____return3612_8_, n____return3612_7_, 
        n____return3612_6_, n____return3612_5_, n____return3612_4_, 
        n____return3612_3_, n____return3612_2_, n____return3612_1_, 
        n____return3612_0_}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n6110, 
        s_dvd_zeros_3_, n6089, s_dvd_zeros_1_, s_dvd_zeros_0_}), .CI(1'b0), 
        .DIFF({n____return3652_9_, n3654_8_, n____return3652_7_, 
        n____return3652_6_, n____return3652_5_, n____return3652_4_, 
        n____return3652_3_, n____return3652_2_, n____return3652_1_, 
        n____return3652_0_}) );
  pre_norm_div_DW01_add_10_1 add_1_root_add_118_plus_plus_431 ( .A({n5729, 
        n5695, n5697, n5692, n5693, n5562, n5563, n5564, n5561, 
        n____return3540_0_}), .B({n____return3578_9_, n____return3578_8_, 
        n____return3578_7_, n____return3578_6_, n____return3578_5_, 
        n____return3578_4_, n____return3578_3_, n____return3578_2_, 
        n____return3578_1_, n____return3578_0_}), .CI(1'b0), .SUM({
        n____return3612_9_, n____return3612_8_, n____return3612_7_, 
        n____return3612_6_, n____return3612_5_, n____return3612_4_, 
        n____return3612_3_, n____return3612_2_, n____return3612_1_, 
        n____return3612_0_}) );
  pre_norm_div_DW01_sub_10_0 sub_2_root_add_118_plus_plus_431 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, n6118, n6081, n6111, n6047, s_div_zeros_0_}), .B({
        s_expb_in_9_, s_expb_in_8_, s_expb_in_7_, s_expb_in_6_, s_expb_in_5_, 
        s_expb_in_4_, s_expb_in_3_, s_expb_in_2_, s_expb_in_1_, s_expb_in_0_}), 
        .CI(1'b0), .DIFF({n____return3578_9_, n____return3578_8_, 
        n____return3578_7_, n____return3578_6_, n____return3578_5_, 
        n____return3578_4_, n____return3578_3_, n____return3578_2_, 
        n____return3578_1_, n____return3578_0_}) );
endmodule


module post_norm_div_DW01_inc_9_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;
  wire   carry_8_, carry_7_, carry_6_, carry_5_, carry_4_, carry_3_, carry_2_;

  inv01 U5 ( .Y(SUM[0]), .A(A[0]) );
  xor2 U6 ( .Y(SUM[8]), .A0(carry_8_), .A1(A[8]) );
  hadd1 U1_1_1 ( .S(SUM[1]), .CO(carry_2_), .A(A[1]), .B(A[0]) );
  hadd1 U1_1_2 ( .S(SUM[2]), .CO(carry_3_), .A(A[2]), .B(carry_2_) );
  hadd1 U1_1_3 ( .S(SUM[3]), .CO(carry_4_), .A(A[3]), .B(carry_3_) );
  hadd1 U1_1_4 ( .S(SUM[4]), .CO(carry_5_), .A(A[4]), .B(carry_4_) );
  hadd1 U1_1_5 ( .S(SUM[5]), .CO(carry_6_), .A(A[5]), .B(carry_5_) );
  hadd1 U1_1_6 ( .S(SUM[6]), .CO(carry_7_), .A(A[6]), .B(carry_6_) );
  hadd1 U1_1_7 ( .S(SUM[7]), .CO(carry_8_), .A(A[7]), .B(carry_7_) );
endmodule


module post_norm_div_DW01_cmp2_6_0 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [5:0] A;
  input [5:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41;

  inv01 U6 ( .Y(n41), .A(B[0]) );
  inv01 U7 ( .Y(n30), .A(n15) );
  nor02 U8 ( .Y(n16), .A0(B[4]), .A1(n32) );
  nor02 U9 ( .Y(n17), .A0(B[3]), .A1(n33) );
  inv01 U10 ( .Y(n18), .A(n34) );
  nor02 U11 ( .Y(n15), .A0(n18), .A1(n19) );
  nor02 U12 ( .Y(n20), .A0(n16), .A1(n17) );
  inv01 U13 ( .Y(n19), .A(n20) );
  inv02 U14 ( .Y(n33), .A(A[3]) );
  inv02 U15 ( .Y(n32), .A(A[4]) );
  nand02 U16 ( .Y(n37), .A0(n40), .A1(n21) );
  inv01 U17 ( .Y(n22), .A(n35) );
  inv01 U18 ( .Y(n23), .A(B[2]) );
  inv01 U19 ( .Y(n24), .A(n39) );
  inv01 U20 ( .Y(n25), .A(n38) );
  nand02 U21 ( .Y(n26), .A0(n22), .A1(n23) );
  nand02 U22 ( .Y(n27), .A0(n24), .A1(n25) );
  nand02 U23 ( .Y(n28), .A0(n26), .A1(n27) );
  inv01 U24 ( .Y(n21), .A(n28) );
  inv01 U25 ( .Y(n36), .A(n37) );
  inv02 U26 ( .Y(n39), .A(A[1]) );
  inv02 U27 ( .Y(n35), .A(A[2]) );
  or02 U28 ( .Y(LT_LE), .A0(n29), .A1(B[5]) );
  nand02 U29 ( .Y(n29), .A0(n30), .A1(n31) );
  nand02 U30 ( .Y(n31), .A0(B[4]), .A1(n32) );
  ao221 U31 ( .Y(n34), .A0(n35), .A1(B[2]), .B0(n33), .B1(B[3]), .C0(n36) );
  ao21 U32 ( .Y(n40), .A0(n38), .A1(n39), .B0(B[1]) );
  nor02 U33 ( .Y(n38), .A0(n41), .A1(A[0]) );
endmodule


module post_norm_div_DW01_inc_25_0 ( A, SUM );
  input [24:0] A;
  output [24:0] SUM;
  wire   carry_23_, carry_22_, carry_21_, carry_20_, carry_19_, carry_18_,
         carry_17_, carry_16_, carry_15_, carry_14_, carry_13_, carry_12_,
         carry_11_, carry_10_, carry_9_, carry_8_, carry_7_, carry_6_,
         carry_5_, carry_4_, carry_3_, carry_2_;

  inv04 U5 ( .Y(SUM[0]), .A(A[0]) );
  hadd1 U1_1_1 ( .S(SUM[1]), .CO(carry_2_), .A(A[1]), .B(A[0]) );
  hadd1 U1_1_2 ( .S(SUM[2]), .CO(carry_3_), .A(A[2]), .B(carry_2_) );
  hadd1 U1_1_3 ( .S(SUM[3]), .CO(carry_4_), .A(A[3]), .B(carry_3_) );
  hadd1 U1_1_4 ( .S(SUM[4]), .CO(carry_5_), .A(A[4]), .B(carry_4_) );
  hadd1 U1_1_5 ( .S(SUM[5]), .CO(carry_6_), .A(A[5]), .B(carry_5_) );
  hadd1 U1_1_6 ( .S(SUM[6]), .CO(carry_7_), .A(A[6]), .B(carry_6_) );
  hadd1 U1_1_7 ( .S(SUM[7]), .CO(carry_8_), .A(A[7]), .B(carry_7_) );
  hadd1 U1_1_8 ( .S(SUM[8]), .CO(carry_9_), .A(A[8]), .B(carry_8_) );
  hadd1 U1_1_9 ( .S(SUM[9]), .CO(carry_10_), .A(A[9]), .B(carry_9_) );
  hadd1 U1_1_10 ( .S(SUM[10]), .CO(carry_11_), .A(A[10]), .B(carry_10_) );
  hadd1 U1_1_11 ( .S(SUM[11]), .CO(carry_12_), .A(A[11]), .B(carry_11_) );
  hadd1 U1_1_12 ( .S(SUM[12]), .CO(carry_13_), .A(A[12]), .B(carry_12_) );
  hadd1 U1_1_13 ( .S(SUM[13]), .CO(carry_14_), .A(A[13]), .B(carry_13_) );
  hadd1 U1_1_14 ( .S(SUM[14]), .CO(carry_15_), .A(A[14]), .B(carry_14_) );
  hadd1 U1_1_15 ( .S(SUM[15]), .CO(carry_16_), .A(A[15]), .B(carry_15_) );
  hadd1 U1_1_16 ( .S(SUM[16]), .CO(carry_17_), .A(A[16]), .B(carry_16_) );
  hadd1 U1_1_17 ( .S(SUM[17]), .CO(carry_18_), .A(A[17]), .B(carry_17_) );
  hadd1 U1_1_18 ( .S(SUM[18]), .CO(carry_19_), .A(A[18]), .B(carry_18_) );
  hadd1 U1_1_19 ( .S(SUM[19]), .CO(carry_20_), .A(A[19]), .B(carry_19_) );
  hadd1 U1_1_20 ( .S(SUM[20]), .CO(carry_21_), .A(A[20]), .B(carry_20_) );
  hadd1 U1_1_21 ( .S(SUM[21]), .CO(carry_22_), .A(A[21]), .B(carry_21_) );
  hadd1 U1_1_22 ( .S(SUM[22]), .CO(carry_23_), .A(A[22]), .B(carry_22_) );
  hadd1 U1_1_23 ( .S(SUM[23]), .CO(SUM[24]), .A(A[23]), .B(carry_23_) );
endmodule


module post_norm_div_DW01_dec_9_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;
  wire   carry_8_, carry_7_, carry_6_, carry_5_, carry_4_, carry_3_, n5, n7,
         n9, n11, n13, n15, n17, n19, n21, n22, n23, n24, n25, n26, n27;

  xor2 U6 ( .Y(n5), .A0(carry_8_), .A1(A[8]) );
  inv01 U7 ( .Y(SUM[8]), .A(n5) );
  xor2 U8 ( .Y(n7), .A0(A[2]), .A1(n22) );
  inv01 U9 ( .Y(SUM[2]), .A(n7) );
  xor2 U10 ( .Y(n9), .A0(A[6]), .A1(n27) );
  inv01 U11 ( .Y(SUM[6]), .A(n9) );
  xor2 U12 ( .Y(n11), .A0(A[7]), .A1(n26) );
  inv01 U13 ( .Y(SUM[7]), .A(n11) );
  xor2 U14 ( .Y(n13), .A0(A[3]), .A1(n23) );
  inv01 U15 ( .Y(SUM[3]), .A(n13) );
  xor2 U16 ( .Y(n15), .A0(A[5]), .A1(n25) );
  inv01 U17 ( .Y(SUM[5]), .A(n15) );
  xor2 U18 ( .Y(n17), .A0(A[1]), .A1(A[0]) );
  inv01 U19 ( .Y(SUM[1]), .A(n17) );
  xor2 U20 ( .Y(n19), .A0(A[4]), .A1(n24) );
  inv01 U21 ( .Y(SUM[4]), .A(n19) );
  nor02 U22 ( .Y(n21), .A0(A[1]), .A1(A[0]) );
  inv02 U23 ( .Y(n22), .A(n21) );
  buf02 U24 ( .Y(n23), .A(carry_3_) );
  buf02 U25 ( .Y(n24), .A(carry_4_) );
  buf02 U26 ( .Y(n25), .A(carry_5_) );
  buf02 U27 ( .Y(n26), .A(carry_7_) );
  buf02 U28 ( .Y(n27), .A(carry_6_) );
  inv01 U29 ( .Y(SUM[0]), .A(A[0]) );
  or02 U1_B_2 ( .Y(carry_3_), .A0(A[2]), .A1(n22) );
  or02 U1_B_3 ( .Y(carry_4_), .A0(A[3]), .A1(n23) );
  or02 U1_B_4 ( .Y(carry_5_), .A0(A[4]), .A1(n24) );
  or02 U1_B_5 ( .Y(carry_6_), .A0(A[5]), .A1(n25) );
  or02 U1_B_6 ( .Y(carry_7_), .A0(A[6]), .A1(n27) );
  or02 U1_B_7 ( .Y(carry_8_), .A0(A[7]), .A1(n26) );
endmodule


module post_norm_div ( clk_i, opa_i, opb_i, qutnt_i, rmndr_i, exp_10_i, sign_i, 
        rmode_i, output_o, ine_o );
  input [31:0] opa_i;
  input [31:0] opb_i;
  input [26:0] qutnt_i;
  input [26:0] rmndr_i;
  input [9:0] exp_10_i;
  input [1:0] rmode_i;
  output [31:0] output_o;
  input clk_i, sign_i;
  output ine_o;
  wire   s_output_o_31_, s_output_o_30_, s_output_o_29_, s_output_o_28_,
         s_output_o_27_, s_output_o_26_, s_output_o_25_, s_output_o_24_,
         s_output_o_23_, s_output_o_22_, s_ine_o, v_shl433_0_, s_fraco1_26_,
         s_fraco1_25_, s_fraco1_24_, s_fraco1_23_, s_fraco1_22_, s_fraco1_21_,
         s_fraco1_20_, s_fraco1_19_, s_fraco1_18_, s_fraco1_17_, s_fraco1_16_,
         s_fraco1_15_, s_fraco1_14_, s_fraco1_13_, s_fraco1_12_, s_fraco1_11_,
         s_fraco1_10_, s_fraco1_9_, s_fraco1_8_, s_fraco1_7_, s_fraco1_6_,
         s_fraco1_5_, s_fraco1_4_, s_fraco1_3_, s_fraco1_0_, s_round, s_sign_i,
         s_expo3_7_, s_expo3_6_, s_expo3_5_, s_expo3_4_, s_expo3_3_,
         s_expo3_2_, s_expo3_1_, s_expo3_0_, s_fraco2_22_, s_opa_i_30_,
         s_opa_i_29_, s_opa_i_28_, s_opa_i_25_, s_opa_i_24_, s_opa_i_23_,
         s_opa_i_21_, s_opa_i_20_, s_opa_i_16_, s_opa_i_15_, s_opa_i_14_,
         s_opa_i_11_, s_opa_i_10_, s_opa_i_6_, s_opa_i_5_, s_opa_i_4_,
         s_opa_i_1_, s_opa_i_0_, s_opb_i_30_, s_opb_i_29_, s_opb_i_28_,
         s_opb_i_25_, s_opb_i_24_, s_opb_i_23_, s_opb_i_21_, s_opb_i_20_,
         s_opb_i_16_, s_opb_i_15_, s_opb_i_14_, s_opb_i_11_, s_opb_i_10_,
         s_opb_i_6_, s_opb_i_5_, s_opb_i_4_, s_opb_i_1_, s_opb_i_0_,
         s_rmndr_i_23_, s_rmndr_i_22_, s_rmndr_i_21_, s_rmndr_i_17_,
         s_rmndr_i_16_, s_rmndr_i_15_, s_rmndr_i_10_, s_rmndr_i_5_,
         s_rmndr_i_4_, s_rmndr_i_3_, s_rmndr_i_0_, s_exp_10_i_8_,
         s_exp_10_i_7_, s_exp_10_i_6_, s_exp_10_i_5_, s_exp_10_i_4_,
         s_exp_10_i_3_, s_exp_10_i_2_, s_exp_10_i_1_, s_exp_10_i_0_,
         s_rmode_i_1_, s_rmode_i_0_, s_expo1480_0_, s_shr1482_5_, s_shr1482_4_,
         s_shr1482_3_, s_shr1482_2_, s_shr1482_1_, s_shr1482_0_, s_shr1_5_,
         s_shr1_4_, s_shr1_3_, s_shr1_2_, s_shr1_1_, s_shr1_0_, s_shl1_4_,
         s_shl1_3_, s_shl1_2_, s_shl1_1_, s_shl1_0_, s_fraco1812_26_,
         s_fraco1812_25_, s_fraco1812_24_, s_fraco1812_23_, s_fraco1812_22_,
         s_fraco1812_21_, s_fraco1812_20_, s_fraco1812_19_, s_fraco1812_18_,
         s_fraco1812_17_, s_fraco1812_16_, s_fraco1812_15_, s_fraco1812_14_,
         s_fraco1812_13_, s_fraco1812_12_, s_fraco1812_11_, s_fraco1812_10_,
         s_fraco1812_9_, s_fraco1812_8_, s_fraco1812_7_, s_fraco1812_6_,
         s_fraco1812_5_, s_fraco1812_4_, s_fraco1812_3_, s_fraco1812_2_,
         s_fraco1812_1_, s_fraco1812_0_, n1238_8_, n____return1236_7_,
         n____return1236_6_, n____return1236_5_, n____return1236_4_,
         n____return1236_3_, n____return1236_2_, n____return1236_1_,
         n____return1236_0_, s_r_zeros_4_, s_r_zeros_3_, s_r_zeros_2_,
         s_r_zeros_1_, s_r_zeros_0_, n____return2916, n____return2878_3_,
         n____return2878_1_, n3243_24_, n____return3241_23_,
         n____return3241_22_, n____return3241_21_, n____return3241_20_,
         n____return3241_19_, n____return3241_18_, n____return3241_17_,
         n____return3241_16_, n____return3241_15_, n____return3241_14_,
         n____return3241_13_, n____return3241_12_, n____return3241_11_,
         n____return3241_10_, n____return3241_9_, n____return3241_8_,
         n____return3241_7_, n____return3241_6_, n____return3241_5_,
         n____return3241_4_, n____return3241_3_, n____return3241_2_,
         n____return3241_1_, n____return3241_0_, s_expo33281_8_,
         s_expo33281_7_, s_expo33281_6_, s_expo33281_5_, s_expo33281_4_,
         s_expo33281_3_, s_expo33281_2_, s_expo33281_1_, s_expo33281_0_,
         s_fraco23289_22_, s_fraco23289_21_, s_fraco23289_20_,
         s_fraco23289_19_, s_fraco23289_18_, s_fraco23289_17_,
         s_fraco23289_16_, s_fraco23289_15_, s_fraco23289_14_,
         s_fraco23289_13_, s_fraco23289_12_, s_fraco23289_11_,
         s_fraco23289_10_, s_fraco23289_9_, s_fraco23289_8_, s_fraco23289_7_,
         s_fraco23289_6_, s_fraco23289_5_, s_fraco23289_4_, s_fraco23289_3_,
         s_fraco23289_2_, s_fraco23289_1_, s_fraco23289_0_, n3318_7_,
         n____return3316_8_, n____return3316_6_, n____return3316_5_,
         n____return3316_4_, n____return3316_3_, n____return3316_2_,
         n____return3316_1_, n____return3316_0_, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900;
  wire   [26:0] s_qutnt_i;
  wire   [8:0] s_expo1;
  wire   [8:0] s_expo2;

  dff s_shl1_reg_5_ ( .QB(n8882), .D(1'b0), .CLK(clk_i) );
  dff s_shl1_reg_4_ ( .Q(s_shl1_4_), .D(1'b0), .CLK(clk_i) );
  dff s_shl1_reg_3_ ( .Q(s_shl1_3_), .D(1'b0), .CLK(clk_i) );
  dff s_shl1_reg_2_ ( .Q(s_shl1_2_), .D(1'b0), .CLK(clk_i) );
  dff s_shl1_reg_1_ ( .Q(s_shl1_1_), .D(1'b0), .CLK(clk_i) );
  dff s_expa_reg_7_ ( .QB(n8841), .D(opa_i[30]), .CLK(clk_i) );
  dff s_expa_reg_6_ ( .QB(n8840), .D(opa_i[29]), .CLK(clk_i) );
  dff s_expa_reg_5_ ( .QB(n8839), .D(opa_i[28]), .CLK(clk_i) );
  dff s_expa_reg_4_ ( .QB(n8838), .D(opa_i[27]), .CLK(clk_i) );
  dff s_expa_reg_3_ ( .QB(n8845), .D(opa_i[26]), .CLK(clk_i) );
  dff s_expa_reg_2_ ( .QB(n8844), .D(opa_i[25]), .CLK(clk_i) );
  dff s_expa_reg_1_ ( .QB(n8843), .D(opa_i[24]), .CLK(clk_i) );
  dff s_expa_reg_0_ ( .QB(n8842), .D(opa_i[23]), .CLK(clk_i) );
  dff s_expb_reg_7_ ( .QB(n8833), .D(opb_i[30]), .CLK(clk_i) );
  dff s_expb_reg_6_ ( .QB(n8832), .D(opb_i[29]), .CLK(clk_i) );
  dff s_expb_reg_5_ ( .QB(n8831), .D(opb_i[28]), .CLK(clk_i) );
  dff s_expb_reg_4_ ( .QB(n8830), .D(opb_i[27]), .CLK(clk_i) );
  dff s_expb_reg_3_ ( .QB(n8837), .D(opb_i[26]), .CLK(clk_i) );
  dff s_expb_reg_2_ ( .QB(n8836), .D(opb_i[25]), .CLK(clk_i) );
  dff s_expb_reg_1_ ( .QB(n8835), .D(opb_i[24]), .CLK(clk_i) );
  dff s_expb_reg_0_ ( .QB(n8834), .D(opb_i[23]), .CLK(clk_i) );
  dff s_qutnt_i_reg_26_ ( .Q(s_qutnt_i[26]), .D(qutnt_i[26]), .CLK(clk_i) );
  dff s_qutnt_i_reg_25_ ( .Q(s_qutnt_i[25]), .D(qutnt_i[25]), .CLK(clk_i) );
  dff s_qutnt_i_reg_24_ ( .Q(s_qutnt_i[24]), .D(qutnt_i[24]), .CLK(clk_i) );
  dff s_qutnt_i_reg_23_ ( .Q(s_qutnt_i[23]), .D(qutnt_i[23]), .CLK(clk_i) );
  dff s_qutnt_i_reg_22_ ( .Q(s_qutnt_i[22]), .D(qutnt_i[22]), .CLK(clk_i) );
  dff s_qutnt_i_reg_21_ ( .Q(s_qutnt_i[21]), .D(qutnt_i[21]), .CLK(clk_i) );
  dff s_qutnt_i_reg_20_ ( .Q(s_qutnt_i[20]), .D(qutnt_i[20]), .CLK(clk_i) );
  dff s_qutnt_i_reg_19_ ( .Q(s_qutnt_i[19]), .D(qutnt_i[19]), .CLK(clk_i) );
  dff s_qutnt_i_reg_18_ ( .Q(s_qutnt_i[18]), .D(qutnt_i[18]), .CLK(clk_i) );
  dff s_qutnt_i_reg_17_ ( .Q(s_qutnt_i[17]), .D(qutnt_i[17]), .CLK(clk_i) );
  dff s_qutnt_i_reg_16_ ( .Q(s_qutnt_i[16]), .D(qutnt_i[16]), .CLK(clk_i) );
  dff s_qutnt_i_reg_15_ ( .Q(s_qutnt_i[15]), .D(qutnt_i[15]), .CLK(clk_i) );
  dff s_qutnt_i_reg_14_ ( .Q(s_qutnt_i[14]), .D(qutnt_i[14]), .CLK(clk_i) );
  dff s_qutnt_i_reg_13_ ( .Q(s_qutnt_i[13]), .D(qutnt_i[13]), .CLK(clk_i) );
  dff s_qutnt_i_reg_12_ ( .Q(s_qutnt_i[12]), .D(qutnt_i[12]), .CLK(clk_i) );
  dff s_qutnt_i_reg_11_ ( .Q(s_qutnt_i[11]), .D(qutnt_i[11]), .CLK(clk_i) );
  dff s_qutnt_i_reg_10_ ( .Q(s_qutnt_i[10]), .D(qutnt_i[10]), .CLK(clk_i) );
  dff s_qutnt_i_reg_9_ ( .Q(s_qutnt_i[9]), .D(qutnt_i[9]), .CLK(clk_i) );
  dff s_qutnt_i_reg_8_ ( .Q(s_qutnt_i[8]), .D(qutnt_i[8]), .CLK(clk_i) );
  dff s_qutnt_i_reg_7_ ( .Q(s_qutnt_i[7]), .D(qutnt_i[7]), .CLK(clk_i) );
  dff s_qutnt_i_reg_6_ ( .Q(s_qutnt_i[6]), .QB(n8308), .D(qutnt_i[6]), .CLK(
        clk_i) );
  dff s_qutnt_i_reg_5_ ( .Q(s_qutnt_i[5]), .D(qutnt_i[5]), .CLK(clk_i) );
  dff s_qutnt_i_reg_4_ ( .Q(s_qutnt_i[4]), .D(qutnt_i[4]), .CLK(clk_i) );
  dff s_qutnt_i_reg_3_ ( .Q(s_qutnt_i[3]), .D(qutnt_i[3]), .CLK(clk_i) );
  dff s_qutnt_i_reg_2_ ( .Q(s_qutnt_i[2]), .D(qutnt_i[2]), .CLK(clk_i) );
  dff s_qutnt_i_reg_1_ ( .Q(s_qutnt_i[1]), .D(qutnt_i[1]), .CLK(clk_i) );
  dff s_qutnt_i_reg_0_ ( .Q(s_qutnt_i[0]), .D(qutnt_i[0]), .CLK(clk_i) );
  dff s_rmndr_i_reg_26_ ( .QB(n8890), .D(rmndr_i[26]), .CLK(clk_i) );
  dff s_rmndr_i_reg_25_ ( .QB(n8889), .D(rmndr_i[25]), .CLK(clk_i) );
  dff s_rmndr_i_reg_24_ ( .QB(n8888), .D(rmndr_i[24]), .CLK(clk_i) );
  dff s_rmndr_i_reg_23_ ( .Q(s_rmndr_i_23_), .D(rmndr_i[23]), .CLK(clk_i) );
  dff s_rmndr_i_reg_22_ ( .Q(s_rmndr_i_22_), .D(rmndr_i[22]), .CLK(clk_i) );
  dff s_rmndr_i_reg_21_ ( .Q(s_rmndr_i_21_), .D(rmndr_i[21]), .CLK(clk_i) );
  dff s_rmndr_i_reg_20_ ( .QB(n8893), .D(rmndr_i[20]), .CLK(clk_i) );
  dff s_rmndr_i_reg_19_ ( .QB(n8895), .D(rmndr_i[19]), .CLK(clk_i) );
  dff s_rmndr_i_reg_18_ ( .QB(n8894), .D(rmndr_i[18]), .CLK(clk_i) );
  dff s_rmndr_i_reg_17_ ( .Q(s_rmndr_i_17_), .D(rmndr_i[17]), .CLK(clk_i) );
  dff s_rmndr_i_reg_16_ ( .Q(s_rmndr_i_16_), .D(rmndr_i[16]), .CLK(clk_i) );
  dff s_rmndr_i_reg_15_ ( .Q(s_rmndr_i_15_), .D(rmndr_i[15]), .CLK(clk_i) );
  dff s_rmndr_i_reg_14_ ( .QB(n8899), .D(rmndr_i[14]), .CLK(clk_i) );
  dff s_rmndr_i_reg_13_ ( .QB(n8898), .D(rmndr_i[13]), .CLK(clk_i) );
  dff s_rmndr_i_reg_12_ ( .QB(n8897), .D(rmndr_i[12]), .CLK(clk_i) );
  dff s_rmndr_i_reg_11_ ( .QB(n8896), .D(rmndr_i[11]), .CLK(clk_i) );
  dff s_rmndr_i_reg_10_ ( .Q(s_rmndr_i_10_), .D(rmndr_i[10]), .CLK(clk_i) );
  dff s_rmndr_i_reg_9_ ( .QB(n8887), .D(rmndr_i[9]), .CLK(clk_i) );
  dff s_rmndr_i_reg_8_ ( .QB(n8886), .D(rmndr_i[8]), .CLK(clk_i) );
  dff s_rmndr_i_reg_7_ ( .QB(n8885), .D(rmndr_i[7]), .CLK(clk_i) );
  dff s_rmndr_i_reg_6_ ( .QB(n8884), .D(rmndr_i[6]), .CLK(clk_i) );
  dff s_rmndr_i_reg_5_ ( .Q(s_rmndr_i_5_), .D(rmndr_i[5]), .CLK(clk_i) );
  dff s_rmndr_i_reg_4_ ( .Q(s_rmndr_i_4_), .D(rmndr_i[4]), .CLK(clk_i) );
  dff s_rmndr_i_reg_3_ ( .Q(s_rmndr_i_3_), .D(rmndr_i[3]), .CLK(clk_i) );
  dff s_rmndr_i_reg_2_ ( .QB(n8891), .D(rmndr_i[2]), .CLK(clk_i) );
  dff s_rmndr_i_reg_1_ ( .QB(n8892), .D(rmndr_i[1]), .CLK(clk_i) );
  dff s_rmndr_i_reg_0_ ( .Q(s_rmndr_i_0_), .D(rmndr_i[0]), .CLK(clk_i) );
  dff s_exp_10_i_reg_9_ ( .QB(n8900), .D(exp_10_i[9]), .CLK(clk_i) );
  dff s_exp_10_i_reg_8_ ( .Q(s_exp_10_i_8_), .D(exp_10_i[8]), .CLK(clk_i) );
  dff s_exp_10_i_reg_7_ ( .Q(s_exp_10_i_7_), .D(exp_10_i[7]), .CLK(clk_i) );
  dff s_exp_10_i_reg_6_ ( .Q(s_exp_10_i_6_), .D(exp_10_i[6]), .CLK(clk_i) );
  dff s_exp_10_i_reg_5_ ( .Q(s_exp_10_i_5_), .D(exp_10_i[5]), .CLK(clk_i) );
  dff s_exp_10_i_reg_4_ ( .Q(s_exp_10_i_4_), .D(exp_10_i[4]), .CLK(clk_i) );
  dff s_exp_10_i_reg_3_ ( .Q(s_exp_10_i_3_), .D(exp_10_i[3]), .CLK(clk_i) );
  dff s_exp_10_i_reg_2_ ( .Q(s_exp_10_i_2_), .D(exp_10_i[2]), .CLK(clk_i) );
  dff s_exp_10_i_reg_1_ ( .Q(s_exp_10_i_1_), .D(exp_10_i[1]), .CLK(clk_i) );
  dff s_exp_10_i_reg_0_ ( .Q(s_exp_10_i_0_), .D(exp_10_i[0]), .CLK(clk_i) );
  dff s_rmode_i_reg_1_ ( .Q(s_rmode_i_1_), .D(rmode_i[1]), .CLK(clk_i) );
  dff s_rmode_i_reg_0_ ( .Q(s_rmode_i_0_), .D(rmode_i[0]), .CLK(clk_i) );
  dff output_o_reg_31_ ( .Q(output_o[31]), .D(s_output_o_31_), .CLK(clk_i) );
  dff output_o_reg_30_ ( .Q(output_o[30]), .D(s_output_o_30_), .CLK(clk_i) );
  dff output_o_reg_29_ ( .Q(output_o[29]), .D(s_output_o_29_), .CLK(clk_i) );
  dff output_o_reg_28_ ( .Q(output_o[28]), .D(s_output_o_28_), .CLK(clk_i) );
  dff output_o_reg_27_ ( .Q(output_o[27]), .D(s_output_o_27_), .CLK(clk_i) );
  dff output_o_reg_26_ ( .Q(output_o[26]), .D(s_output_o_26_), .CLK(clk_i) );
  dff output_o_reg_25_ ( .Q(output_o[25]), .D(s_output_o_25_), .CLK(clk_i) );
  dff output_o_reg_24_ ( .Q(output_o[24]), .D(s_output_o_24_), .CLK(clk_i) );
  dff output_o_reg_23_ ( .Q(output_o[23]), .D(s_output_o_23_), .CLK(clk_i) );
  dff output_o_reg_22_ ( .Q(output_o[22]), .D(s_output_o_22_), .CLK(clk_i) );
  dff output_o_reg_21_ ( .Q(output_o[21]), .D(n5211), .CLK(clk_i) );
  dff output_o_reg_20_ ( .Q(output_o[20]), .D(n5197), .CLK(clk_i) );
  dff output_o_reg_19_ ( .Q(output_o[19]), .D(n5221), .CLK(clk_i) );
  dff output_o_reg_18_ ( .Q(output_o[18]), .D(n5193), .CLK(clk_i) );
  dff output_o_reg_17_ ( .Q(output_o[17]), .D(n5189), .CLK(clk_i) );
  dff output_o_reg_16_ ( .Q(output_o[16]), .D(n5215), .CLK(clk_i) );
  dff output_o_reg_15_ ( .Q(output_o[15]), .D(n5225), .CLK(clk_i) );
  dff output_o_reg_14_ ( .Q(output_o[14]), .D(n5227), .CLK(clk_i) );
  dff output_o_reg_13_ ( .Q(output_o[13]), .D(n5207), .CLK(clk_i) );
  dff output_o_reg_12_ ( .Q(output_o[12]), .D(n5209), .CLK(clk_i) );
  dff output_o_reg_11_ ( .Q(output_o[11]), .D(n5187), .CLK(clk_i) );
  dff output_o_reg_10_ ( .Q(output_o[10]), .D(n5223), .CLK(clk_i) );
  dff output_o_reg_9_ ( .Q(output_o[9]), .D(n5217), .CLK(clk_i) );
  dff output_o_reg_8_ ( .Q(output_o[8]), .D(n5205), .CLK(clk_i) );
  dff output_o_reg_7_ ( .Q(output_o[7]), .D(n5219), .CLK(clk_i) );
  dff output_o_reg_6_ ( .Q(output_o[6]), .D(n5199), .CLK(clk_i) );
  dff output_o_reg_5_ ( .Q(output_o[5]), .D(n5231), .CLK(clk_i) );
  dff output_o_reg_4_ ( .Q(output_o[4]), .D(n5201), .CLK(clk_i) );
  dff output_o_reg_3_ ( .Q(output_o[3]), .D(n5233), .CLK(clk_i) );
  dff output_o_reg_2_ ( .Q(output_o[2]), .D(n5191), .CLK(clk_i) );
  dff output_o_reg_1_ ( .Q(output_o[1]), .D(n5203), .CLK(clk_i) );
  dff output_o_reg_0_ ( .Q(output_o[0]), .D(n5229), .CLK(clk_i) );
  dff s_expo1_reg_8_ ( .Q(s_expo1[8]), .D(n5175), .CLK(clk_i) );
  dff s_expo1_reg_7_ ( .Q(s_expo1[7]), .D(n5173), .CLK(clk_i) );
  dff s_expo1_reg_6_ ( .Q(s_expo1[6]), .D(n5182), .CLK(clk_i) );
  dff s_expo1_reg_5_ ( .Q(s_expo1[5]), .D(n5400), .CLK(clk_i) );
  dff s_expo1_reg_4_ ( .Q(s_expo1[4]), .D(n5184), .CLK(clk_i) );
  dff s_expo1_reg_3_ ( .Q(s_expo1[3]), .D(n5171), .CLK(clk_i) );
  dff s_expo1_reg_2_ ( .Q(s_expo1[2]), .D(n5474), .CLK(clk_i) );
  dff s_expo1_reg_1_ ( .Q(s_expo1[1]), .D(n5466), .CLK(clk_i) );
  dff s_expo1_reg_0_ ( .Q(s_expo1[0]), .D(s_expo1480_0_), .CLK(clk_i) );
  dff s_shr1_reg_5_ ( .Q(s_shr1_5_), .D(s_shr1482_5_), .CLK(clk_i) );
  dff s_shr1_reg_4_ ( .Q(s_shr1_4_), .D(s_shr1482_4_), .CLK(clk_i) );
  dff s_shr1_reg_3_ ( .Q(s_shr1_3_), .D(s_shr1482_3_), .CLK(clk_i) );
  dff s_shr1_reg_2_ ( .Q(s_shr1_2_), .D(s_shr1482_2_), .CLK(clk_i) );
  dff s_shr1_reg_1_ ( .Q(s_shr1_1_), .D(s_shr1482_1_), .CLK(clk_i) );
  dff s_shr1_reg_0_ ( .Q(s_shr1_0_), .D(s_shr1482_0_), .CLK(clk_i) );
  dff s_fraco1_reg_26_ ( .Q(s_fraco1_26_), .QB(n8324), .D(s_fraco1812_26_), 
        .CLK(clk_i) );
  dff s_fraco1_reg_25_ ( .Q(s_fraco1_25_), .QB(n8868), .D(s_fraco1812_25_), 
        .CLK(clk_i) );
  dff s_fraco1_reg_24_ ( .Q(s_fraco1_24_), .QB(n8869), .D(s_fraco1812_24_), 
        .CLK(clk_i) );
  dff s_fraco1_reg_23_ ( .Q(s_fraco1_23_), .QB(n8870), .D(s_fraco1812_23_), 
        .CLK(clk_i) );
  dff s_fraco1_reg_22_ ( .Q(s_fraco1_22_), .QB(n8872), .D(s_fraco1812_22_), 
        .CLK(clk_i) );
  dff s_fraco1_reg_21_ ( .Q(s_fraco1_21_), .QB(n8873), .D(s_fraco1812_21_), 
        .CLK(clk_i) );
  dff s_fraco1_reg_20_ ( .Q(s_fraco1_20_), .QB(n8874), .D(s_fraco1812_20_), 
        .CLK(clk_i) );
  dff s_fraco1_reg_19_ ( .Q(s_fraco1_19_), .QB(n8875), .D(s_fraco1812_19_), 
        .CLK(clk_i) );
  dff s_fraco1_reg_18_ ( .Q(s_fraco1_18_), .QB(n8876), .D(s_fraco1812_18_), 
        .CLK(clk_i) );
  dff s_fraco1_reg_17_ ( .Q(s_fraco1_17_), .QB(n8877), .D(s_fraco1812_17_), 
        .CLK(clk_i) );
  dff s_fraco1_reg_16_ ( .Q(s_fraco1_16_), .QB(n8878), .D(s_fraco1812_16_), 
        .CLK(clk_i) );
  dff s_fraco1_reg_15_ ( .Q(s_fraco1_15_), .QB(n8879), .D(s_fraco1812_15_), 
        .CLK(clk_i) );
  dff s_fraco1_reg_14_ ( .Q(s_fraco1_14_), .QB(n8880), .D(s_fraco1812_14_), 
        .CLK(clk_i) );
  dff s_fraco1_reg_13_ ( .Q(s_fraco1_13_), .QB(n8881), .D(s_fraco1812_13_), 
        .CLK(clk_i) );
  dff s_fraco1_reg_12_ ( .Q(s_fraco1_12_), .QB(n8860), .D(s_fraco1812_12_), 
        .CLK(clk_i) );
  dff s_fraco1_reg_11_ ( .Q(s_fraco1_11_), .QB(n8861), .D(s_fraco1812_11_), 
        .CLK(clk_i) );
  dff s_fraco1_reg_10_ ( .Q(s_fraco1_10_), .QB(n8862), .D(s_fraco1812_10_), 
        .CLK(clk_i) );
  dff s_fraco1_reg_9_ ( .Q(s_fraco1_9_), .QB(n8863), .D(s_fraco1812_9_), .CLK(
        clk_i) );
  dff s_fraco1_reg_8_ ( .Q(s_fraco1_8_), .QB(n8864), .D(s_fraco1812_8_), .CLK(
        clk_i) );
  dff s_fraco1_reg_7_ ( .Q(s_fraco1_7_), .QB(n8865), .D(s_fraco1812_7_), .CLK(
        clk_i) );
  dff s_fraco1_reg_6_ ( .Q(s_fraco1_6_), .QB(n8866), .D(s_fraco1812_6_), .CLK(
        clk_i) );
  dff s_fraco1_reg_5_ ( .Q(s_fraco1_5_), .QB(n8867), .D(s_fraco1812_5_), .CLK(
        clk_i) );
  dff s_fraco1_reg_4_ ( .Q(s_fraco1_4_), .QB(n8871), .D(s_fraco1812_4_), .CLK(
        clk_i) );
  dff s_fraco1_reg_3_ ( .Q(s_fraco1_3_), .D(s_fraco1812_3_), .CLK(clk_i) );
  dff s_fraco1_reg_2_ ( .Q(n8883), .D(s_fraco1812_2_), .CLK(clk_i) );
  dff s_fraco1_reg_1_ ( .Q(s_round), .D(s_fraco1812_1_), .CLK(clk_i) );
  dff s_fraco1_reg_0_ ( .Q(s_fraco1_0_), .D(s_fraco1812_0_), .CLK(clk_i) );
  dff s_expo3_reg_8_ ( .QB(n8859), .D(s_expo33281_8_), .CLK(clk_i) );
  dff s_expo3_reg_7_ ( .Q(s_expo3_7_), .D(s_expo33281_7_), .CLK(clk_i) );
  dff s_expo3_reg_6_ ( .Q(s_expo3_6_), .D(s_expo33281_6_), .CLK(clk_i) );
  dff s_expo3_reg_5_ ( .Q(s_expo3_5_), .D(s_expo33281_5_), .CLK(clk_i) );
  dff s_expo3_reg_4_ ( .Q(s_expo3_4_), .D(s_expo33281_4_), .CLK(clk_i) );
  dff s_expo3_reg_3_ ( .Q(s_expo3_3_), .D(s_expo33281_3_), .CLK(clk_i) );
  dff s_expo3_reg_2_ ( .Q(s_expo3_2_), .D(s_expo33281_2_), .CLK(clk_i) );
  dff s_expo3_reg_1_ ( .Q(s_expo3_1_), .D(s_expo33281_1_), .CLK(clk_i) );
  dff s_expo3_reg_0_ ( .Q(s_expo3_0_), .D(s_expo33281_0_), .CLK(clk_i) );
  dff s_opa_i_reg_30_ ( .Q(s_opa_i_30_), .D(opa_i[30]), .CLK(clk_i) );
  dff s_opa_i_reg_29_ ( .Q(s_opa_i_29_), .D(opa_i[29]), .CLK(clk_i) );
  dff s_opa_i_reg_28_ ( .Q(s_opa_i_28_), .D(opa_i[28]), .CLK(clk_i) );
  dff s_opa_i_reg_27_ ( .QB(n8829), .D(opa_i[27]), .CLK(clk_i) );
  dff s_opa_i_reg_26_ ( .QB(n8828), .D(opa_i[26]), .CLK(clk_i) );
  dff s_opa_i_reg_25_ ( .Q(s_opa_i_25_), .D(opa_i[25]), .CLK(clk_i) );
  dff s_opa_i_reg_24_ ( .Q(s_opa_i_24_), .D(opa_i[24]), .CLK(clk_i) );
  dff s_opa_i_reg_23_ ( .Q(s_opa_i_23_), .D(opa_i[23]), .CLK(clk_i) );
  dff s_opa_i_reg_22_ ( .QB(n8820), .D(opa_i[22]), .CLK(clk_i) );
  dff s_opa_i_reg_21_ ( .Q(s_opa_i_21_), .D(opa_i[21]), .CLK(clk_i) );
  dff s_opa_i_reg_20_ ( .Q(s_opa_i_20_), .D(opa_i[20]), .CLK(clk_i) );
  dff s_opa_i_reg_19_ ( .QB(n8825), .D(opa_i[19]), .CLK(clk_i) );
  dff s_opa_i_reg_18_ ( .QB(n8824), .D(opa_i[18]), .CLK(clk_i) );
  dff s_opa_i_reg_17_ ( .QB(n8823), .D(opa_i[17]), .CLK(clk_i) );
  dff s_opa_i_reg_16_ ( .Q(s_opa_i_16_), .D(opa_i[16]), .CLK(clk_i) );
  dff s_opa_i_reg_15_ ( .Q(s_opa_i_15_), .D(opa_i[15]), .CLK(clk_i) );
  dff s_opa_i_reg_14_ ( .Q(s_opa_i_14_), .D(opa_i[14]), .CLK(clk_i) );
  dff s_opa_i_reg_13_ ( .QB(n8827), .D(opa_i[13]), .CLK(clk_i) );
  dff s_opa_i_reg_12_ ( .QB(n8826), .D(opa_i[12]), .CLK(clk_i) );
  dff s_opa_i_reg_11_ ( .Q(s_opa_i_11_), .D(opa_i[11]), .CLK(clk_i) );
  dff s_opa_i_reg_10_ ( .Q(s_opa_i_10_), .D(opa_i[10]), .CLK(clk_i) );
  dff s_opa_i_reg_9_ ( .QB(n8819), .D(opa_i[9]), .CLK(clk_i) );
  dff s_opa_i_reg_8_ ( .QB(n8818), .D(opa_i[8]), .CLK(clk_i) );
  dff s_opa_i_reg_7_ ( .QB(n8817), .D(opa_i[7]), .CLK(clk_i) );
  dff s_opa_i_reg_6_ ( .Q(s_opa_i_6_), .D(opa_i[6]), .CLK(clk_i) );
  dff s_opa_i_reg_5_ ( .Q(s_opa_i_5_), .D(opa_i[5]), .CLK(clk_i) );
  dff s_opa_i_reg_4_ ( .Q(s_opa_i_4_), .D(opa_i[4]), .CLK(clk_i) );
  dff s_opa_i_reg_3_ ( .QB(n8822), .D(opa_i[3]), .CLK(clk_i) );
  dff s_opa_i_reg_2_ ( .QB(n8821), .D(opa_i[2]), .CLK(clk_i) );
  dff s_opa_i_reg_1_ ( .Q(s_opa_i_1_), .D(opa_i[1]), .CLK(clk_i) );
  dff s_opa_i_reg_0_ ( .Q(s_opa_i_0_), .D(opa_i[0]), .CLK(clk_i) );
  dff s_opb_i_reg_30_ ( .Q(s_opb_i_30_), .D(opb_i[30]), .CLK(clk_i) );
  dff s_opb_i_reg_29_ ( .Q(s_opb_i_29_), .D(opb_i[29]), .CLK(clk_i) );
  dff s_opb_i_reg_28_ ( .Q(s_opb_i_28_), .D(opb_i[28]), .CLK(clk_i) );
  dff s_opb_i_reg_27_ ( .QB(n8858), .D(opb_i[27]), .CLK(clk_i) );
  dff s_opb_i_reg_26_ ( .QB(n8857), .D(opb_i[26]), .CLK(clk_i) );
  dff s_opb_i_reg_25_ ( .Q(s_opb_i_25_), .D(opb_i[25]), .CLK(clk_i) );
  dff s_opb_i_reg_24_ ( .Q(s_opb_i_24_), .D(opb_i[24]), .CLK(clk_i) );
  dff s_opb_i_reg_23_ ( .Q(s_opb_i_23_), .D(opb_i[23]), .CLK(clk_i) );
  dff s_opb_i_reg_22_ ( .QB(n8849), .D(opb_i[22]), .CLK(clk_i) );
  dff s_opb_i_reg_21_ ( .Q(s_opb_i_21_), .D(opb_i[21]), .CLK(clk_i) );
  dff s_opb_i_reg_20_ ( .Q(s_opb_i_20_), .D(opb_i[20]), .CLK(clk_i) );
  dff s_opb_i_reg_19_ ( .QB(n8854), .D(opb_i[19]), .CLK(clk_i) );
  dff s_opb_i_reg_18_ ( .QB(n8853), .D(opb_i[18]), .CLK(clk_i) );
  dff s_opb_i_reg_17_ ( .QB(n8852), .D(opb_i[17]), .CLK(clk_i) );
  dff s_opb_i_reg_16_ ( .Q(s_opb_i_16_), .D(opb_i[16]), .CLK(clk_i) );
  dff s_opb_i_reg_15_ ( .Q(s_opb_i_15_), .D(opb_i[15]), .CLK(clk_i) );
  dff s_opb_i_reg_14_ ( .Q(s_opb_i_14_), .D(opb_i[14]), .CLK(clk_i) );
  dff s_opb_i_reg_13_ ( .QB(n8856), .D(opb_i[13]), .CLK(clk_i) );
  dff s_opb_i_reg_12_ ( .QB(n8855), .D(opb_i[12]), .CLK(clk_i) );
  dff s_opb_i_reg_11_ ( .Q(s_opb_i_11_), .D(opb_i[11]), .CLK(clk_i) );
  dff s_opb_i_reg_10_ ( .Q(s_opb_i_10_), .D(opb_i[10]), .CLK(clk_i) );
  dff s_opb_i_reg_9_ ( .QB(n8848), .D(opb_i[9]), .CLK(clk_i) );
  dff s_opb_i_reg_8_ ( .QB(n8847), .D(opb_i[8]), .CLK(clk_i) );
  dff s_opb_i_reg_7_ ( .QB(n8846), .D(opb_i[7]), .CLK(clk_i) );
  dff s_opb_i_reg_6_ ( .Q(s_opb_i_6_), .D(opb_i[6]), .CLK(clk_i) );
  dff s_opb_i_reg_5_ ( .Q(s_opb_i_5_), .D(opb_i[5]), .CLK(clk_i) );
  dff s_opb_i_reg_4_ ( .Q(s_opb_i_4_), .D(opb_i[4]), .CLK(clk_i) );
  dff s_opb_i_reg_3_ ( .QB(n8851), .D(opb_i[3]), .CLK(clk_i) );
  dff s_opb_i_reg_2_ ( .QB(n8850), .D(opb_i[2]), .CLK(clk_i) );
  dff s_opb_i_reg_1_ ( .Q(s_opb_i_1_), .D(opb_i[1]), .CLK(clk_i) );
  dff s_opb_i_reg_0_ ( .Q(s_opb_i_0_), .D(opb_i[0]), .CLK(clk_i) );
  dff s_sign_i_reg ( .Q(s_sign_i), .D(sign_i), .CLK(clk_i) );
  dff ine_o_reg ( .Q(ine_o), .D(s_ine_o), .CLK(clk_i) );
  dff s_shl1_reg_0_ ( .Q(s_shl1_0_), .D(v_shl433_0_), .CLK(clk_i) );
  dff s_fraco2_reg_22_ ( .Q(s_fraco2_22_), .D(s_fraco23289_22_), .CLK(clk_i)
         );
  dff s_fraco2_reg_21_ ( .QB(n8803), .D(s_fraco23289_21_), .CLK(clk_i) );
  dff s_fraco2_reg_20_ ( .QB(n8804), .D(s_fraco23289_20_), .CLK(clk_i) );
  dff s_fraco2_reg_19_ ( .QB(n8806), .D(s_fraco23289_19_), .CLK(clk_i) );
  dff s_fraco2_reg_18_ ( .QB(n8807), .D(s_fraco23289_18_), .CLK(clk_i) );
  dff s_fraco2_reg_17_ ( .QB(n8808), .D(s_fraco23289_17_), .CLK(clk_i) );
  dff s_fraco2_reg_16_ ( .QB(n8809), .D(s_fraco23289_16_), .CLK(clk_i) );
  dff s_fraco2_reg_15_ ( .QB(n8810), .D(s_fraco23289_15_), .CLK(clk_i) );
  dff s_fraco2_reg_14_ ( .QB(n8811), .D(s_fraco23289_14_), .CLK(clk_i) );
  dff s_fraco2_reg_13_ ( .QB(n8812), .D(s_fraco23289_13_), .CLK(clk_i) );
  dff s_fraco2_reg_12_ ( .QB(n8813), .D(s_fraco23289_12_), .CLK(clk_i) );
  dff s_fraco2_reg_11_ ( .QB(n8814), .D(s_fraco23289_11_), .CLK(clk_i) );
  dff s_fraco2_reg_10_ ( .QB(n8815), .D(s_fraco23289_10_), .CLK(clk_i) );
  dff s_fraco2_reg_9_ ( .QB(n8795), .D(s_fraco23289_9_), .CLK(clk_i) );
  dff s_fraco2_reg_8_ ( .QB(n8796), .D(s_fraco23289_8_), .CLK(clk_i) );
  dff s_fraco2_reg_7_ ( .QB(n8797), .D(s_fraco23289_7_), .CLK(clk_i) );
  dff s_fraco2_reg_6_ ( .QB(n8798), .D(s_fraco23289_6_), .CLK(clk_i) );
  dff s_fraco2_reg_5_ ( .QB(n8799), .D(s_fraco23289_5_), .CLK(clk_i) );
  dff s_fraco2_reg_4_ ( .QB(n8800), .D(s_fraco23289_4_), .CLK(clk_i) );
  dff s_fraco2_reg_3_ ( .QB(n8801), .D(s_fraco23289_3_), .CLK(clk_i) );
  dff s_fraco2_reg_2_ ( .QB(n8802), .D(s_fraco23289_2_), .CLK(clk_i) );
  dff s_fraco2_reg_1_ ( .QB(n8805), .D(s_fraco23289_1_), .CLK(clk_i) );
  dff s_fraco2_reg_0_ ( .QB(n8816), .D(s_fraco23289_0_), .CLK(clk_i) );
  xor2 U1535 ( .Y(n5150), .A0(n5539), .A1(n8746) );
  inv01 U1536 ( .Y(n5151), .A(n5150) );
  xor2 U1537 ( .Y(n5152), .A0(n5534), .A1(n8900) );
  inv01 U1538 ( .Y(n5153), .A(n5152) );
  inv01 U1539 ( .Y(n5154), .A(n8775) );
  inv02 U1540 ( .Y(n8775), .A(n8776) );
  inv01 U1541 ( .Y(n5155), .A(n8779) );
  inv01 U1542 ( .Y(n5156), .A(n8777) );
  xor2 U1543 ( .Y(n5157), .A0(n7964), .A1(n5605) );
  inv01 U1544 ( .Y(n5158), .A(n5157) );
  inv01 U1545 ( .Y(n5159), .A(n8767) );
  nand02 U1546 ( .Y(n5160), .A0(s_shl1_1_), .A1(s_shl1_0_) );
  inv02 U1547 ( .Y(n5161), .A(n5160) );
  inv02 U1548 ( .Y(n8416), .A(n8761) );
  or02 U1549 ( .Y(n5162), .A0(n8417), .A1(n8418) );
  inv01 U1550 ( .Y(n5163), .A(n5162) );
  inv02 U1551 ( .Y(n8330), .A(n8514) );
  xor2 U1552 ( .Y(n5164), .A0(n8414), .A1(n8415) );
  inv01 U1553 ( .Y(n5165), .A(n5164) );
  ao22 U1554 ( .Y(n5166), .A0(n8365), .A1(s_qutnt_i[4]), .B0(n8374), .B1(
        s_qutnt_i[7]) );
  inv01 U1555 ( .Y(n5167), .A(n5166) );
  inv02 U1556 ( .Y(n5490), .A(n8609) );
  inv01 U1557 ( .Y(n5168), .A(n8397) );
  inv02 U1558 ( .Y(n8397), .A(n8398) );
  inv01 U1559 ( .Y(n5169), .A(n8403) );
  or02 U1560 ( .Y(n5170), .A0(n8167), .A1(n8339) );
  inv01 U1561 ( .Y(n5171), .A(n5170) );
  or02 U1562 ( .Y(n5172), .A0(n7732), .A1(n8341) );
  inv01 U1563 ( .Y(n5173), .A(n5172) );
  or02 U1564 ( .Y(n5174), .A0(n8071), .A1(n8341) );
  inv01 U1565 ( .Y(n5175), .A(n5174) );
  ao22 U1566 ( .Y(n5176), .A0(n8367), .A1(s_qutnt_i[3]), .B0(n8372), .B1(
        s_qutnt_i[6]) );
  inv01 U1567 ( .Y(n5177), .A(n5176) );
  inv01 U1568 ( .Y(n5178), .A(n8773) );
  ao22 U1569 ( .Y(n5179), .A0(n8352), .A1(n8578), .B0(n8359), .B1(n8654) );
  inv01 U1570 ( .Y(n5180), .A(n5179) );
  or02 U1571 ( .Y(n5181), .A0(n8414), .A1(n8339) );
  inv01 U1572 ( .Y(n5182), .A(n5181) );
  or02 U1573 ( .Y(n5183), .A0(n8399), .A1(n8341) );
  inv01 U1574 ( .Y(n5184), .A(n5183) );
  buf02 U1575 ( .Y(n5185), .A(n8748) );
  or02 U1576 ( .Y(n5186), .A0(n8362), .A1(n8814) );
  inv01 U1577 ( .Y(n5187), .A(n5186) );
  or02 U1578 ( .Y(n5188), .A0(n8362), .A1(n8808) );
  inv01 U1579 ( .Y(n5189), .A(n5188) );
  or02 U1580 ( .Y(n5190), .A0(n8362), .A1(n8802) );
  inv01 U1581 ( .Y(n5191), .A(n5190) );
  or02 U1582 ( .Y(n5192), .A0(n8362), .A1(n8807) );
  inv01 U1583 ( .Y(n5193), .A(n5192) );
  ao22 U1584 ( .Y(n5194), .A0(n8369), .A1(s_qutnt_i[18]), .B0(n8361), .B1(
        s_qutnt_i[19]) );
  inv01 U1585 ( .Y(n5195), .A(n5194) );
  or02 U1586 ( .Y(n5196), .A0(n8362), .A1(n8804) );
  inv01 U1587 ( .Y(n5197), .A(n5196) );
  or02 U1588 ( .Y(n5198), .A0(n8362), .A1(n8798) );
  inv01 U1589 ( .Y(n5199), .A(n5198) );
  or02 U1590 ( .Y(n5200), .A0(n8362), .A1(n8800) );
  inv01 U1591 ( .Y(n5201), .A(n5200) );
  or02 U1592 ( .Y(n5202), .A0(n8362), .A1(n8805) );
  inv01 U1593 ( .Y(n5203), .A(n5202) );
  or02 U1594 ( .Y(n5204), .A0(n8362), .A1(n8796) );
  inv01 U1595 ( .Y(n5205), .A(n5204) );
  or02 U1596 ( .Y(n5206), .A0(n8362), .A1(n8812) );
  inv01 U1597 ( .Y(n5207), .A(n5206) );
  or02 U1598 ( .Y(n5208), .A0(n8362), .A1(n8813) );
  inv01 U1599 ( .Y(n5209), .A(n5208) );
  or02 U1600 ( .Y(n5210), .A0(n8362), .A1(n8803) );
  inv01 U1601 ( .Y(n5211), .A(n5210) );
  ao22 U1602 ( .Y(n5212), .A0(s_qutnt_i[4]), .A1(n8369), .B0(n8361), .B1(
        s_qutnt_i[5]) );
  inv01 U1603 ( .Y(n5213), .A(n5212) );
  or02 U1604 ( .Y(n5214), .A0(n8362), .A1(n8809) );
  inv01 U1605 ( .Y(n5215), .A(n5214) );
  or02 U1606 ( .Y(n5216), .A0(n8362), .A1(n8795) );
  inv01 U1607 ( .Y(n5217), .A(n5216) );
  or02 U1608 ( .Y(n5218), .A0(n8362), .A1(n8797) );
  inv01 U1609 ( .Y(n5219), .A(n5218) );
  or02 U1610 ( .Y(n5220), .A0(n8362), .A1(n8806) );
  inv01 U1611 ( .Y(n5221), .A(n5220) );
  or02 U1612 ( .Y(n5222), .A0(n8362), .A1(n8815) );
  inv01 U1613 ( .Y(n5223), .A(n5222) );
  or02 U1614 ( .Y(n5224), .A0(n8362), .A1(n8810) );
  inv01 U1615 ( .Y(n5225), .A(n5224) );
  or02 U1616 ( .Y(n5226), .A0(n8362), .A1(n8811) );
  inv01 U1617 ( .Y(n5227), .A(n5226) );
  or02 U1618 ( .Y(n5228), .A0(n8362), .A1(n8816) );
  inv01 U1619 ( .Y(n5229), .A(n5228) );
  or02 U1620 ( .Y(n5230), .A0(n8362), .A1(n8799) );
  inv01 U1621 ( .Y(n5231), .A(n5230) );
  or02 U1622 ( .Y(n5232), .A0(n8362), .A1(n8801) );
  inv01 U1623 ( .Y(n5233), .A(n5232) );
  ao22 U1624 ( .Y(n5234), .A0(n____return3241_22_), .A1(n8552), .B0(
        n____return3241_23_), .B1(n8553) );
  inv01 U1625 ( .Y(n5235), .A(n5234) );
  nand02 U1626 ( .Y(n8729), .A0(n5236), .A1(n5237) );
  inv01 U1627 ( .Y(n5238), .A(s_qutnt_i[12]) );
  inv01 U1628 ( .Y(n5239), .A(s_qutnt_i[9]) );
  inv01 U1629 ( .Y(n5240), .A(n8366) );
  inv01 U1630 ( .Y(n5241), .A(n8372) );
  nand02 U1631 ( .Y(n5242), .A0(n5238), .A1(n5239) );
  nand02 U1632 ( .Y(n5243), .A0(n5238), .A1(n5240) );
  nand02 U1633 ( .Y(n5244), .A0(n5239), .A1(n5241) );
  nand02 U1634 ( .Y(n5245), .A0(n5240), .A1(n5241) );
  nand02 U1635 ( .Y(n5246), .A0(n5242), .A1(n5243) );
  inv01 U1636 ( .Y(n5236), .A(n5246) );
  nand02 U1637 ( .Y(n5247), .A0(n5244), .A1(n5245) );
  inv01 U1638 ( .Y(n5237), .A(n5247) );
  nand02 U1639 ( .Y(n8732), .A0(n5248), .A1(n5249) );
  inv01 U1640 ( .Y(n5250), .A(s_qutnt_i[24]) );
  inv01 U1641 ( .Y(n5251), .A(s_qutnt_i[23]) );
  inv01 U1642 ( .Y(n5252), .A(n8369) );
  inv01 U1643 ( .Y(n5253), .A(n8361) );
  nand02 U1644 ( .Y(n5254), .A0(n5250), .A1(n5251) );
  nand02 U1645 ( .Y(n5255), .A0(n5250), .A1(n5252) );
  nand02 U1646 ( .Y(n5256), .A0(n5251), .A1(n5253) );
  nand02 U1647 ( .Y(n5257), .A0(n5252), .A1(n5253) );
  nand02 U1648 ( .Y(n5258), .A0(n5254), .A1(n5255) );
  inv01 U1649 ( .Y(n5248), .A(n5258) );
  nand02 U1650 ( .Y(n5259), .A0(n5256), .A1(n5257) );
  inv01 U1651 ( .Y(n5249), .A(n5259) );
  ao22 U1652 ( .Y(n5260), .A0(n8369), .A1(s_qutnt_i[9]), .B0(n8361), .B1(
        s_qutnt_i[10]) );
  inv01 U1653 ( .Y(n5261), .A(n5260) );
  ao22 U1654 ( .Y(n5262), .A0(n8367), .A1(s_qutnt_i[23]), .B0(n8373), .B1(
        s_qutnt_i[26]) );
  inv01 U1655 ( .Y(n5263), .A(n5262) );
  inv02 U1656 ( .Y(n8366), .A(n8364) );
  nand02 U1657 ( .Y(n8708), .A0(n5264), .A1(n5265) );
  inv01 U1658 ( .Y(n5266), .A(s_qutnt_i[17]) );
  inv01 U1659 ( .Y(n5267), .A(s_qutnt_i[14]) );
  inv01 U1660 ( .Y(n5268), .A(n8367) );
  inv01 U1661 ( .Y(n5269), .A(n8374) );
  nand02 U1662 ( .Y(n5270), .A0(n5266), .A1(n5267) );
  nand02 U1663 ( .Y(n5271), .A0(n5266), .A1(n5268) );
  nand02 U1664 ( .Y(n5272), .A0(n5267), .A1(n5269) );
  nand02 U1665 ( .Y(n5273), .A0(n5268), .A1(n5269) );
  nand02 U1666 ( .Y(n5274), .A0(n5270), .A1(n5271) );
  inv01 U1667 ( .Y(n5264), .A(n5274) );
  nand02 U1668 ( .Y(n5275), .A0(n5272), .A1(n5273) );
  inv01 U1669 ( .Y(n5265), .A(n5275) );
  ao22 U1670 ( .Y(n5276), .A0(n8370), .A1(s_qutnt_i[14]), .B0(n8361), .B1(
        s_qutnt_i[15]) );
  inv01 U1671 ( .Y(n5277), .A(n5276) );
  ao22 U1672 ( .Y(n5278), .A0(n8369), .A1(s_qutnt_i[21]), .B0(n8361), .B1(
        s_qutnt_i[22]) );
  inv01 U1673 ( .Y(n5279), .A(n5278) );
  nand02 U1674 ( .Y(n8701), .A0(n5280), .A1(n5281) );
  inv01 U1675 ( .Y(n5282), .A(s_qutnt_i[18]) );
  inv01 U1676 ( .Y(n5283), .A(s_qutnt_i[15]) );
  inv01 U1677 ( .Y(n5284), .A(n8365) );
  inv01 U1678 ( .Y(n5285), .A(n8373) );
  nand02 U1679 ( .Y(n5286), .A0(n5282), .A1(n5283) );
  nand02 U1680 ( .Y(n5287), .A0(n5282), .A1(n5284) );
  nand02 U1681 ( .Y(n5288), .A0(n5283), .A1(n5285) );
  nand02 U1682 ( .Y(n5289), .A0(n5284), .A1(n5285) );
  nand02 U1683 ( .Y(n5290), .A0(n5286), .A1(n5287) );
  inv01 U1684 ( .Y(n5280), .A(n5290) );
  nand02 U1685 ( .Y(n5291), .A0(n5288), .A1(n5289) );
  inv01 U1686 ( .Y(n5281), .A(n5291) );
  ao22 U1687 ( .Y(n5292), .A0(n8370), .A1(s_qutnt_i[15]), .B0(n8361), .B1(
        s_qutnt_i[16]) );
  inv01 U1688 ( .Y(n5293), .A(n5292) );
  nand02 U1689 ( .Y(n8743), .A0(n5294), .A1(n5295) );
  inv01 U1690 ( .Y(n5296), .A(s_qutnt_i[17]) );
  inv01 U1691 ( .Y(n5297), .A(s_qutnt_i[16]) );
  inv01 U1692 ( .Y(n5298), .A(n8370) );
  inv01 U1693 ( .Y(n5299), .A(n8361) );
  nand02 U1694 ( .Y(n5300), .A0(n5296), .A1(n5297) );
  nand02 U1695 ( .Y(n5301), .A0(n5296), .A1(n5298) );
  nand02 U1696 ( .Y(n5302), .A0(n5297), .A1(n5299) );
  nand02 U1697 ( .Y(n5303), .A0(n5298), .A1(n5299) );
  nand02 U1698 ( .Y(n5304), .A0(n5300), .A1(n5301) );
  inv01 U1699 ( .Y(n5294), .A(n5304) );
  nand02 U1700 ( .Y(n5305), .A0(n5302), .A1(n5303) );
  inv01 U1701 ( .Y(n5295), .A(n5305) );
  ao22 U1702 ( .Y(n5306), .A0(n8367), .A1(s_qutnt_i[16]), .B0(n8373), .B1(
        s_qutnt_i[19]) );
  inv01 U1703 ( .Y(n5307), .A(n5306) );
  ao22 U1704 ( .Y(n5308), .A0(n8370), .A1(s_qutnt_i[12]), .B0(n8361), .B1(
        s_qutnt_i[13]) );
  inv01 U1705 ( .Y(n5309), .A(n5308) );
  nand02 U1706 ( .Y(n8737), .A0(n5310), .A1(n5311) );
  inv01 U1707 ( .Y(n5312), .A(s_qutnt_i[10]) );
  inv01 U1708 ( .Y(n5313), .A(s_qutnt_i[7]) );
  inv01 U1709 ( .Y(n5314), .A(n8366) );
  inv01 U1710 ( .Y(n5315), .A(n8374) );
  nand02 U1711 ( .Y(n5316), .A0(n5312), .A1(n5313) );
  nand02 U1712 ( .Y(n5317), .A0(n5312), .A1(n5314) );
  nand02 U1713 ( .Y(n5318), .A0(n5313), .A1(n5315) );
  nand02 U1714 ( .Y(n5319), .A0(n5314), .A1(n5315) );
  nand02 U1715 ( .Y(n5320), .A0(n5316), .A1(n5317) );
  inv01 U1716 ( .Y(n5310), .A(n5320) );
  nand02 U1717 ( .Y(n5321), .A0(n5318), .A1(n5319) );
  inv01 U1718 ( .Y(n5311), .A(n5321) );
  ao22 U1719 ( .Y(n5322), .A0(n8369), .A1(s_qutnt_i[7]), .B0(n8361), .B1(
        s_qutnt_i[8]) );
  inv01 U1720 ( .Y(n5323), .A(n5322) );
  ao22 U1721 ( .Y(n5324), .A0(n8367), .A1(s_qutnt_i[22]), .B0(n8373), .B1(
        s_qutnt_i[25]) );
  inv01 U1722 ( .Y(n5325), .A(n5324) );
  ao22 U1723 ( .Y(n5326), .A0(n8366), .A1(s_qutnt_i[12]), .B0(n8374), .B1(
        s_qutnt_i[15]) );
  inv01 U1724 ( .Y(n5327), .A(n5326) );
  nand02 U1725 ( .Y(n8685), .A0(n5328), .A1(n5329) );
  inv01 U1726 ( .Y(n5330), .A(s_qutnt_i[21]) );
  inv01 U1727 ( .Y(n5331), .A(s_qutnt_i[18]) );
  inv01 U1728 ( .Y(n5332), .A(n8365) );
  inv01 U1729 ( .Y(n5333), .A(n8373) );
  nand02 U1730 ( .Y(n5334), .A0(n5330), .A1(n5331) );
  nand02 U1731 ( .Y(n5335), .A0(n5330), .A1(n5332) );
  nand02 U1732 ( .Y(n5336), .A0(n5331), .A1(n5333) );
  nand02 U1733 ( .Y(n5337), .A0(n5332), .A1(n5333) );
  nand02 U1734 ( .Y(n5338), .A0(n5334), .A1(n5335) );
  inv01 U1735 ( .Y(n5328), .A(n5338) );
  nand02 U1736 ( .Y(n5339), .A0(n5336), .A1(n5337) );
  inv01 U1737 ( .Y(n5329), .A(n5339) );
  ao22 U1738 ( .Y(n5340), .A0(n8370), .A1(s_qutnt_i[22]), .B0(n8361), .B1(
        s_qutnt_i[23]) );
  inv01 U1739 ( .Y(n5341), .A(n5340) );
  ao22 U1740 ( .Y(n5342), .A0(n8365), .A1(s_qutnt_i[21]), .B0(n8373), .B1(
        s_qutnt_i[24]) );
  inv01 U1741 ( .Y(n5343), .A(n5342) );
  inv01 U1742 ( .Y(n8731), .A(n5344) );
  nor02 U1743 ( .Y(n5345), .A0(n8366), .A1(s_qutnt_i[3]) );
  nor02 U1744 ( .Y(n5346), .A0(s_qutnt_i[0]), .A1(s_qutnt_i[3]) );
  nor02 U1745 ( .Y(n5347), .A0(n8366), .A1(n8374) );
  nor02 U1746 ( .Y(n5348), .A0(s_qutnt_i[0]), .A1(n8374) );
  nor02 U1747 ( .Y(n5344), .A0(n5349), .A1(n5350) );
  nor02 U1748 ( .Y(n5351), .A0(n5345), .A1(n5346) );
  inv01 U1749 ( .Y(n5349), .A(n5351) );
  nor02 U1750 ( .Y(n5352), .A0(n5347), .A1(n5348) );
  inv01 U1751 ( .Y(n5350), .A(n5352) );
  nand02 U1752 ( .Y(n8728), .A0(n5353), .A1(n5354) );
  inv01 U1753 ( .Y(n5355), .A(s_qutnt_i[4]) );
  inv01 U1754 ( .Y(n5356), .A(n8366) );
  inv01 U1755 ( .Y(n5357), .A(s_qutnt_i[1]) );
  inv01 U1756 ( .Y(n5358), .A(n8374) );
  nand02 U1757 ( .Y(n5359), .A0(n5355), .A1(n5356) );
  nand02 U1758 ( .Y(n5360), .A0(n5355), .A1(n5357) );
  nand02 U1759 ( .Y(n5361), .A0(n5356), .A1(n5358) );
  nand02 U1760 ( .Y(n5362), .A0(n5357), .A1(n5358) );
  nand02 U1761 ( .Y(n5363), .A0(n5359), .A1(n5360) );
  inv01 U1762 ( .Y(n5353), .A(n5363) );
  nand02 U1763 ( .Y(n5364), .A0(n5361), .A1(n5362) );
  inv01 U1764 ( .Y(n5354), .A(n5364) );
  ao22 U1765 ( .Y(n5365), .A0(s_qutnt_i[2]), .A1(n8366), .B0(n8374), .B1(
        s_qutnt_i[5]) );
  inv01 U1766 ( .Y(n5366), .A(n5365) );
  nand02 U1767 ( .Y(n8724), .A0(n5367), .A1(n5368) );
  inv01 U1768 ( .Y(n5369), .A(s_qutnt_i[13]) );
  inv01 U1769 ( .Y(n5370), .A(s_qutnt_i[10]) );
  inv01 U1770 ( .Y(n5371), .A(n8366) );
  inv01 U1771 ( .Y(n5372), .A(n8372) );
  nand02 U1772 ( .Y(n5373), .A0(n5369), .A1(n5370) );
  nand02 U1773 ( .Y(n5374), .A0(n5369), .A1(n5371) );
  nand02 U1774 ( .Y(n5375), .A0(n5370), .A1(n5372) );
  nand02 U1775 ( .Y(n5376), .A0(n5371), .A1(n5372) );
  nand02 U1776 ( .Y(n5377), .A0(n5373), .A1(n5374) );
  inv01 U1777 ( .Y(n5367), .A(n5377) );
  nand02 U1778 ( .Y(n5378), .A0(n5375), .A1(n5376) );
  inv01 U1779 ( .Y(n5368), .A(n5378) );
  ao22 U1780 ( .Y(n5379), .A0(n8369), .A1(s_qutnt_i[10]), .B0(n8361), .B1(
        s_qutnt_i[11]) );
  inv01 U1781 ( .Y(n5380), .A(n5379) );
  ao22 U1782 ( .Y(n5381), .A0(n8365), .A1(s_qutnt_i[19]), .B0(n8373), .B1(
        s_qutnt_i[22]) );
  inv01 U1783 ( .Y(n5382), .A(n5381) );
  ao22 U1784 ( .Y(n5383), .A0(n8369), .A1(s_qutnt_i[19]), .B0(n8361), .B1(
        s_qutnt_i[20]) );
  inv01 U1785 ( .Y(n5384), .A(n5383) );
  nand02 U1786 ( .Y(n8694), .A0(n5385), .A1(n5386) );
  inv01 U1787 ( .Y(n5387), .A(s_qutnt_i[6]) );
  inv01 U1788 ( .Y(n5388), .A(s_qutnt_i[5]) );
  inv01 U1789 ( .Y(n5389), .A(n8369) );
  inv01 U1790 ( .Y(n5390), .A(n8361) );
  nand02 U1791 ( .Y(n5391), .A0(n5387), .A1(n5388) );
  nand02 U1792 ( .Y(n5392), .A0(n5387), .A1(n5389) );
  nand02 U1793 ( .Y(n5393), .A0(n5388), .A1(n5390) );
  nand02 U1794 ( .Y(n5394), .A0(n5389), .A1(n5390) );
  nand02 U1795 ( .Y(n5395), .A0(n5391), .A1(n5392) );
  inv01 U1796 ( .Y(n5385), .A(n5395) );
  nand02 U1797 ( .Y(n5396), .A0(n5393), .A1(n5394) );
  inv01 U1798 ( .Y(n5386), .A(n5396) );
  ao22 U1799 ( .Y(n5397), .A0(n8367), .A1(s_qutnt_i[5]), .B0(n8372), .B1(
        s_qutnt_i[8]) );
  inv01 U1800 ( .Y(n5398), .A(n5397) );
  or02 U1801 ( .Y(n5399), .A0(n8395), .A1(n8340) );
  inv01 U1802 ( .Y(n5400), .A(n5399) );
  ao22 U1803 ( .Y(n5401), .A0(n8370), .A1(s_qutnt_i[11]), .B0(n8361), .B1(
        s_qutnt_i[12]) );
  inv01 U1804 ( .Y(n5402), .A(n5401) );
  nand02 U1805 ( .Y(n8723), .A0(n5403), .A1(n5404) );
  inv01 U1806 ( .Y(n5405), .A(s_qutnt_i[14]) );
  inv01 U1807 ( .Y(n5406), .A(s_qutnt_i[13]) );
  inv01 U1808 ( .Y(n5407), .A(n8370) );
  inv01 U1809 ( .Y(n5408), .A(n8361) );
  nand02 U1810 ( .Y(n5409), .A0(n5405), .A1(n5406) );
  nand02 U1811 ( .Y(n5410), .A0(n5405), .A1(n5407) );
  nand02 U1812 ( .Y(n5411), .A0(n5406), .A1(n5408) );
  nand02 U1813 ( .Y(n5412), .A0(n5407), .A1(n5408) );
  nand02 U1814 ( .Y(n5413), .A0(n5409), .A1(n5410) );
  inv01 U1815 ( .Y(n5403), .A(n5413) );
  nand02 U1816 ( .Y(n5414), .A0(n5411), .A1(n5412) );
  inv01 U1817 ( .Y(n5404), .A(n5414) );
  ao22 U1818 ( .Y(n5415), .A0(n8365), .A1(s_qutnt_i[13]), .B0(n8372), .B1(
        s_qutnt_i[16]) );
  inv01 U1819 ( .Y(n5416), .A(n5415) );
  ao22 U1820 ( .Y(n5417), .A0(n8365), .A1(s_qutnt_i[11]), .B0(n8372), .B1(
        s_qutnt_i[14]) );
  inv01 U1821 ( .Y(n5418), .A(n5417) );
  buf02 U1822 ( .Y(n5419), .A(n8751) );
  buf02 U1823 ( .Y(n5420), .A(n8754) );
  buf02 U1824 ( .Y(n5421), .A(n8752) );
  buf02 U1825 ( .Y(n5422), .A(n8749) );
  nand02 U1826 ( .Y(n8671), .A0(n5423), .A1(n5424) );
  inv01 U1827 ( .Y(n5425), .A(s_qutnt_i[23]) );
  inv01 U1828 ( .Y(n5426), .A(s_qutnt_i[20]) );
  inv01 U1829 ( .Y(n5427), .A(n8365) );
  inv01 U1830 ( .Y(n5428), .A(n8373) );
  nand02 U1831 ( .Y(n5429), .A0(n5425), .A1(n5426) );
  nand02 U1832 ( .Y(n5430), .A0(n5425), .A1(n5427) );
  nand02 U1833 ( .Y(n5431), .A0(n5426), .A1(n5428) );
  nand02 U1834 ( .Y(n5432), .A0(n5427), .A1(n5428) );
  nand02 U1835 ( .Y(n5433), .A0(n5429), .A1(n5430) );
  inv01 U1836 ( .Y(n5423), .A(n5433) );
  nand02 U1837 ( .Y(n5434), .A0(n5431), .A1(n5432) );
  inv01 U1838 ( .Y(n5424), .A(n5434) );
  ao22 U1839 ( .Y(n5435), .A0(n8369), .A1(s_qutnt_i[20]), .B0(n8361), .B1(
        s_qutnt_i[21]) );
  inv01 U1840 ( .Y(n5436), .A(n5435) );
  buf02 U1841 ( .Y(n5437), .A(n8753) );
  buf02 U1842 ( .Y(n5438), .A(n8750) );
  ao22 U1843 ( .Y(n5439), .A0(n8370), .A1(s_qutnt_i[8]), .B0(n8361), .B1(
        s_qutnt_i[9]) );
  inv01 U1844 ( .Y(n5440), .A(n5439) );
  ao22 U1845 ( .Y(n5441), .A0(n8369), .A1(s_qutnt_i[17]), .B0(n8361), .B1(
        s_qutnt_i[18]) );
  inv01 U1846 ( .Y(n5442), .A(n5441) );
  ao22 U1847 ( .Y(n5443), .A0(n8367), .A1(s_qutnt_i[17]), .B0(n8372), .B1(
        s_qutnt_i[20]) );
  inv01 U1848 ( .Y(n5444), .A(n5443) );
  ao22 U1849 ( .Y(n5445), .A0(n8366), .A1(s_qutnt_i[8]), .B0(n8372), .B1(
        s_qutnt_i[11]) );
  inv01 U1850 ( .Y(n5446), .A(n5445) );
  buf02 U1851 ( .Y(n5447), .A(n8755) );
  inv01 U1852 ( .Y(n5448), .A(n8769) );
  nand02 U1853 ( .Y(n8725), .A0(n5449), .A1(n5450) );
  inv01 U1854 ( .Y(n5451), .A(s_qutnt_i[9]) );
  inv01 U1855 ( .Y(n5452), .A(s_qutnt_i[6]) );
  inv01 U1856 ( .Y(n5453), .A(n8367) );
  inv01 U1857 ( .Y(n5454), .A(n8374) );
  nand02 U1858 ( .Y(n5455), .A0(n5451), .A1(n5452) );
  nand02 U1859 ( .Y(n5456), .A0(n5451), .A1(n5453) );
  nand02 U1860 ( .Y(n5457), .A0(n5452), .A1(n5454) );
  nand02 U1861 ( .Y(n5458), .A0(n5453), .A1(n5454) );
  nand02 U1862 ( .Y(n5459), .A0(n5455), .A1(n5456) );
  inv01 U1863 ( .Y(n5449), .A(n5459) );
  nand02 U1864 ( .Y(n5460), .A0(n5457), .A1(n5458) );
  inv01 U1865 ( .Y(n5450), .A(n5460) );
  ao22 U1866 ( .Y(n5461), .A0(n8370), .A1(s_qutnt_i[6]), .B0(n8361), .B1(
        s_qutnt_i[7]) );
  inv01 U1867 ( .Y(n5462), .A(n5461) );
  ao22 U1868 ( .Y(n5463), .A0(n8361), .A1(n8553), .B0(s_shr1_1_), .B1(n8382)
         );
  inv01 U1869 ( .Y(n5464), .A(n5463) );
  or02 U1870 ( .Y(n5465), .A0(n8410), .A1(n8340) );
  inv01 U1871 ( .Y(n5466), .A(n5465) );
  buf02 U1872 ( .Y(n5467), .A(n8756) );
  ao21 U1873 ( .Y(n5468), .A0(n7947), .A1(n8520), .B0(n8521) );
  inv01 U1874 ( .Y(n5469), .A(n5468) );
  buf02 U1875 ( .Y(n5470), .A(n8727) );
  nand02 U1876 ( .Y(n8405), .A0(n5471), .A1(n5472) );
  nand02 U1877 ( .Y(n5471), .A0(s_exp_10_i_2_), .A1(n8773) );
  inv01 U1878 ( .Y(n5472), .A(n8774) );
  buf08 U1879 ( .Y(n8337), .A(n8638) );
  or02 U1880 ( .Y(n5473), .A0(n8411), .A1(n8339) );
  inv01 U1881 ( .Y(n5474), .A(n5473) );
  ao22 U1882 ( .Y(n5475), .A0(n8359), .A1(n8672), .B0(n8345), .B1(n8596) );
  inv01 U1883 ( .Y(n5476), .A(n5475) );
  ao22 U1884 ( .Y(n5477), .A0(n8359), .A1(n8674), .B0(n8343), .B1(n8592) );
  inv01 U1885 ( .Y(n5478), .A(n5477) );
  ao22 U1886 ( .Y(n5479), .A0(n8363), .A1(n8666), .B0(n8343), .B1(n8584) );
  inv01 U1887 ( .Y(n5480), .A(n5479) );
  ao22 U1888 ( .Y(n5481), .A0(n8350), .A1(n8576), .B0(n8363), .B1(n8615) );
  inv01 U1889 ( .Y(n5482), .A(n5481) );
  ao22 U1890 ( .Y(n5483), .A0(n8281), .A1(n8603), .B0(n8363), .B1(n8644) );
  inv01 U1891 ( .Y(n5484), .A(n5483) );
  ao22 U1892 ( .Y(n5485), .A0(n8363), .A1(n8650), .B0(n8678), .B1(n8613) );
  inv01 U1893 ( .Y(n5486), .A(n5485) );
  nand02 U1894 ( .Y(n8598), .A0(n5487), .A1(n5488) );
  inv01 U1895 ( .Y(n5489), .A(n8610) );
  inv01 U1896 ( .Y(n5491), .A(n8359) );
  inv01 U1897 ( .Y(n5492), .A(n8352) );
  nand02 U1898 ( .Y(n5493), .A0(n5489), .A1(n5490) );
  nand02 U1899 ( .Y(n5494), .A0(n5489), .A1(n5491) );
  nand02 U1900 ( .Y(n5495), .A0(n5490), .A1(n5492) );
  nand02 U1901 ( .Y(n5496), .A0(n5491), .A1(n5492) );
  nand02 U1902 ( .Y(n5497), .A0(n5493), .A1(n5494) );
  inv01 U1903 ( .Y(n5487), .A(n5497) );
  nand02 U1904 ( .Y(n5498), .A0(n5495), .A1(n5496) );
  inv01 U1905 ( .Y(n5488), .A(n5498) );
  ao22 U1906 ( .Y(n5499), .A0(n8337), .A1(n8609), .B0(n8359), .B1(n8677) );
  inv01 U1907 ( .Y(n5500), .A(n5499) );
  ao22 U1908 ( .Y(n5501), .A0(n8363), .A1(n8673), .B0(n8337), .B1(n8630) );
  inv01 U1909 ( .Y(n5502), .A(n5501) );
  inv01 U1910 ( .Y(n8412), .A(n5503) );
  nor02 U1911 ( .Y(n5504), .A0(n7970), .A1(n8410) );
  inv01 U1912 ( .Y(n5505), .A(n8409) );
  nor02 U1913 ( .Y(n5503), .A0(n5504), .A1(n5505) );
  nand02 U1914 ( .Y(n5506), .A0(n8490), .A1(n8507) );
  inv02 U1915 ( .Y(n5507), .A(n5506) );
  ao22 U1916 ( .Y(n5508), .A0(n8363), .A1(n8674), .B0(n8350), .B1(n8592) );
  inv01 U1917 ( .Y(n5509), .A(n5508) );
  ao22 U1918 ( .Y(n5510), .A0(n8327), .A1(n8613), .B0(n8343), .B1(n8614) );
  inv01 U1919 ( .Y(n5511), .A(n5510) );
  nand03 U1920 ( .Y(n5512), .A0(n8473), .A1(n8486), .A2(s_qutnt_i[13]) );
  inv02 U1921 ( .Y(n5513), .A(n5512) );
  nand03 U1922 ( .Y(n5514), .A0(s_qutnt_i[26]), .A1(n8479), .A2(n5595) );
  inv02 U1923 ( .Y(n5515), .A(n5514) );
  or03 U1924 ( .Y(n5516), .A0(n5538), .A1(s_round), .A2(s_fraco1_3_) );
  inv01 U1925 ( .Y(n5517), .A(n5516) );
  or03 U1926 ( .Y(n5518), .A0(n8529), .A1(n____return2916), .A2(n5563) );
  inv01 U1927 ( .Y(n5519), .A(n5518) );
  inv01 U1928 ( .Y(s_fraco1812_13_), .A(n5520) );
  inv01 U1929 ( .Y(n5521), .A(n5558) );
  inv01 U1930 ( .Y(n5522), .A(n8720) );
  inv01 U1931 ( .Y(n5523), .A(n5533) );
  inv01 U1932 ( .Y(n5524), .A(n5180) );
  nor02 U1933 ( .Y(n5520), .A0(n5525), .A1(n5526) );
  nor02 U1934 ( .Y(n5527), .A0(n5521), .A1(n5522) );
  inv01 U1935 ( .Y(n5525), .A(n5527) );
  nor02 U1936 ( .Y(n5528), .A0(n5523), .A1(n5524) );
  inv01 U1937 ( .Y(n5526), .A(n5528) );
  nand03 U1938 ( .Y(n5529), .A0(n8486), .A1(n8505), .A2(n8473) );
  inv02 U1939 ( .Y(n5530), .A(n5529) );
  inv01 U1940 ( .Y(n5531), .A(n7934) );
  ao22 U1941 ( .Y(n5532), .A0(n8363), .A1(n5555), .B0(n8345), .B1(n8581) );
  inv01 U1942 ( .Y(n5533), .A(n5532) );
  buf08 U1943 ( .Y(n5534), .A(n8764) );
  nor02 U1944 ( .Y(n8762), .A0(n8759), .A1(n5535) );
  nor02 U1945 ( .Y(n5536), .A0(n8761), .A1(n8758) );
  inv01 U1946 ( .Y(n5535), .A(n5536) );
  inv01 U1947 ( .Y(n5537), .A(n5693) );
  buf02 U1948 ( .Y(n5538), .A(n8789) );
  buf08 U1949 ( .Y(n5539), .A(n8781) );
  nand02 U1950 ( .Y(n8720), .A0(n5540), .A1(n5541) );
  inv01 U1951 ( .Y(n5542), .A(n8307) );
  inv01 U1952 ( .Y(n5543), .A(n8579) );
  inv01 U1953 ( .Y(n5544), .A(n8571) );
  inv01 U1954 ( .Y(n5545), .A(n8337) );
  nand02 U1955 ( .Y(n5546), .A0(n5542), .A1(n5543) );
  nand02 U1956 ( .Y(n5547), .A0(n5542), .A1(n5544) );
  nand02 U1957 ( .Y(n5548), .A0(n5543), .A1(n5545) );
  nand02 U1958 ( .Y(n5549), .A0(n5544), .A1(n5545) );
  nand02 U1959 ( .Y(n5550), .A0(n5546), .A1(n5547) );
  inv01 U1960 ( .Y(n5540), .A(n5550) );
  nand02 U1961 ( .Y(n5551), .A0(n5548), .A1(n5549) );
  inv01 U1962 ( .Y(n5541), .A(n5551) );
  buf02 U1963 ( .Y(n5552), .A(n8713) );
  buf02 U1964 ( .Y(n5553), .A(n8656) );
  buf02 U1965 ( .Y(n5555), .A(n8656) );
  buf02 U1966 ( .Y(n5554), .A(n8656) );
  inv01 U1967 ( .Y(n5556), .A(n8381) );
  buf08 U1968 ( .Y(n8381), .A(n8544) );
  ao22 U1969 ( .Y(n5557), .A0(n8348), .A1(n8572), .B0(n8338), .B1(n8615) );
  inv01 U1970 ( .Y(n5558), .A(n5557) );
  buf02 U1971 ( .Y(n5559), .A(n8654) );
  or02 U1972 ( .Y(n5560), .A0(n8405), .A1(n7442) );
  inv01 U1973 ( .Y(n5561), .A(n5560) );
  or03 U1974 ( .Y(n5562), .A0(n8519), .A1(n5699), .A2(n8530) );
  inv01 U1975 ( .Y(n5563), .A(n5562) );
  or03 U1976 ( .Y(n5564), .A0(n8434), .A1(n8432), .A2(n8433) );
  inv01 U1977 ( .Y(n5565), .A(n5564) );
  inv01 U1978 ( .Y(n8482), .A(n5566) );
  inv01 U1979 ( .Y(n5567), .A(n8422) );
  inv01 U1980 ( .Y(n5568), .A(n8423) );
  inv01 U1981 ( .Y(n5569), .A(n8420) );
  nand02 U1982 ( .Y(n5566), .A0(n5569), .A1(n5570) );
  nand02 U1983 ( .Y(n5571), .A0(n5567), .A1(n5568) );
  inv01 U1984 ( .Y(n5570), .A(n5571) );
  ao21 U1985 ( .Y(n5572), .A0(n8388), .A1(n8461), .B0(n8427) );
  inv01 U1986 ( .Y(n5573), .A(n5572) );
  or02 U1987 ( .Y(n5574), .A0(n8317), .A1(n8318) );
  inv02 U1988 ( .Y(n5575), .A(n5574) );
  inv01 U1989 ( .Y(s_fraco23289_22_), .A(n5576) );
  nor02 U1990 ( .Y(n5577), .A0(n8381), .A1(n8868) );
  inv01 U1991 ( .Y(n5578), .A(n5235) );
  nor02 U1992 ( .Y(n5576), .A0(n5577), .A1(n5578) );
  inv01 U1993 ( .Y(n8483), .A(n5579) );
  inv01 U1994 ( .Y(n5580), .A(n8424) );
  inv01 U1995 ( .Y(n5581), .A(n8425) );
  inv01 U1996 ( .Y(n5582), .A(n8421) );
  nand02 U1997 ( .Y(n5579), .A0(n5582), .A1(n5583) );
  nand02 U1998 ( .Y(n5584), .A0(n5580), .A1(n5581) );
  inv01 U1999 ( .Y(n5583), .A(n5584) );
  inv01 U2000 ( .Y(n8458), .A(n5585) );
  inv01 U2001 ( .Y(n5586), .A(n8427) );
  inv01 U2002 ( .Y(n5587), .A(n8428) );
  inv01 U2003 ( .Y(n5588), .A(n8389) );
  nand02 U2004 ( .Y(n5585), .A0(n5588), .A1(n5589) );
  nand02 U2005 ( .Y(n5590), .A0(n5586), .A1(n5587) );
  inv01 U2006 ( .Y(n5589), .A(n5590) );
  or03 U2007 ( .Y(n5591), .A0(n8428), .A1(n8426), .A2(n8427) );
  inv01 U2008 ( .Y(n5592), .A(n5591) );
  nand02 U2009 ( .Y(n5593), .A0(n8497), .A1(n8498) );
  inv02 U2010 ( .Y(n5594), .A(n5593) );
  buf02 U2011 ( .Y(n5595), .A(n8480) );
  buf02 U2012 ( .Y(n5596), .A(n8480) );
  buf02 U2013 ( .Y(n5597), .A(n8782) );
  inv02 U2014 ( .Y(n8399), .A(n8760) );
  inv02 U2015 ( .Y(n8400), .A(n5598) );
  inv01 U2016 ( .Y(n5599), .A(n8410) );
  inv01 U2017 ( .Y(n5600), .A(n8165) );
  inv01 U2018 ( .Y(n5601), .A(n8411) );
  nor02 U2019 ( .Y(n5598), .A0(n5601), .A1(n5602) );
  nor02 U2020 ( .Y(n5603), .A0(n5599), .A1(n5600) );
  inv01 U2021 ( .Y(n5602), .A(n5603) );
  xor2 U2022 ( .Y(n5604), .A0(n8395), .A1(n8161) );
  inv01 U2023 ( .Y(n5605), .A(n5604) );
  inv02 U2024 ( .Y(n8414), .A(n8758) );
  nand02 U2025 ( .Y(n5606), .A0(s_shl1_2_), .A1(n8619) );
  inv02 U2026 ( .Y(n5607), .A(n5606) );
  or03 U2027 ( .Y(n5608), .A0(s_opa_i_28_), .A1(s_opa_i_30_), .A2(s_opa_i_29_)
         );
  inv01 U2028 ( .Y(n5609), .A(n5608) );
  or03 U2029 ( .Y(n5610), .A0(s_opb_i_28_), .A1(s_opb_i_30_), .A2(s_opb_i_29_)
         );
  inv01 U2030 ( .Y(n5611), .A(n5610) );
  inv01 U2031 ( .Y(n8786), .A(n5612) );
  inv01 U2032 ( .Y(n5613), .A(n5517) );
  inv01 U2033 ( .Y(n5614), .A(s_rmode_i_0_) );
  inv01 U2034 ( .Y(n5615), .A(n8790) );
  nand02 U2035 ( .Y(n5612), .A0(n5615), .A1(n5616) );
  nand02 U2036 ( .Y(n5617), .A0(n5613), .A1(n5614) );
  inv01 U2037 ( .Y(n5616), .A(n5617) );
  xor2 U2038 ( .Y(n5618), .A0(s_shr1_0_), .A1(n8382) );
  inv01 U2039 ( .Y(n5619), .A(n5618) );
  inv12 U2040 ( .Y(n5965), .A(n8571) );
  inv04 U2041 ( .Y(n8571), .A(n8353) );
  inv02 U2042 ( .Y(s_expo2[6]), .A(n5438) );
  inv02 U2043 ( .Y(s_expo2[4]), .A(n5421) );
  inv02 U2044 ( .Y(s_expo2[2]), .A(n5420) );
  inv02 U2045 ( .Y(s_expo2[3]), .A(n5437) );
  inv02 U2046 ( .Y(s_expo2[5]), .A(n5419) );
  inv02 U2047 ( .Y(s_expo2[7]), .A(n5422) );
  inv02 U2048 ( .Y(s_expo2[1]), .A(n5447) );
  inv02 U2049 ( .Y(s_expo2[8]), .A(n5185) );
  xor2 U2050 ( .Y(n5620), .A0(n8399), .A1(n8400) );
  inv01 U2051 ( .Y(n5621), .A(n5620) );
  inv01 U2052 ( .Y(n8625), .A(n5622) );
  nor02 U2053 ( .Y(n5623), .A0(n8308), .A1(n8376) );
  nor02 U2054 ( .Y(n5624), .A0(n8493), .A1(n8360) );
  nor02 U2055 ( .Y(n5625), .A0(n8511), .A1(n8379) );
  nor02 U2056 ( .Y(n5622), .A0(n5625), .A1(n5626) );
  nor02 U2057 ( .Y(n5627), .A0(n5623), .A1(n5624) );
  inv01 U2058 ( .Y(n5626), .A(n5627) );
  inv01 U2059 ( .Y(n8634), .A(n5628) );
  nor02 U2060 ( .Y(n5629), .A0(n8511), .A1(n8376) );
  nor02 U2061 ( .Y(n5630), .A0(n8510), .A1(n8360) );
  nor02 U2062 ( .Y(n5631), .A0(n8493), .A1(n8380) );
  nor02 U2063 ( .Y(n5628), .A0(n5631), .A1(n5632) );
  nor02 U2064 ( .Y(n5633), .A0(n5629), .A1(n5630) );
  inv01 U2065 ( .Y(n5632), .A(n5633) );
  inv02 U2066 ( .Y(n8493), .A(s_qutnt_i[4]) );
  inv01 U2067 ( .Y(n8693), .A(n5634) );
  nor02 U2068 ( .Y(n5635), .A0(n8493), .A1(n8376) );
  nor02 U2069 ( .Y(n5636), .A0(n8492), .A1(n8360) );
  nor02 U2070 ( .Y(n5637), .A0(n8510), .A1(n8379) );
  nor02 U2071 ( .Y(n5634), .A0(n5637), .A1(n5638) );
  nor02 U2072 ( .Y(n5639), .A0(n5635), .A1(n5636) );
  inv01 U2073 ( .Y(n5638), .A(n5639) );
  inv01 U2074 ( .Y(n8741), .A(n5640) );
  nor02 U2075 ( .Y(n5641), .A0(n8510), .A1(n8376) );
  nor02 U2076 ( .Y(n5642), .A0(n8462), .A1(n8360) );
  nor02 U2077 ( .Y(n5643), .A0(n8492), .A1(n8380) );
  nor02 U2078 ( .Y(n5640), .A0(n5643), .A1(n5644) );
  nor02 U2079 ( .Y(n5645), .A0(n5641), .A1(n5642) );
  inv01 U2080 ( .Y(n5644), .A(n5645) );
  inv02 U2081 ( .Y(n8492), .A(s_qutnt_i[2]) );
  inv02 U2082 ( .Y(n8510), .A(s_qutnt_i[3]) );
  ao32 U2083 ( .Y(n5646), .A0(s_shl1_3_), .A1(n8618), .A2(n8336), .B0(n8359), 
        .B1(n8663) );
  inv01 U2084 ( .Y(n5647), .A(n5646) );
  nand02 U2085 ( .Y(n8679), .A0(n5648), .A1(n5649) );
  inv01 U2086 ( .Y(n5650), .A(n8615) );
  inv01 U2087 ( .Y(n5651), .A(n8329) );
  inv01 U2088 ( .Y(n5652), .A(n8307) );
  inv01 U2089 ( .Y(n5653), .A(n8653) );
  inv02 U2090 ( .Y(n5654), .A(n8281) );
  nand02 U2091 ( .Y(n5655), .A0(n5650), .A1(n5651) );
  nand02 U2092 ( .Y(n5656), .A0(n5650), .A1(n5652) );
  nand02 U2093 ( .Y(n5657), .A0(n5650), .A1(n5653) );
  nand02 U2094 ( .Y(n5658), .A0(n5651), .A1(n5654) );
  nand02 U2095 ( .Y(n5659), .A0(n5652), .A1(n5654) );
  nand02 U2096 ( .Y(n5660), .A0(n5653), .A1(n5654) );
  nand02 U2097 ( .Y(n5661), .A0(n5655), .A1(n5656) );
  inv01 U2098 ( .Y(n5662), .A(n5661) );
  nand02 U2099 ( .Y(n5663), .A0(n5657), .A1(n5662) );
  inv01 U2100 ( .Y(n5648), .A(n5663) );
  nand02 U2101 ( .Y(n5664), .A0(n5658), .A1(n5659) );
  inv01 U2102 ( .Y(n5665), .A(n5664) );
  nand02 U2103 ( .Y(n5666), .A0(n5660), .A1(n5665) );
  inv01 U2104 ( .Y(n5649), .A(n5666) );
  buf02 U2105 ( .Y(n8307), .A(n8612) );
  inv04 U2106 ( .Y(n8281), .A(n8280) );
  nand02 U2107 ( .Y(n8599), .A0(n5667), .A1(n5668) );
  inv01 U2108 ( .Y(n5669), .A(n8607) );
  inv01 U2109 ( .Y(n5670), .A(n8327) );
  inv01 U2110 ( .Y(n5671), .A(n8606) );
  inv01 U2111 ( .Y(n5672), .A(n8605) );
  inv02 U2112 ( .Y(n5673), .A(n8345) );
  nand02 U2113 ( .Y(n5674), .A0(n5669), .A1(n5670) );
  nand02 U2114 ( .Y(n5675), .A0(n5669), .A1(n5671) );
  nand02 U2115 ( .Y(n5676), .A0(n5669), .A1(n5672) );
  nand02 U2116 ( .Y(n5677), .A0(n5670), .A1(n5673) );
  nand02 U2117 ( .Y(n5678), .A0(n5671), .A1(n5673) );
  nand02 U2118 ( .Y(n5679), .A0(n5672), .A1(n5673) );
  nand02 U2119 ( .Y(n5680), .A0(n5674), .A1(n5675) );
  inv01 U2120 ( .Y(n5681), .A(n5680) );
  nand02 U2121 ( .Y(n5682), .A0(n5676), .A1(n5681) );
  inv01 U2122 ( .Y(n5667), .A(n5682) );
  nand02 U2123 ( .Y(n5683), .A0(n5677), .A1(n5678) );
  inv01 U2124 ( .Y(n5684), .A(n5683) );
  nand02 U2125 ( .Y(n5685), .A0(n5679), .A1(n5684) );
  inv01 U2126 ( .Y(n5668), .A(n5685) );
  ao32 U2127 ( .Y(n5686), .A0(n8678), .A1(n8605), .A2(s_shr1_3_), .B0(n8363), 
        .B1(n8637) );
  inv01 U2128 ( .Y(n5687), .A(n5686) );
  nand02 U2129 ( .Y(n5688), .A0(n8279), .A1(n8509) );
  inv02 U2130 ( .Y(n5689), .A(n5688) );
  nand02 U2131 ( .Y(n5690), .A0(n8476), .A1(n8501) );
  inv02 U2132 ( .Y(n5691), .A(n5690) );
  inv01 U2133 ( .Y(s_ine_o), .A(n5692) );
  inv01 U2134 ( .Y(n5693), .A(n8516) );
  inv01 U2135 ( .Y(n5694), .A(n8517) );
  inv01 U2136 ( .Y(n5695), .A(n5519) );
  nand02 U2137 ( .Y(n5692), .A0(n5695), .A1(n5696) );
  nand02 U2138 ( .Y(n5697), .A0(n5693), .A1(n5694) );
  inv01 U2139 ( .Y(n5696), .A(n5697) );
  ao21 U2140 ( .Y(n5698), .A0(n8531), .A1(n8532), .B0(n8533) );
  inv01 U2141 ( .Y(n5699), .A(n5698) );
  inv01 U2142 ( .Y(s_fraco23289_1_), .A(n5700) );
  nor02 U2143 ( .Y(n5701), .A0(n8381), .A1(n8871) );
  nor02 U2144 ( .Y(n5702), .A0(n8375), .A1(n8557) );
  nor02 U2145 ( .Y(n5703), .A0(n8382), .A1(n8551) );
  nor02 U2146 ( .Y(n5700), .A0(n5703), .A1(n5704) );
  nor02 U2147 ( .Y(n5705), .A0(n5701), .A1(n5702) );
  inv01 U2148 ( .Y(n5704), .A(n5705) );
  inv01 U2149 ( .Y(s_fraco23289_19_), .A(n5706) );
  nor02 U2150 ( .Y(n5707), .A0(n8381), .A1(n8872) );
  nor02 U2151 ( .Y(n5708), .A0(n8375), .A1(n8558) );
  nor02 U2152 ( .Y(n5709), .A0(n8382), .A1(n8556) );
  nor02 U2153 ( .Y(n5706), .A0(n5709), .A1(n5710) );
  nor02 U2154 ( .Y(n5711), .A0(n5707), .A1(n5708) );
  inv01 U2155 ( .Y(n5710), .A(n5711) );
  nand02 U2156 ( .Y(s_fraco23289_11_), .A0(n5712), .A1(n5713) );
  inv01 U2157 ( .Y(n5714), .A(n8880) );
  inv01 U2158 ( .Y(n5715), .A(n8381) );
  inv01 U2159 ( .Y(n5716), .A(n8566) );
  inv01 U2160 ( .Y(n5717), .A(n8375) );
  inv01 U2161 ( .Y(n5718), .A(n8565) );
  inv01 U2162 ( .Y(n5719), .A(n8382) );
  nand02 U2163 ( .Y(n5720), .A0(n5714), .A1(n5715) );
  nand02 U2164 ( .Y(n5721), .A0(n5716), .A1(n5717) );
  nand02 U2165 ( .Y(n5712), .A0(n5718), .A1(n5719) );
  nand02 U2166 ( .Y(n5722), .A0(n5720), .A1(n5721) );
  inv01 U2167 ( .Y(n5713), .A(n5722) );
  nand02 U2168 ( .Y(s_fraco23289_17_), .A0(n5723), .A1(n5724) );
  inv01 U2169 ( .Y(n5725), .A(n8874) );
  inv01 U2170 ( .Y(n5726), .A(n8381) );
  inv01 U2171 ( .Y(n5727), .A(n8560) );
  inv01 U2172 ( .Y(n5728), .A(n8375) );
  inv01 U2173 ( .Y(n5729), .A(n8559) );
  inv01 U2174 ( .Y(n5730), .A(n8382) );
  nand02 U2175 ( .Y(n5731), .A0(n5725), .A1(n5726) );
  nand02 U2176 ( .Y(n5732), .A0(n5727), .A1(n5728) );
  nand02 U2177 ( .Y(n5723), .A0(n5729), .A1(n5730) );
  nand02 U2178 ( .Y(n5733), .A0(n5731), .A1(n5732) );
  inv01 U2179 ( .Y(n5724), .A(n5733) );
  inv01 U2180 ( .Y(s_fraco23289_21_), .A(n5734) );
  nor02 U2181 ( .Y(n5735), .A0(n8381), .A1(n8869) );
  nor02 U2182 ( .Y(n5736), .A0(n8375), .A1(n8555) );
  nor02 U2183 ( .Y(n5737), .A0(n8382), .A1(n8554) );
  nor02 U2184 ( .Y(n5734), .A0(n5737), .A1(n5738) );
  nor02 U2185 ( .Y(n5739), .A0(n5735), .A1(n5736) );
  inv01 U2186 ( .Y(n5738), .A(n5739) );
  nand02 U2187 ( .Y(s_fraco23289_4_), .A0(n5740), .A1(n5741) );
  inv01 U2188 ( .Y(n5742), .A(n8865) );
  inv01 U2189 ( .Y(n5743), .A(n8381) );
  inv01 U2190 ( .Y(n5744), .A(n8549) );
  inv01 U2191 ( .Y(n5745), .A(n8375) );
  inv01 U2192 ( .Y(n5746), .A(n8548) );
  inv01 U2193 ( .Y(n5747), .A(n8382) );
  nand02 U2194 ( .Y(n5748), .A0(n5742), .A1(n5743) );
  nand02 U2195 ( .Y(n5749), .A0(n5744), .A1(n5745) );
  nand02 U2196 ( .Y(n5740), .A0(n5746), .A1(n5747) );
  nand02 U2197 ( .Y(n5750), .A0(n5748), .A1(n5749) );
  inv01 U2198 ( .Y(n5741), .A(n5750) );
  nand02 U2199 ( .Y(s_fraco23289_10_), .A0(n5751), .A1(n5752) );
  inv01 U2200 ( .Y(n5753), .A(n8881) );
  inv01 U2201 ( .Y(n5754), .A(n8381) );
  inv01 U2202 ( .Y(n5755), .A(n8541) );
  inv01 U2203 ( .Y(n5756), .A(n8375) );
  inv01 U2204 ( .Y(n5757), .A(n8566) );
  inv01 U2205 ( .Y(n5758), .A(n8382) );
  nand02 U2206 ( .Y(n5759), .A0(n5753), .A1(n5754) );
  nand02 U2207 ( .Y(n5760), .A0(n5755), .A1(n5756) );
  nand02 U2208 ( .Y(n5751), .A0(n5757), .A1(n5758) );
  nand02 U2209 ( .Y(n5761), .A0(n5759), .A1(n5760) );
  inv01 U2210 ( .Y(n5752), .A(n5761) );
  inv01 U2211 ( .Y(s_fraco23289_20_), .A(n5762) );
  nor02 U2212 ( .Y(n5763), .A0(n8381), .A1(n8870) );
  nor02 U2213 ( .Y(n5764), .A0(n8375), .A1(n8556) );
  nor02 U2214 ( .Y(n5765), .A0(n8382), .A1(n8555) );
  nor02 U2215 ( .Y(n5762), .A0(n5765), .A1(n5766) );
  nor02 U2216 ( .Y(n5767), .A0(n5763), .A1(n5764) );
  inv01 U2217 ( .Y(n5766), .A(n5767) );
  nand02 U2218 ( .Y(s_fraco23289_7_), .A0(n5768), .A1(n5769) );
  inv01 U2219 ( .Y(n5770), .A(n8862) );
  inv01 U2220 ( .Y(n5771), .A(n8381) );
  inv01 U2221 ( .Y(n5772), .A(n8546) );
  inv01 U2222 ( .Y(n5773), .A(n8375) );
  inv01 U2223 ( .Y(n5774), .A(n8545) );
  inv01 U2224 ( .Y(n5775), .A(n8382) );
  nand02 U2225 ( .Y(n5776), .A0(n5770), .A1(n5771) );
  nand02 U2226 ( .Y(n5777), .A0(n5772), .A1(n5773) );
  nand02 U2227 ( .Y(n5768), .A0(n5774), .A1(n5775) );
  nand02 U2228 ( .Y(n5778), .A0(n5776), .A1(n5777) );
  inv01 U2229 ( .Y(n5769), .A(n5778) );
  inv01 U2230 ( .Y(s_fraco23289_6_), .A(n5779) );
  nor02 U2231 ( .Y(n5780), .A0(n8381), .A1(n8863) );
  nor02 U2232 ( .Y(n5781), .A0(n8375), .A1(n8547) );
  nor02 U2233 ( .Y(n5782), .A0(n8382), .A1(n8546) );
  nor02 U2234 ( .Y(n5779), .A0(n5782), .A1(n5783) );
  nor02 U2235 ( .Y(n5784), .A0(n5780), .A1(n5781) );
  inv01 U2236 ( .Y(n5783), .A(n5784) );
  nand02 U2237 ( .Y(s_fraco23289_14_), .A0(n5785), .A1(n5786) );
  inv01 U2238 ( .Y(n5787), .A(n8877) );
  inv01 U2239 ( .Y(n5788), .A(n8381) );
  inv01 U2240 ( .Y(n5789), .A(n8563) );
  inv01 U2241 ( .Y(n5790), .A(n8375) );
  inv01 U2242 ( .Y(n5791), .A(n8562) );
  inv01 U2243 ( .Y(n5792), .A(n8382) );
  nand02 U2244 ( .Y(n5793), .A0(n5787), .A1(n5788) );
  nand02 U2245 ( .Y(n5794), .A0(n5789), .A1(n5790) );
  nand02 U2246 ( .Y(n5785), .A0(n5791), .A1(n5792) );
  nand02 U2247 ( .Y(n5795), .A0(n5793), .A1(n5794) );
  inv01 U2248 ( .Y(n5786), .A(n5795) );
  inv01 U2249 ( .Y(s_fraco23289_18_), .A(n5796) );
  nor02 U2250 ( .Y(n5797), .A0(n8381), .A1(n8873) );
  nor02 U2251 ( .Y(n5798), .A0(n8375), .A1(n8559) );
  nor02 U2252 ( .Y(n5799), .A0(n8382), .A1(n8558) );
  nor02 U2253 ( .Y(n5796), .A0(n5799), .A1(n5800) );
  nor02 U2254 ( .Y(n5801), .A0(n5797), .A1(n5798) );
  inv01 U2255 ( .Y(n5800), .A(n5801) );
  inv01 U2256 ( .Y(s_fraco23289_13_), .A(n5802) );
  nor02 U2257 ( .Y(n5803), .A0(n8381), .A1(n8878) );
  nor02 U2258 ( .Y(n5804), .A0(n8375), .A1(n8564) );
  nor02 U2259 ( .Y(n5805), .A0(n8382), .A1(n8563) );
  nor02 U2260 ( .Y(n5802), .A0(n5805), .A1(n5806) );
  nor02 U2261 ( .Y(n5807), .A0(n5803), .A1(n5804) );
  inv01 U2262 ( .Y(n5806), .A(n5807) );
  inv01 U2263 ( .Y(s_fraco23289_3_), .A(n5808) );
  nor02 U2264 ( .Y(n5809), .A0(n8381), .A1(n8866) );
  nor02 U2265 ( .Y(n5810), .A0(n8375), .A1(n8550) );
  nor02 U2266 ( .Y(n5811), .A0(n8382), .A1(n8549) );
  nor02 U2267 ( .Y(n5808), .A0(n5811), .A1(n5812) );
  nor02 U2268 ( .Y(n5813), .A0(n5809), .A1(n5810) );
  inv01 U2269 ( .Y(n5812), .A(n5813) );
  nand02 U2270 ( .Y(s_fraco23289_2_), .A0(n5814), .A1(n5815) );
  inv01 U2271 ( .Y(n5816), .A(n8867) );
  inv01 U2272 ( .Y(n5817), .A(n8381) );
  inv01 U2273 ( .Y(n5818), .A(n8551) );
  inv01 U2274 ( .Y(n5819), .A(n8375) );
  inv01 U2275 ( .Y(n5820), .A(n8550) );
  inv01 U2276 ( .Y(n5821), .A(n8382) );
  nand02 U2277 ( .Y(n5822), .A0(n5816), .A1(n5817) );
  nand02 U2278 ( .Y(n5823), .A0(n5818), .A1(n5819) );
  nand02 U2279 ( .Y(n5814), .A0(n5820), .A1(n5821) );
  nand02 U2280 ( .Y(n5824), .A0(n5822), .A1(n5823) );
  inv01 U2281 ( .Y(n5815), .A(n5824) );
  nand02 U2282 ( .Y(s_fraco23289_5_), .A0(n5825), .A1(n5826) );
  inv01 U2283 ( .Y(n5827), .A(n8864) );
  inv01 U2284 ( .Y(n5828), .A(n8381) );
  inv01 U2285 ( .Y(n5829), .A(n8548) );
  inv01 U2286 ( .Y(n5830), .A(n8375) );
  inv01 U2287 ( .Y(n5831), .A(n8547) );
  inv01 U2288 ( .Y(n5832), .A(n8382) );
  nand02 U2289 ( .Y(n5833), .A0(n5827), .A1(n5828) );
  nand02 U2290 ( .Y(n5834), .A0(n5829), .A1(n5830) );
  nand02 U2291 ( .Y(n5825), .A0(n5831), .A1(n5832) );
  nand02 U2292 ( .Y(n5835), .A0(n5833), .A1(n5834) );
  inv01 U2293 ( .Y(n5826), .A(n5835) );
  inv01 U2294 ( .Y(s_fraco23289_9_), .A(n5836) );
  nor02 U2295 ( .Y(n5837), .A0(n8381), .A1(n8860) );
  nor02 U2296 ( .Y(n5838), .A0(n8375), .A1(n8543) );
  nor02 U2297 ( .Y(n5839), .A0(n8382), .A1(n8541) );
  nor02 U2298 ( .Y(n5836), .A0(n5839), .A1(n5840) );
  nor02 U2299 ( .Y(n5841), .A0(n5837), .A1(n5838) );
  inv01 U2300 ( .Y(n5840), .A(n5841) );
  nand02 U2301 ( .Y(n8613), .A0(n5842), .A1(n5843) );
  inv01 U2302 ( .Y(n5844), .A(n8328) );
  inv01 U2303 ( .Y(n5845), .A(n8683) );
  inv01 U2304 ( .Y(n5846), .A(n8322) );
  inv01 U2305 ( .Y(n5847), .A(n8681) );
  nand02 U2306 ( .Y(n5842), .A0(n5844), .A1(n5845) );
  nand02 U2307 ( .Y(n5843), .A0(n5846), .A1(n5847) );
  buf02 U2308 ( .Y(n8328), .A(n8684) );
  nand02 U2309 ( .Y(s_fraco23289_15_), .A0(n5848), .A1(n5849) );
  inv01 U2310 ( .Y(n5850), .A(n8876) );
  inv01 U2311 ( .Y(n5851), .A(n8381) );
  inv01 U2312 ( .Y(n5852), .A(n8562) );
  inv01 U2313 ( .Y(n5853), .A(n8375) );
  inv01 U2314 ( .Y(n5854), .A(n8561) );
  inv01 U2315 ( .Y(n5855), .A(n8382) );
  nand02 U2316 ( .Y(n5856), .A0(n5850), .A1(n5851) );
  nand02 U2317 ( .Y(n5857), .A0(n5852), .A1(n5853) );
  nand02 U2318 ( .Y(n5848), .A0(n5854), .A1(n5855) );
  nand02 U2319 ( .Y(n5858), .A0(n5856), .A1(n5857) );
  inv01 U2320 ( .Y(n5849), .A(n5858) );
  nand02 U2321 ( .Y(s_fraco23289_16_), .A0(n5859), .A1(n5860) );
  inv01 U2322 ( .Y(n5861), .A(n8875) );
  inv01 U2323 ( .Y(n5862), .A(n8381) );
  inv01 U2324 ( .Y(n5863), .A(n8561) );
  inv01 U2325 ( .Y(n5864), .A(n8375) );
  inv01 U2326 ( .Y(n5865), .A(n8560) );
  inv01 U2327 ( .Y(n5866), .A(n8382) );
  nand02 U2328 ( .Y(n5867), .A0(n5861), .A1(n5862) );
  nand02 U2329 ( .Y(n5868), .A0(n5863), .A1(n5864) );
  nand02 U2330 ( .Y(n5859), .A0(n5865), .A1(n5866) );
  nand02 U2331 ( .Y(n5869), .A0(n5867), .A1(n5868) );
  inv01 U2332 ( .Y(n5860), .A(n5869) );
  inv01 U2333 ( .Y(s_fraco23289_12_), .A(n5870) );
  nor02 U2334 ( .Y(n5871), .A0(n8381), .A1(n8879) );
  nor02 U2335 ( .Y(n5872), .A0(n8375), .A1(n8565) );
  nor02 U2336 ( .Y(n5873), .A0(n8382), .A1(n8564) );
  nor02 U2337 ( .Y(n5870), .A0(n5873), .A1(n5874) );
  nor02 U2338 ( .Y(n5875), .A0(n5871), .A1(n5872) );
  inv01 U2339 ( .Y(n5874), .A(n5875) );
  inv02 U2340 ( .Y(n8561), .A(n____return3241_16_) );
  nand02 U2341 ( .Y(n8408), .A0(n5876), .A1(n5877) );
  inv01 U2342 ( .Y(n5878), .A(n8411) );
  inv01 U2343 ( .Y(n5879), .A(n8405) );
  inv01 U2344 ( .Y(n5880), .A(n8406) );
  inv01 U2345 ( .Y(n5881), .A(n8410) );
  nand02 U2346 ( .Y(n5882), .A0(n5878), .A1(n5879) );
  nand02 U2347 ( .Y(n5883), .A0(n5878), .A1(n5880) );
  nand02 U2348 ( .Y(n5884), .A0(n5879), .A1(n5881) );
  nand02 U2349 ( .Y(n5885), .A0(n5880), .A1(n5881) );
  nand02 U2350 ( .Y(n5886), .A0(n5882), .A1(n5883) );
  inv01 U2351 ( .Y(n5876), .A(n5886) );
  nand02 U2352 ( .Y(n5887), .A0(n5884), .A1(n5885) );
  inv01 U2353 ( .Y(n5877), .A(n5887) );
  inv01 U2354 ( .Y(s_fraco23289_8_), .A(n5888) );
  nor02 U2355 ( .Y(n5889), .A0(n8381), .A1(n8861) );
  nor02 U2356 ( .Y(n5890), .A0(n8375), .A1(n8545) );
  nor02 U2357 ( .Y(n5891), .A0(n8543), .A1(n8382) );
  nor02 U2358 ( .Y(n5888), .A0(n5891), .A1(n5892) );
  nor02 U2359 ( .Y(n5893), .A0(n5889), .A1(n5890) );
  inv01 U2360 ( .Y(n5892), .A(n5893) );
  inv01 U2361 ( .Y(n8661), .A(n5894) );
  nor02 U2362 ( .Y(n5895), .A0(n8495), .A1(n8377) );
  nor02 U2363 ( .Y(n5896), .A0(n8496), .A1(n8386) );
  inv01 U2364 ( .Y(n5897), .A(n5343) );
  nor02 U2365 ( .Y(n5894), .A0(n5897), .A1(n5898) );
  nor02 U2366 ( .Y(n5899), .A0(n5895), .A1(n5896) );
  inv01 U2367 ( .Y(n5898), .A(n5899) );
  inv01 U2368 ( .Y(n8651), .A(n5900) );
  nor02 U2369 ( .Y(n5901), .A0(n8496), .A1(n8377) );
  nor02 U2370 ( .Y(n5902), .A0(n8494), .A1(n8387) );
  inv01 U2371 ( .Y(n5903), .A(n5325) );
  nor02 U2372 ( .Y(n5900), .A0(n5903), .A1(n5904) );
  nor02 U2373 ( .Y(n5905), .A0(n5901), .A1(n5902) );
  inv01 U2374 ( .Y(n5904), .A(n5905) );
  buf02 U2375 ( .Y(n8387), .A(n8384) );
  inv01 U2376 ( .Y(n8670), .A(n5906) );
  nor02 U2377 ( .Y(n5907), .A0(n8498), .A1(n8377) );
  nor02 U2378 ( .Y(n5908), .A0(n8495), .A1(n8385) );
  inv01 U2379 ( .Y(n5909), .A(n8671) );
  nor02 U2380 ( .Y(n5906), .A0(n5909), .A1(n5910) );
  nor02 U2381 ( .Y(n5911), .A0(n5907), .A1(n5908) );
  inv01 U2382 ( .Y(n5910), .A(n5911) );
  inv01 U2383 ( .Y(n8643), .A(n5912) );
  nor02 U2384 ( .Y(n5913), .A0(n8494), .A1(n8377) );
  nor02 U2385 ( .Y(n5914), .A0(n8479), .A1(n8385) );
  inv01 U2386 ( .Y(n5915), .A(n5263) );
  nor02 U2387 ( .Y(n5912), .A0(n5915), .A1(n5916) );
  nor02 U2388 ( .Y(n5917), .A0(n5913), .A1(n5914) );
  inv01 U2389 ( .Y(n5916), .A(n5917) );
  inv02 U2390 ( .Y(n8495), .A(s_qutnt_i[22]) );
  nand02 U2391 ( .Y(n8582), .A0(n5918), .A1(n5919) );
  inv02 U2392 ( .Y(n5920), .A(n8589) );
  inv02 U2393 ( .Y(n5921), .A(n8588) );
  inv02 U2394 ( .Y(n5922), .A(n8587) );
  inv02 U2395 ( .Y(n5923), .A(n8069) );
  inv02 U2396 ( .Y(n5924), .A(n8347) );
  nand02 U2397 ( .Y(n5925), .A0(n5922), .A1(n5926) );
  nand02 U2398 ( .Y(n5927), .A0(n5923), .A1(n5928) );
  nand02 U2399 ( .Y(n5929), .A0(n5924), .A1(n5930) );
  nand02 U2400 ( .Y(n5931), .A0(n5924), .A1(n5932) );
  nand02 U2401 ( .Y(n5933), .A0(n5965), .A1(n5934) );
  nand02 U2402 ( .Y(n5935), .A0(n5965), .A1(n5936) );
  nand02 U2403 ( .Y(n5937), .A0(n5965), .A1(n5938) );
  nand02 U2404 ( .Y(n5939), .A0(n5965), .A1(n5940) );
  nand02 U2405 ( .Y(n5941), .A0(n5920), .A1(n5921) );
  inv01 U2406 ( .Y(n5926), .A(n5941) );
  nand02 U2407 ( .Y(n5942), .A0(n5920), .A1(n5921) );
  inv01 U2408 ( .Y(n5928), .A(n5942) );
  nand02 U2409 ( .Y(n5943), .A0(n5920), .A1(n5922) );
  inv01 U2410 ( .Y(n5930), .A(n5943) );
  nand02 U2411 ( .Y(n5944), .A0(n5920), .A1(n5923) );
  inv01 U2412 ( .Y(n5932), .A(n5944) );
  nand02 U2413 ( .Y(n5945), .A0(n5921), .A1(n5922) );
  inv01 U2414 ( .Y(n5934), .A(n5945) );
  nand02 U2415 ( .Y(n5946), .A0(n5921), .A1(n5923) );
  inv01 U2416 ( .Y(n5936), .A(n5946) );
  nand02 U2417 ( .Y(n5947), .A0(n5922), .A1(n5924) );
  inv01 U2418 ( .Y(n5938), .A(n5947) );
  nand02 U2419 ( .Y(n5948), .A0(n5923), .A1(n5924) );
  inv01 U2420 ( .Y(n5940), .A(n5948) );
  nand02 U2421 ( .Y(n5949), .A0(n5925), .A1(n5927) );
  inv01 U2422 ( .Y(n5950), .A(n5949) );
  nand02 U2423 ( .Y(n5951), .A0(n5929), .A1(n5931) );
  inv01 U2424 ( .Y(n5952), .A(n5951) );
  nand02 U2425 ( .Y(n5953), .A0(n5950), .A1(n5952) );
  inv01 U2426 ( .Y(n5918), .A(n5953) );
  nand02 U2427 ( .Y(n5954), .A0(n5933), .A1(n5935) );
  inv01 U2428 ( .Y(n5955), .A(n5954) );
  nand02 U2429 ( .Y(n5956), .A0(n5937), .A1(n5939) );
  inv01 U2430 ( .Y(n5957), .A(n5956) );
  nand02 U2431 ( .Y(n5958), .A0(n5955), .A1(n5957) );
  inv01 U2432 ( .Y(n5919), .A(n5958) );
  nand02 U2433 ( .Y(n8622), .A0(n5959), .A1(n5960) );
  inv02 U2434 ( .Y(n5961), .A(n8596) );
  inv02 U2435 ( .Y(n5962), .A(n8592) );
  inv02 U2436 ( .Y(n5963), .A(n8630) );
  inv02 U2437 ( .Y(n5964), .A(n8363) );
  inv02 U2438 ( .Y(n5966), .A(n8348) );
  nand02 U2439 ( .Y(n5967), .A0(n5963), .A1(n5968) );
  nand02 U2440 ( .Y(n5969), .A0(n5964), .A1(n5970) );
  nand02 U2441 ( .Y(n5971), .A0(n5965), .A1(n5972) );
  nand02 U2442 ( .Y(n5973), .A0(n5965), .A1(n5974) );
  nand02 U2443 ( .Y(n5975), .A0(n5966), .A1(n5976) );
  nand02 U2444 ( .Y(n5977), .A0(n5966), .A1(n5978) );
  nand02 U2445 ( .Y(n5979), .A0(n5966), .A1(n5980) );
  nand02 U2446 ( .Y(n5981), .A0(n5966), .A1(n5982) );
  nand02 U2447 ( .Y(n5983), .A0(n5961), .A1(n5962) );
  inv01 U2448 ( .Y(n5968), .A(n5983) );
  nand02 U2449 ( .Y(n5984), .A0(n5961), .A1(n5962) );
  inv01 U2450 ( .Y(n5970), .A(n5984) );
  nand02 U2451 ( .Y(n5985), .A0(n5961), .A1(n5963) );
  inv01 U2452 ( .Y(n5972), .A(n5985) );
  nand02 U2453 ( .Y(n5986), .A0(n5961), .A1(n5964) );
  inv01 U2454 ( .Y(n5974), .A(n5986) );
  nand02 U2455 ( .Y(n5987), .A0(n5962), .A1(n5963) );
  inv01 U2456 ( .Y(n5976), .A(n5987) );
  nand02 U2457 ( .Y(n5988), .A0(n5962), .A1(n5964) );
  inv01 U2458 ( .Y(n5978), .A(n5988) );
  nand02 U2459 ( .Y(n5989), .A0(n5963), .A1(n5965) );
  inv01 U2460 ( .Y(n5980), .A(n5989) );
  nand02 U2461 ( .Y(n5990), .A0(n5964), .A1(n5965) );
  inv01 U2462 ( .Y(n5982), .A(n5990) );
  nand02 U2463 ( .Y(n5991), .A0(n5967), .A1(n5969) );
  inv01 U2464 ( .Y(n5992), .A(n5991) );
  nand02 U2465 ( .Y(n5993), .A0(n5971), .A1(n5973) );
  inv01 U2466 ( .Y(n5994), .A(n5993) );
  nand02 U2467 ( .Y(n5995), .A0(n5992), .A1(n5994) );
  inv01 U2468 ( .Y(n5959), .A(n5995) );
  nand02 U2469 ( .Y(n5996), .A0(n5975), .A1(n5977) );
  inv01 U2470 ( .Y(n5997), .A(n5996) );
  nand02 U2471 ( .Y(n5998), .A0(n5979), .A1(n5981) );
  inv01 U2472 ( .Y(n5999), .A(n5998) );
  nand02 U2473 ( .Y(n6000), .A0(n5997), .A1(n5999) );
  inv01 U2474 ( .Y(n5960), .A(n6000) );
  nand02 U2475 ( .Y(n8569), .A0(n6001), .A1(n6002) );
  inv02 U2476 ( .Y(n6003), .A(n8581) );
  inv02 U2477 ( .Y(n6004), .A(n8579) );
  inv02 U2478 ( .Y(n6005), .A(n8578) );
  inv02 U2479 ( .Y(n6006), .A(n8348) );
  inv02 U2480 ( .Y(n6007), .A(n8069) );
  inv02 U2481 ( .Y(n6008), .A(n8350) );
  nand02 U2482 ( .Y(n6009), .A0(n6005), .A1(n6010) );
  nand02 U2483 ( .Y(n6011), .A0(n6006), .A1(n6012) );
  nand02 U2484 ( .Y(n6013), .A0(n6007), .A1(n6014) );
  nand02 U2485 ( .Y(n6015), .A0(n6007), .A1(n6016) );
  nand02 U2486 ( .Y(n6017), .A0(n6008), .A1(n6018) );
  nand02 U2487 ( .Y(n6019), .A0(n6008), .A1(n6020) );
  nand02 U2488 ( .Y(n6021), .A0(n6008), .A1(n6022) );
  nand02 U2489 ( .Y(n6023), .A0(n6008), .A1(n6024) );
  nand02 U2490 ( .Y(n6025), .A0(n6003), .A1(n6004) );
  inv01 U2491 ( .Y(n6010), .A(n6025) );
  nand02 U2492 ( .Y(n6026), .A0(n6003), .A1(n6004) );
  inv01 U2493 ( .Y(n6012), .A(n6026) );
  nand02 U2494 ( .Y(n6027), .A0(n6003), .A1(n6005) );
  inv01 U2495 ( .Y(n6014), .A(n6027) );
  nand02 U2496 ( .Y(n6028), .A0(n6003), .A1(n6006) );
  inv01 U2497 ( .Y(n6016), .A(n6028) );
  nand02 U2498 ( .Y(n6029), .A0(n6004), .A1(n6005) );
  inv01 U2499 ( .Y(n6018), .A(n6029) );
  nand02 U2500 ( .Y(n6030), .A0(n6004), .A1(n6006) );
  inv01 U2501 ( .Y(n6020), .A(n6030) );
  nand02 U2502 ( .Y(n6031), .A0(n6005), .A1(n6007) );
  inv01 U2503 ( .Y(n6022), .A(n6031) );
  nand02 U2504 ( .Y(n6032), .A0(n6006), .A1(n6007) );
  inv01 U2505 ( .Y(n6024), .A(n6032) );
  nand02 U2506 ( .Y(n6033), .A0(n6009), .A1(n6011) );
  inv01 U2507 ( .Y(n6034), .A(n6033) );
  nand02 U2508 ( .Y(n6035), .A0(n6013), .A1(n6015) );
  inv01 U2509 ( .Y(n6036), .A(n6035) );
  nand02 U2510 ( .Y(n6037), .A0(n6034), .A1(n6036) );
  inv01 U2511 ( .Y(n6001), .A(n6037) );
  nand02 U2512 ( .Y(n6038), .A0(n6017), .A1(n6019) );
  inv01 U2513 ( .Y(n6039), .A(n6038) );
  nand02 U2514 ( .Y(n6040), .A0(n6021), .A1(n6023) );
  inv01 U2515 ( .Y(n6041), .A(n6040) );
  nand02 U2516 ( .Y(n6042), .A0(n6039), .A1(n6041) );
  inv01 U2517 ( .Y(n6002), .A(n6042) );
  nand02 U2518 ( .Y(n8590), .A0(n6043), .A1(n6044) );
  inv02 U2519 ( .Y(n6045), .A(n8597) );
  inv02 U2520 ( .Y(n6046), .A(n8596) );
  inv02 U2521 ( .Y(n6047), .A(n8595) );
  inv02 U2522 ( .Y(n6048), .A(n8069) );
  inv02 U2523 ( .Y(n6049), .A(n8351) );
  nand02 U2524 ( .Y(n6050), .A0(n6047), .A1(n6051) );
  nand02 U2525 ( .Y(n6052), .A0(n6048), .A1(n6053) );
  nand02 U2526 ( .Y(n6054), .A0(n6049), .A1(n6055) );
  nand02 U2527 ( .Y(n6056), .A0(n6049), .A1(n6057) );
  nand02 U2528 ( .Y(n6058), .A0(n5965), .A1(n6059) );
  nand02 U2529 ( .Y(n6060), .A0(n5965), .A1(n6061) );
  nand02 U2530 ( .Y(n6062), .A0(n5965), .A1(n6063) );
  nand02 U2531 ( .Y(n6064), .A0(n5965), .A1(n6065) );
  nand02 U2532 ( .Y(n6066), .A0(n6045), .A1(n6046) );
  inv01 U2533 ( .Y(n6051), .A(n6066) );
  nand02 U2534 ( .Y(n6067), .A0(n6045), .A1(n6046) );
  inv01 U2535 ( .Y(n6053), .A(n6067) );
  nand02 U2536 ( .Y(n6068), .A0(n6045), .A1(n6047) );
  inv01 U2537 ( .Y(n6055), .A(n6068) );
  nand02 U2538 ( .Y(n6069), .A0(n6045), .A1(n6048) );
  inv01 U2539 ( .Y(n6057), .A(n6069) );
  nand02 U2540 ( .Y(n6070), .A0(n6046), .A1(n6047) );
  inv01 U2541 ( .Y(n6059), .A(n6070) );
  nand02 U2542 ( .Y(n6071), .A0(n6046), .A1(n6048) );
  inv01 U2543 ( .Y(n6061), .A(n6071) );
  nand02 U2544 ( .Y(n6072), .A0(n6047), .A1(n6049) );
  inv01 U2545 ( .Y(n6063), .A(n6072) );
  nand02 U2546 ( .Y(n6073), .A0(n6048), .A1(n6049) );
  inv01 U2547 ( .Y(n6065), .A(n6073) );
  nand02 U2548 ( .Y(n6074), .A0(n6050), .A1(n6052) );
  inv01 U2549 ( .Y(n6075), .A(n6074) );
  nand02 U2550 ( .Y(n6076), .A0(n6054), .A1(n6056) );
  inv01 U2551 ( .Y(n6077), .A(n6076) );
  nand02 U2552 ( .Y(n6078), .A0(n6075), .A1(n6077) );
  inv01 U2553 ( .Y(n6043), .A(n6078) );
  nand02 U2554 ( .Y(n6079), .A0(n6058), .A1(n6060) );
  inv01 U2555 ( .Y(n6080), .A(n6079) );
  nand02 U2556 ( .Y(n6081), .A0(n6062), .A1(n6064) );
  inv01 U2557 ( .Y(n6082), .A(n6081) );
  nand02 U2558 ( .Y(n6083), .A0(n6080), .A1(n6082) );
  inv01 U2559 ( .Y(n6044), .A(n6083) );
  nand02 U2560 ( .Y(n8710), .A0(n6084), .A1(n6085) );
  inv02 U2561 ( .Y(n6086), .A(n8666) );
  inv02 U2562 ( .Y(n6087), .A(n8663) );
  inv02 U2563 ( .Y(n6088), .A(n8714) );
  inv02 U2564 ( .Y(n6089), .A(n8678) );
  inv02 U2565 ( .Y(n6090), .A(n8338) );
  inv02 U2566 ( .Y(n6091), .A(n8359) );
  nand02 U2567 ( .Y(n6092), .A0(n6088), .A1(n6093) );
  nand02 U2568 ( .Y(n6094), .A0(n6089), .A1(n6095) );
  nand02 U2569 ( .Y(n6096), .A0(n6090), .A1(n6097) );
  nand02 U2570 ( .Y(n6098), .A0(n6090), .A1(n6099) );
  nand02 U2571 ( .Y(n6100), .A0(n6091), .A1(n6101) );
  nand02 U2572 ( .Y(n6102), .A0(n6091), .A1(n6103) );
  nand02 U2573 ( .Y(n6104), .A0(n6091), .A1(n6105) );
  nand02 U2574 ( .Y(n6106), .A0(n6091), .A1(n6107) );
  nand02 U2575 ( .Y(n6108), .A0(n6086), .A1(n6087) );
  inv01 U2576 ( .Y(n6093), .A(n6108) );
  nand02 U2577 ( .Y(n6109), .A0(n6086), .A1(n6087) );
  inv01 U2578 ( .Y(n6095), .A(n6109) );
  nand02 U2579 ( .Y(n6110), .A0(n6086), .A1(n6088) );
  inv01 U2580 ( .Y(n6097), .A(n6110) );
  nand02 U2581 ( .Y(n6111), .A0(n6086), .A1(n6089) );
  inv01 U2582 ( .Y(n6099), .A(n6111) );
  nand02 U2583 ( .Y(n6112), .A0(n6087), .A1(n6088) );
  inv01 U2584 ( .Y(n6101), .A(n6112) );
  nand02 U2585 ( .Y(n6113), .A0(n6087), .A1(n6089) );
  inv01 U2586 ( .Y(n6103), .A(n6113) );
  nand02 U2587 ( .Y(n6114), .A0(n6088), .A1(n6090) );
  inv01 U2588 ( .Y(n6105), .A(n6114) );
  nand02 U2589 ( .Y(n6115), .A0(n6089), .A1(n6090) );
  inv01 U2590 ( .Y(n6107), .A(n6115) );
  nand02 U2591 ( .Y(n6116), .A0(n6092), .A1(n6094) );
  inv01 U2592 ( .Y(n6117), .A(n6116) );
  nand02 U2593 ( .Y(n6118), .A0(n6096), .A1(n6098) );
  inv01 U2594 ( .Y(n6119), .A(n6118) );
  nand02 U2595 ( .Y(n6120), .A0(n6117), .A1(n6119) );
  inv01 U2596 ( .Y(n6084), .A(n6120) );
  nand02 U2597 ( .Y(n6121), .A0(n6100), .A1(n6102) );
  inv01 U2598 ( .Y(n6122), .A(n6121) );
  nand02 U2599 ( .Y(n6123), .A0(n6104), .A1(n6106) );
  inv01 U2600 ( .Y(n6124), .A(n6123) );
  nand02 U2601 ( .Y(n6125), .A0(n6122), .A1(n6124) );
  inv01 U2602 ( .Y(n6085), .A(n6125) );
  nand02 U2603 ( .Y(n8640), .A0(n6126), .A1(n6127) );
  inv02 U2604 ( .Y(n6128), .A(n8644) );
  inv02 U2605 ( .Y(n6129), .A(n8643) );
  inv02 U2606 ( .Y(n6130), .A(n8642) );
  inv02 U2607 ( .Y(n6131), .A(n8338) );
  inv02 U2608 ( .Y(n6132), .A(n8363) );
  inv02 U2609 ( .Y(n6133), .A(n8359) );
  nand02 U2610 ( .Y(n6134), .A0(n6130), .A1(n6135) );
  nand02 U2611 ( .Y(n6136), .A0(n6131), .A1(n6137) );
  nand02 U2612 ( .Y(n6138), .A0(n6132), .A1(n6139) );
  nand02 U2613 ( .Y(n6140), .A0(n6132), .A1(n6141) );
  nand02 U2614 ( .Y(n6142), .A0(n6133), .A1(n6143) );
  nand02 U2615 ( .Y(n6144), .A0(n6133), .A1(n6145) );
  nand02 U2616 ( .Y(n6146), .A0(n6133), .A1(n6147) );
  nand02 U2617 ( .Y(n6148), .A0(n6133), .A1(n6149) );
  nand02 U2618 ( .Y(n6150), .A0(n6128), .A1(n6129) );
  inv01 U2619 ( .Y(n6135), .A(n6150) );
  nand02 U2620 ( .Y(n6151), .A0(n6128), .A1(n6129) );
  inv01 U2621 ( .Y(n6137), .A(n6151) );
  nand02 U2622 ( .Y(n6152), .A0(n6128), .A1(n6130) );
  inv01 U2623 ( .Y(n6139), .A(n6152) );
  nand02 U2624 ( .Y(n6153), .A0(n6128), .A1(n6131) );
  inv01 U2625 ( .Y(n6141), .A(n6153) );
  nand02 U2626 ( .Y(n6154), .A0(n6129), .A1(n6130) );
  inv01 U2627 ( .Y(n6143), .A(n6154) );
  nand02 U2628 ( .Y(n6155), .A0(n6129), .A1(n6131) );
  inv01 U2629 ( .Y(n6145), .A(n6155) );
  nand02 U2630 ( .Y(n6156), .A0(n6130), .A1(n6132) );
  inv01 U2631 ( .Y(n6147), .A(n6156) );
  nand02 U2632 ( .Y(n6157), .A0(n6131), .A1(n6132) );
  inv01 U2633 ( .Y(n6149), .A(n6157) );
  nand02 U2634 ( .Y(n6158), .A0(n6134), .A1(n6136) );
  inv01 U2635 ( .Y(n6159), .A(n6158) );
  nand02 U2636 ( .Y(n6160), .A0(n6138), .A1(n6140) );
  inv01 U2637 ( .Y(n6161), .A(n6160) );
  nand02 U2638 ( .Y(n6162), .A0(n6159), .A1(n6161) );
  inv01 U2639 ( .Y(n6126), .A(n6162) );
  nand02 U2640 ( .Y(n6163), .A0(n6142), .A1(n6144) );
  inv01 U2641 ( .Y(n6164), .A(n6163) );
  nand02 U2642 ( .Y(n6165), .A0(n6146), .A1(n6148) );
  inv01 U2643 ( .Y(n6166), .A(n6165) );
  nand02 U2644 ( .Y(n6167), .A0(n6164), .A1(n6166) );
  inv01 U2645 ( .Y(n6127), .A(n6167) );
  nand02 U2646 ( .Y(n8648), .A0(n6168), .A1(n6169) );
  inv02 U2647 ( .Y(n6170), .A(n8579) );
  inv02 U2648 ( .Y(n6171), .A(n8657) );
  inv02 U2649 ( .Y(n6172), .A(n5554) );
  inv02 U2650 ( .Y(n6173), .A(n8337) );
  inv02 U2651 ( .Y(n6174), .A(n8641) );
  inv02 U2652 ( .Y(n6175), .A(n8344) );
  nand02 U2653 ( .Y(n6176), .A0(n6172), .A1(n6177) );
  nand02 U2654 ( .Y(n6178), .A0(n6173), .A1(n6179) );
  nand02 U2655 ( .Y(n6180), .A0(n6174), .A1(n6181) );
  nand02 U2656 ( .Y(n6182), .A0(n6174), .A1(n6183) );
  nand02 U2657 ( .Y(n6184), .A0(n6175), .A1(n6185) );
  nand02 U2658 ( .Y(n6186), .A0(n6175), .A1(n6187) );
  nand02 U2659 ( .Y(n6188), .A0(n6175), .A1(n6189) );
  nand02 U2660 ( .Y(n6190), .A0(n6175), .A1(n6191) );
  nand02 U2661 ( .Y(n6192), .A0(n6170), .A1(n6171) );
  inv01 U2662 ( .Y(n6177), .A(n6192) );
  nand02 U2663 ( .Y(n6193), .A0(n6170), .A1(n6171) );
  inv01 U2664 ( .Y(n6179), .A(n6193) );
  nand02 U2665 ( .Y(n6194), .A0(n6170), .A1(n6172) );
  inv01 U2666 ( .Y(n6181), .A(n6194) );
  nand02 U2667 ( .Y(n6195), .A0(n6170), .A1(n6173) );
  inv01 U2668 ( .Y(n6183), .A(n6195) );
  nand02 U2669 ( .Y(n6196), .A0(n6171), .A1(n6172) );
  inv01 U2670 ( .Y(n6185), .A(n6196) );
  nand02 U2671 ( .Y(n6197), .A0(n6171), .A1(n6173) );
  inv01 U2672 ( .Y(n6187), .A(n6197) );
  nand02 U2673 ( .Y(n6198), .A0(n6172), .A1(n6174) );
  inv01 U2674 ( .Y(n6189), .A(n6198) );
  nand02 U2675 ( .Y(n6199), .A0(n6173), .A1(n6174) );
  inv01 U2676 ( .Y(n6191), .A(n6199) );
  nand02 U2677 ( .Y(n6200), .A0(n6176), .A1(n6178) );
  inv01 U2678 ( .Y(n6201), .A(n6200) );
  nand02 U2679 ( .Y(n6202), .A0(n6180), .A1(n6182) );
  inv01 U2680 ( .Y(n6203), .A(n6202) );
  nand02 U2681 ( .Y(n6204), .A0(n6201), .A1(n6203) );
  inv01 U2682 ( .Y(n6168), .A(n6204) );
  nand02 U2683 ( .Y(n6205), .A0(n6184), .A1(n6186) );
  inv01 U2684 ( .Y(n6206), .A(n6205) );
  nand02 U2685 ( .Y(n6207), .A0(n6188), .A1(n6190) );
  inv01 U2686 ( .Y(n6208), .A(n6207) );
  nand02 U2687 ( .Y(n6209), .A0(n6206), .A1(n6208) );
  inv01 U2688 ( .Y(n6169), .A(n6209) );
  nand02 U2689 ( .Y(n8706), .A0(n6210), .A1(n6211) );
  inv02 U2690 ( .Y(n6212), .A(n5553) );
  inv02 U2691 ( .Y(n6213), .A(n8615) );
  inv02 U2692 ( .Y(n6214), .A(n8654) );
  inv02 U2693 ( .Y(n6215), .A(n8338) );
  inv02 U2694 ( .Y(n6216), .A(n8337) );
  inv02 U2695 ( .Y(n6217), .A(n8359) );
  nand02 U2696 ( .Y(n6218), .A0(n6214), .A1(n6219) );
  nand02 U2697 ( .Y(n6220), .A0(n6215), .A1(n6221) );
  nand02 U2698 ( .Y(n6222), .A0(n6216), .A1(n6223) );
  nand02 U2699 ( .Y(n6224), .A0(n6216), .A1(n6225) );
  nand02 U2700 ( .Y(n6226), .A0(n6217), .A1(n6227) );
  nand02 U2701 ( .Y(n6228), .A0(n6217), .A1(n6229) );
  nand02 U2702 ( .Y(n6230), .A0(n6217), .A1(n6231) );
  nand02 U2703 ( .Y(n6232), .A0(n6217), .A1(n6233) );
  nand02 U2704 ( .Y(n6234), .A0(n6212), .A1(n6213) );
  inv01 U2705 ( .Y(n6219), .A(n6234) );
  nand02 U2706 ( .Y(n6235), .A0(n6212), .A1(n6213) );
  inv01 U2707 ( .Y(n6221), .A(n6235) );
  nand02 U2708 ( .Y(n6236), .A0(n6212), .A1(n6214) );
  inv01 U2709 ( .Y(n6223), .A(n6236) );
  nand02 U2710 ( .Y(n6237), .A0(n6212), .A1(n6215) );
  inv01 U2711 ( .Y(n6225), .A(n6237) );
  nand02 U2712 ( .Y(n6238), .A0(n6213), .A1(n6214) );
  inv01 U2713 ( .Y(n6227), .A(n6238) );
  nand02 U2714 ( .Y(n6239), .A0(n6213), .A1(n6215) );
  inv01 U2715 ( .Y(n6229), .A(n6239) );
  nand02 U2716 ( .Y(n6240), .A0(n6214), .A1(n6216) );
  inv01 U2717 ( .Y(n6231), .A(n6240) );
  nand02 U2718 ( .Y(n6241), .A0(n6215), .A1(n6216) );
  inv01 U2719 ( .Y(n6233), .A(n6241) );
  nand02 U2720 ( .Y(n6242), .A0(n6218), .A1(n6220) );
  inv01 U2721 ( .Y(n6243), .A(n6242) );
  nand02 U2722 ( .Y(n6244), .A0(n6222), .A1(n6224) );
  inv01 U2723 ( .Y(n6245), .A(n6244) );
  nand02 U2724 ( .Y(n6246), .A0(n6243), .A1(n6245) );
  inv01 U2725 ( .Y(n6210), .A(n6246) );
  nand02 U2726 ( .Y(n6247), .A0(n6226), .A1(n6228) );
  inv01 U2727 ( .Y(n6248), .A(n6247) );
  nand02 U2728 ( .Y(n6249), .A0(n6230), .A1(n6232) );
  inv01 U2729 ( .Y(n6250), .A(n6249) );
  nand02 U2730 ( .Y(n6251), .A0(n6248), .A1(n6250) );
  inv01 U2731 ( .Y(n6211), .A(n6251) );
  nand02 U2732 ( .Y(n8658), .A0(n6252), .A1(n6253) );
  inv02 U2733 ( .Y(n6254), .A(n8666) );
  inv02 U2734 ( .Y(n6255), .A(n8665) );
  inv02 U2735 ( .Y(n6256), .A(n8587) );
  inv02 U2736 ( .Y(n6257), .A(n8343) );
  inv02 U2737 ( .Y(n6258), .A(n8338) );
  inv02 U2738 ( .Y(n6259), .A(n8337) );
  nand02 U2739 ( .Y(n6260), .A0(n6256), .A1(n6261) );
  nand02 U2740 ( .Y(n6262), .A0(n6257), .A1(n6263) );
  nand02 U2741 ( .Y(n6264), .A0(n6258), .A1(n6265) );
  nand02 U2742 ( .Y(n6266), .A0(n6258), .A1(n6267) );
  nand02 U2743 ( .Y(n6268), .A0(n6259), .A1(n6269) );
  nand02 U2744 ( .Y(n6270), .A0(n6259), .A1(n6271) );
  nand02 U2745 ( .Y(n6272), .A0(n6259), .A1(n6273) );
  nand02 U2746 ( .Y(n6274), .A0(n6259), .A1(n6275) );
  nand02 U2747 ( .Y(n6276), .A0(n6254), .A1(n6255) );
  inv01 U2748 ( .Y(n6261), .A(n6276) );
  nand02 U2749 ( .Y(n6277), .A0(n6254), .A1(n6255) );
  inv01 U2750 ( .Y(n6263), .A(n6277) );
  nand02 U2751 ( .Y(n6278), .A0(n6254), .A1(n6256) );
  inv01 U2752 ( .Y(n6265), .A(n6278) );
  nand02 U2753 ( .Y(n6279), .A0(n6254), .A1(n6257) );
  inv01 U2754 ( .Y(n6267), .A(n6279) );
  nand02 U2755 ( .Y(n6280), .A0(n6255), .A1(n6256) );
  inv01 U2756 ( .Y(n6269), .A(n6280) );
  nand02 U2757 ( .Y(n6281), .A0(n6255), .A1(n6257) );
  inv01 U2758 ( .Y(n6271), .A(n6281) );
  nand02 U2759 ( .Y(n6282), .A0(n6256), .A1(n6258) );
  inv01 U2760 ( .Y(n6273), .A(n6282) );
  nand02 U2761 ( .Y(n6283), .A0(n6257), .A1(n6258) );
  inv01 U2762 ( .Y(n6275), .A(n6283) );
  nand02 U2763 ( .Y(n6284), .A0(n6260), .A1(n6262) );
  inv01 U2764 ( .Y(n6285), .A(n6284) );
  nand02 U2765 ( .Y(n6286), .A0(n6264), .A1(n6266) );
  inv01 U2766 ( .Y(n6287), .A(n6286) );
  nand02 U2767 ( .Y(n6288), .A0(n6285), .A1(n6287) );
  inv01 U2768 ( .Y(n6252), .A(n6288) );
  nand02 U2769 ( .Y(n6289), .A0(n6268), .A1(n6270) );
  inv01 U2770 ( .Y(n6290), .A(n6289) );
  nand02 U2771 ( .Y(n6291), .A0(n6272), .A1(n6274) );
  inv01 U2772 ( .Y(n6292), .A(n6291) );
  nand02 U2773 ( .Y(n6293), .A0(n6290), .A1(n6292) );
  inv01 U2774 ( .Y(n6253), .A(n6293) );
  nand02 U2775 ( .Y(n8699), .A0(n6294), .A1(n6295) );
  inv02 U2776 ( .Y(n6296), .A(n8603) );
  inv02 U2777 ( .Y(n6297), .A(n8637) );
  inv02 U2778 ( .Y(n6298), .A(n8677) );
  inv02 U2779 ( .Y(n6299), .A(n8338) );
  inv02 U2780 ( .Y(n6300), .A(n8359) );
  inv02 U2781 ( .Y(n6301), .A(n8337) );
  nand02 U2782 ( .Y(n6302), .A0(n6298), .A1(n6303) );
  nand02 U2783 ( .Y(n6304), .A0(n6299), .A1(n6305) );
  nand02 U2784 ( .Y(n6306), .A0(n6300), .A1(n6307) );
  nand02 U2785 ( .Y(n6308), .A0(n6300), .A1(n6309) );
  nand02 U2786 ( .Y(n6310), .A0(n6301), .A1(n6311) );
  nand02 U2787 ( .Y(n6312), .A0(n6301), .A1(n6313) );
  nand02 U2788 ( .Y(n6314), .A0(n6301), .A1(n6315) );
  nand02 U2789 ( .Y(n6316), .A0(n6301), .A1(n6317) );
  nand02 U2790 ( .Y(n6318), .A0(n6296), .A1(n6297) );
  inv01 U2791 ( .Y(n6303), .A(n6318) );
  nand02 U2792 ( .Y(n6319), .A0(n6296), .A1(n6297) );
  inv01 U2793 ( .Y(n6305), .A(n6319) );
  nand02 U2794 ( .Y(n6320), .A0(n6296), .A1(n6298) );
  inv01 U2795 ( .Y(n6307), .A(n6320) );
  nand02 U2796 ( .Y(n6321), .A0(n6296), .A1(n6299) );
  inv01 U2797 ( .Y(n6309), .A(n6321) );
  nand02 U2798 ( .Y(n6322), .A0(n6297), .A1(n6298) );
  inv01 U2799 ( .Y(n6311), .A(n6322) );
  nand02 U2800 ( .Y(n6323), .A0(n6297), .A1(n6299) );
  inv01 U2801 ( .Y(n6313), .A(n6323) );
  nand02 U2802 ( .Y(n6324), .A0(n6298), .A1(n6300) );
  inv01 U2803 ( .Y(n6315), .A(n6324) );
  nand02 U2804 ( .Y(n6325), .A0(n6299), .A1(n6300) );
  inv01 U2805 ( .Y(n6317), .A(n6325) );
  nand02 U2806 ( .Y(n6326), .A0(n6302), .A1(n6304) );
  inv01 U2807 ( .Y(n6327), .A(n6326) );
  nand02 U2808 ( .Y(n6328), .A0(n6306), .A1(n6308) );
  inv01 U2809 ( .Y(n6329), .A(n6328) );
  nand02 U2810 ( .Y(n6330), .A0(n6327), .A1(n6329) );
  inv01 U2811 ( .Y(n6294), .A(n6330) );
  nand02 U2812 ( .Y(n6331), .A0(n6310), .A1(n6312) );
  inv01 U2813 ( .Y(n6332), .A(n6331) );
  nand02 U2814 ( .Y(n6333), .A0(n6314), .A1(n6316) );
  inv01 U2815 ( .Y(n6334), .A(n6333) );
  nand02 U2816 ( .Y(n6335), .A0(n6332), .A1(n6334) );
  inv01 U2817 ( .Y(n6295), .A(n6335) );
  nand02 U2818 ( .Y(n8695), .A0(n6336), .A1(n6337) );
  inv02 U2819 ( .Y(n6338), .A(n8672) );
  inv02 U2820 ( .Y(n6339), .A(n8673) );
  inv02 U2821 ( .Y(n6340), .A(n8674) );
  inv02 U2822 ( .Y(n6341), .A(n8338) );
  inv02 U2823 ( .Y(n6342), .A(n8359) );
  inv02 U2824 ( .Y(n6343), .A(n8337) );
  nand02 U2825 ( .Y(n6344), .A0(n6340), .A1(n6345) );
  nand02 U2826 ( .Y(n6346), .A0(n6341), .A1(n6347) );
  nand02 U2827 ( .Y(n6348), .A0(n6342), .A1(n6349) );
  nand02 U2828 ( .Y(n6350), .A0(n6342), .A1(n6351) );
  nand02 U2829 ( .Y(n6352), .A0(n6343), .A1(n6353) );
  nand02 U2830 ( .Y(n6354), .A0(n6343), .A1(n6355) );
  nand02 U2831 ( .Y(n6356), .A0(n6343), .A1(n6357) );
  nand02 U2832 ( .Y(n6358), .A0(n6343), .A1(n6359) );
  nand02 U2833 ( .Y(n6360), .A0(n6338), .A1(n6339) );
  inv01 U2834 ( .Y(n6345), .A(n6360) );
  nand02 U2835 ( .Y(n6361), .A0(n6338), .A1(n6339) );
  inv01 U2836 ( .Y(n6347), .A(n6361) );
  nand02 U2837 ( .Y(n6362), .A0(n6338), .A1(n6340) );
  inv01 U2838 ( .Y(n6349), .A(n6362) );
  nand02 U2839 ( .Y(n6363), .A0(n6338), .A1(n6341) );
  inv01 U2840 ( .Y(n6351), .A(n6363) );
  nand02 U2841 ( .Y(n6364), .A0(n6339), .A1(n6340) );
  inv01 U2842 ( .Y(n6353), .A(n6364) );
  nand02 U2843 ( .Y(n6365), .A0(n6339), .A1(n6341) );
  inv01 U2844 ( .Y(n6355), .A(n6365) );
  nand02 U2845 ( .Y(n6366), .A0(n6340), .A1(n6342) );
  inv01 U2846 ( .Y(n6357), .A(n6366) );
  nand02 U2847 ( .Y(n6367), .A0(n6341), .A1(n6342) );
  inv01 U2848 ( .Y(n6359), .A(n6367) );
  nand02 U2849 ( .Y(n6368), .A0(n6344), .A1(n6346) );
  inv01 U2850 ( .Y(n6369), .A(n6368) );
  nand02 U2851 ( .Y(n6370), .A0(n6348), .A1(n6350) );
  inv01 U2852 ( .Y(n6371), .A(n6370) );
  nand02 U2853 ( .Y(n6372), .A0(n6369), .A1(n6371) );
  inv01 U2854 ( .Y(n6336), .A(n6372) );
  nand02 U2855 ( .Y(n6373), .A0(n6352), .A1(n6354) );
  inv01 U2856 ( .Y(n6374), .A(n6373) );
  nand02 U2857 ( .Y(n6375), .A0(n6356), .A1(n6358) );
  inv01 U2858 ( .Y(n6376), .A(n6375) );
  nand02 U2859 ( .Y(n6377), .A0(n6374), .A1(n6376) );
  inv01 U2860 ( .Y(n6337), .A(n6377) );
  nand02 U2861 ( .Y(n8686), .A0(n6378), .A1(n6379) );
  inv02 U2862 ( .Y(n6380), .A(n8663) );
  inv02 U2863 ( .Y(n6381), .A(n8665) );
  inv02 U2864 ( .Y(n6382), .A(n8666) );
  inv02 U2865 ( .Y(n6383), .A(n8338) );
  inv02 U2866 ( .Y(n6384), .A(n8359) );
  inv02 U2867 ( .Y(n6385), .A(n8337) );
  nand02 U2868 ( .Y(n6386), .A0(n6382), .A1(n6387) );
  nand02 U2869 ( .Y(n6388), .A0(n6383), .A1(n6389) );
  nand02 U2870 ( .Y(n6390), .A0(n6384), .A1(n6391) );
  nand02 U2871 ( .Y(n6392), .A0(n6384), .A1(n6393) );
  nand02 U2872 ( .Y(n6394), .A0(n6385), .A1(n6395) );
  nand02 U2873 ( .Y(n6396), .A0(n6385), .A1(n6397) );
  nand02 U2874 ( .Y(n6398), .A0(n6385), .A1(n6399) );
  nand02 U2875 ( .Y(n6400), .A0(n6385), .A1(n6401) );
  nand02 U2876 ( .Y(n6402), .A0(n6380), .A1(n6381) );
  inv01 U2877 ( .Y(n6387), .A(n6402) );
  nand02 U2878 ( .Y(n6403), .A0(n6380), .A1(n6381) );
  inv01 U2879 ( .Y(n6389), .A(n6403) );
  nand02 U2880 ( .Y(n6404), .A0(n6380), .A1(n6382) );
  inv01 U2881 ( .Y(n6391), .A(n6404) );
  nand02 U2882 ( .Y(n6405), .A0(n6380), .A1(n6383) );
  inv01 U2883 ( .Y(n6393), .A(n6405) );
  nand02 U2884 ( .Y(n6406), .A0(n6381), .A1(n6382) );
  inv01 U2885 ( .Y(n6395), .A(n6406) );
  nand02 U2886 ( .Y(n6407), .A0(n6381), .A1(n6383) );
  inv01 U2887 ( .Y(n6397), .A(n6407) );
  nand02 U2888 ( .Y(n6408), .A0(n6382), .A1(n6384) );
  inv01 U2889 ( .Y(n6399), .A(n6408) );
  nand02 U2890 ( .Y(n6409), .A0(n6383), .A1(n6384) );
  inv01 U2891 ( .Y(n6401), .A(n6409) );
  nand02 U2892 ( .Y(n6410), .A0(n6386), .A1(n6388) );
  inv01 U2893 ( .Y(n6411), .A(n6410) );
  nand02 U2894 ( .Y(n6412), .A0(n6390), .A1(n6392) );
  inv01 U2895 ( .Y(n6413), .A(n6412) );
  nand02 U2896 ( .Y(n6414), .A0(n6411), .A1(n6413) );
  inv01 U2897 ( .Y(n6378), .A(n6414) );
  nand02 U2898 ( .Y(n6415), .A0(n6394), .A1(n6396) );
  inv01 U2899 ( .Y(n6416), .A(n6415) );
  nand02 U2900 ( .Y(n6417), .A0(n6398), .A1(n6400) );
  inv01 U2901 ( .Y(n6418), .A(n6417) );
  nand02 U2902 ( .Y(n6419), .A0(n6416), .A1(n6418) );
  inv01 U2903 ( .Y(n6379), .A(n6419) );
  nand02 U2904 ( .Y(n8690), .A0(n6420), .A1(n6421) );
  inv02 U2905 ( .Y(n6422), .A(n8307) );
  inv02 U2906 ( .Y(n6423), .A(n8576) );
  inv02 U2907 ( .Y(n6424), .A(n8581) );
  inv02 U2908 ( .Y(n6425), .A(n8347) );
  inv02 U2909 ( .Y(n6426), .A(n8363) );
  nand02 U2910 ( .Y(n6427), .A0(n6424), .A1(n6428) );
  nand02 U2911 ( .Y(n6429), .A0(n5965), .A1(n6430) );
  nand02 U2912 ( .Y(n6431), .A0(n6425), .A1(n6432) );
  nand02 U2913 ( .Y(n6433), .A0(n6425), .A1(n6434) );
  nand02 U2914 ( .Y(n6435), .A0(n6426), .A1(n6436) );
  nand02 U2915 ( .Y(n6437), .A0(n6426), .A1(n6438) );
  nand02 U2916 ( .Y(n6439), .A0(n6426), .A1(n6440) );
  nand02 U2917 ( .Y(n6441), .A0(n6426), .A1(n6442) );
  nand02 U2918 ( .Y(n6443), .A0(n6422), .A1(n6423) );
  inv01 U2919 ( .Y(n6428), .A(n6443) );
  nand02 U2920 ( .Y(n6444), .A0(n6422), .A1(n6423) );
  inv01 U2921 ( .Y(n6430), .A(n6444) );
  nand02 U2922 ( .Y(n6445), .A0(n6422), .A1(n6424) );
  inv01 U2923 ( .Y(n6432), .A(n6445) );
  nand02 U2924 ( .Y(n6446), .A0(n6422), .A1(n5965) );
  inv01 U2925 ( .Y(n6434), .A(n6446) );
  nand02 U2926 ( .Y(n6447), .A0(n6423), .A1(n6424) );
  inv01 U2927 ( .Y(n6436), .A(n6447) );
  nand02 U2928 ( .Y(n6448), .A0(n6423), .A1(n5965) );
  inv01 U2929 ( .Y(n6438), .A(n6448) );
  nand02 U2930 ( .Y(n6449), .A0(n6424), .A1(n6425) );
  inv01 U2931 ( .Y(n6440), .A(n6449) );
  nand02 U2932 ( .Y(n6450), .A0(n5965), .A1(n6425) );
  inv01 U2933 ( .Y(n6442), .A(n6450) );
  nand02 U2934 ( .Y(n6451), .A0(n6427), .A1(n6429) );
  inv01 U2935 ( .Y(n6452), .A(n6451) );
  nand02 U2936 ( .Y(n6453), .A0(n6431), .A1(n6433) );
  inv01 U2937 ( .Y(n6454), .A(n6453) );
  nand02 U2938 ( .Y(n6455), .A0(n6452), .A1(n6454) );
  inv01 U2939 ( .Y(n6420), .A(n6455) );
  nand02 U2940 ( .Y(n6456), .A0(n6435), .A1(n6437) );
  inv01 U2941 ( .Y(n6457), .A(n6456) );
  nand02 U2942 ( .Y(n6458), .A0(n6439), .A1(n6441) );
  inv01 U2943 ( .Y(n6459), .A(n6458) );
  nand02 U2944 ( .Y(n6460), .A0(n6457), .A1(n6459) );
  inv01 U2945 ( .Y(n6421), .A(n6460) );
  nand02 U2946 ( .Y(n8616), .A0(n6461), .A1(n6462) );
  inv02 U2947 ( .Y(n6463), .A(n8584) );
  inv02 U2948 ( .Y(n6464), .A(n8586) );
  inv02 U2949 ( .Y(n6465), .A(n8588) );
  inv02 U2950 ( .Y(n6466), .A(n8351) );
  inv02 U2951 ( .Y(n6467), .A(n8348) );
  nand02 U2952 ( .Y(n6468), .A0(n6465), .A1(n6469) );
  nand02 U2953 ( .Y(n6470), .A0(n5965), .A1(n6471) );
  nand02 U2954 ( .Y(n6472), .A0(n6466), .A1(n6473) );
  nand02 U2955 ( .Y(n6474), .A0(n6466), .A1(n6475) );
  nand02 U2956 ( .Y(n6476), .A0(n6467), .A1(n6477) );
  nand02 U2957 ( .Y(n6478), .A0(n6467), .A1(n6479) );
  nand02 U2958 ( .Y(n6480), .A0(n6467), .A1(n6481) );
  nand02 U2959 ( .Y(n6482), .A0(n6467), .A1(n6483) );
  nand02 U2960 ( .Y(n6484), .A0(n6463), .A1(n6464) );
  inv01 U2961 ( .Y(n6469), .A(n6484) );
  nand02 U2962 ( .Y(n6485), .A0(n6463), .A1(n6464) );
  inv01 U2963 ( .Y(n6471), .A(n6485) );
  nand02 U2964 ( .Y(n6486), .A0(n6463), .A1(n6465) );
  inv01 U2965 ( .Y(n6473), .A(n6486) );
  nand02 U2966 ( .Y(n6487), .A0(n6463), .A1(n5965) );
  inv01 U2967 ( .Y(n6475), .A(n6487) );
  nand02 U2968 ( .Y(n6488), .A0(n6464), .A1(n6465) );
  inv01 U2969 ( .Y(n6477), .A(n6488) );
  nand02 U2970 ( .Y(n6489), .A0(n6464), .A1(n5965) );
  inv01 U2971 ( .Y(n6479), .A(n6489) );
  nand02 U2972 ( .Y(n6490), .A0(n6465), .A1(n6466) );
  inv01 U2973 ( .Y(n6481), .A(n6490) );
  nand02 U2974 ( .Y(n6491), .A0(n5965), .A1(n6466) );
  inv01 U2975 ( .Y(n6483), .A(n6491) );
  nand02 U2976 ( .Y(n6492), .A0(n6468), .A1(n6470) );
  inv01 U2977 ( .Y(n6493), .A(n6492) );
  nand02 U2978 ( .Y(n6494), .A0(n6472), .A1(n6474) );
  inv01 U2979 ( .Y(n6495), .A(n6494) );
  nand02 U2980 ( .Y(n6496), .A0(n6493), .A1(n6495) );
  inv01 U2981 ( .Y(n6461), .A(n6496) );
  nand02 U2982 ( .Y(n6497), .A0(n6476), .A1(n6478) );
  inv01 U2983 ( .Y(n6498), .A(n6497) );
  nand02 U2984 ( .Y(n6499), .A0(n6480), .A1(n6482) );
  inv01 U2985 ( .Y(n6500), .A(n6499) );
  nand02 U2986 ( .Y(n6501), .A0(n6498), .A1(n6500) );
  inv01 U2987 ( .Y(n6462), .A(n6501) );
  nand02 U2988 ( .Y(n8631), .A0(n6502), .A1(n6503) );
  inv02 U2989 ( .Y(n6504), .A(n8609) );
  inv02 U2990 ( .Y(n6505), .A(n8610) );
  inv02 U2991 ( .Y(n6506), .A(n8604) );
  inv02 U2992 ( .Y(n6507), .A(n8347) );
  inv02 U2993 ( .Y(n6508), .A(n8363) );
  nand02 U2994 ( .Y(n6509), .A0(n6506), .A1(n6510) );
  nand02 U2995 ( .Y(n6511), .A0(n5965), .A1(n6512) );
  nand02 U2996 ( .Y(n6513), .A0(n6507), .A1(n6514) );
  nand02 U2997 ( .Y(n6515), .A0(n6507), .A1(n6516) );
  nand02 U2998 ( .Y(n6517), .A0(n6508), .A1(n6518) );
  nand02 U2999 ( .Y(n6519), .A0(n6508), .A1(n6520) );
  nand02 U3000 ( .Y(n6521), .A0(n6508), .A1(n6522) );
  nand02 U3001 ( .Y(n6523), .A0(n6508), .A1(n6524) );
  nand02 U3002 ( .Y(n6525), .A0(n6504), .A1(n6505) );
  inv01 U3003 ( .Y(n6510), .A(n6525) );
  nand02 U3004 ( .Y(n6526), .A0(n6504), .A1(n6505) );
  inv01 U3005 ( .Y(n6512), .A(n6526) );
  nand02 U3006 ( .Y(n6527), .A0(n6504), .A1(n6506) );
  inv01 U3007 ( .Y(n6514), .A(n6527) );
  nand02 U3008 ( .Y(n6528), .A0(n6504), .A1(n5965) );
  inv01 U3009 ( .Y(n6516), .A(n6528) );
  nand02 U3010 ( .Y(n6529), .A0(n6505), .A1(n6506) );
  inv01 U3011 ( .Y(n6518), .A(n6529) );
  nand02 U3012 ( .Y(n6530), .A0(n6505), .A1(n5965) );
  inv01 U3013 ( .Y(n6520), .A(n6530) );
  nand02 U3014 ( .Y(n6531), .A0(n6506), .A1(n6507) );
  inv01 U3015 ( .Y(n6522), .A(n6531) );
  nand02 U3016 ( .Y(n6532), .A0(n5965), .A1(n6507) );
  inv01 U3017 ( .Y(n6524), .A(n6532) );
  nand02 U3018 ( .Y(n6533), .A0(n6509), .A1(n6511) );
  inv01 U3019 ( .Y(n6534), .A(n6533) );
  nand02 U3020 ( .Y(n6535), .A0(n6513), .A1(n6515) );
  inv01 U3021 ( .Y(n6536), .A(n6535) );
  nand02 U3022 ( .Y(n6537), .A0(n6534), .A1(n6536) );
  inv01 U3023 ( .Y(n6502), .A(n6537) );
  nand02 U3024 ( .Y(n6538), .A0(n6517), .A1(n6519) );
  inv01 U3025 ( .Y(n6539), .A(n6538) );
  nand02 U3026 ( .Y(n6540), .A0(n6521), .A1(n6523) );
  inv01 U3027 ( .Y(n6541), .A(n6540) );
  nand02 U3028 ( .Y(n6542), .A0(n6539), .A1(n6541) );
  inv01 U3029 ( .Y(n6503), .A(n6542) );
  nand02 U3030 ( .Y(n8733), .A0(n6543), .A1(n6544) );
  inv02 U3031 ( .Y(n6545), .A(n8601) );
  inv02 U3032 ( .Y(n6546), .A(n8604) );
  inv02 U3033 ( .Y(n6547), .A(n8718) );
  inv02 U3034 ( .Y(n6548), .A(n8351) );
  inv02 U3035 ( .Y(n6549), .A(n8348) );
  nand02 U3036 ( .Y(n6550), .A0(n6547), .A1(n6551) );
  nand02 U3037 ( .Y(n6552), .A0(n5965), .A1(n6553) );
  nand02 U3038 ( .Y(n6554), .A0(n6548), .A1(n6555) );
  nand02 U3039 ( .Y(n6556), .A0(n6548), .A1(n6557) );
  nand02 U3040 ( .Y(n6558), .A0(n6549), .A1(n6559) );
  nand02 U3041 ( .Y(n6560), .A0(n6549), .A1(n6561) );
  nand02 U3042 ( .Y(n6562), .A0(n6549), .A1(n6563) );
  nand02 U3043 ( .Y(n6564), .A0(n6549), .A1(n6565) );
  nand02 U3044 ( .Y(n6566), .A0(n6545), .A1(n6546) );
  inv01 U3045 ( .Y(n6551), .A(n6566) );
  nand02 U3046 ( .Y(n6567), .A0(n6545), .A1(n6546) );
  inv01 U3047 ( .Y(n6553), .A(n6567) );
  nand02 U3048 ( .Y(n6568), .A0(n6545), .A1(n6547) );
  inv01 U3049 ( .Y(n6555), .A(n6568) );
  nand02 U3050 ( .Y(n6569), .A0(n6545), .A1(n5965) );
  inv01 U3051 ( .Y(n6557), .A(n6569) );
  nand02 U3052 ( .Y(n6570), .A0(n6546), .A1(n6547) );
  inv01 U3053 ( .Y(n6559), .A(n6570) );
  nand02 U3054 ( .Y(n6571), .A0(n6546), .A1(n5965) );
  inv01 U3055 ( .Y(n6561), .A(n6571) );
  nand02 U3056 ( .Y(n6572), .A0(n6547), .A1(n6548) );
  inv01 U3057 ( .Y(n6563), .A(n6572) );
  nand02 U3058 ( .Y(n6573), .A0(n5965), .A1(n6548) );
  inv01 U3059 ( .Y(n6565), .A(n6573) );
  nand02 U3060 ( .Y(n6574), .A0(n6550), .A1(n6552) );
  inv01 U3061 ( .Y(n6575), .A(n6574) );
  nand02 U3062 ( .Y(n6576), .A0(n6554), .A1(n6556) );
  inv01 U3063 ( .Y(n6577), .A(n6576) );
  nand02 U3064 ( .Y(n6578), .A0(n6575), .A1(n6577) );
  inv01 U3065 ( .Y(n6543), .A(n6578) );
  nand02 U3066 ( .Y(n6579), .A0(n6558), .A1(n6560) );
  inv01 U3067 ( .Y(n6580), .A(n6579) );
  nand02 U3068 ( .Y(n6581), .A0(n6562), .A1(n6564) );
  inv01 U3069 ( .Y(n6582), .A(n6581) );
  nand02 U3070 ( .Y(n6583), .A0(n6580), .A1(n6582) );
  inv01 U3071 ( .Y(n6544), .A(n6583) );
  inv02 U3072 ( .Y(n8609), .A(n8309) );
  nand02 U3073 ( .Y(n8739), .A0(n6584), .A1(n6585) );
  inv02 U3074 ( .Y(n6586), .A(n8586) );
  inv02 U3075 ( .Y(n6587), .A(n8620) );
  inv02 U3076 ( .Y(n6588), .A(n8584) );
  inv02 U3077 ( .Y(n6589), .A(n8351) );
  inv02 U3078 ( .Y(n6590), .A(n8348) );
  nand02 U3079 ( .Y(n6591), .A0(n6588), .A1(n6592) );
  nand02 U3080 ( .Y(n6593), .A0(n5965), .A1(n6594) );
  nand02 U3081 ( .Y(n6595), .A0(n6589), .A1(n6596) );
  nand02 U3082 ( .Y(n6597), .A0(n6589), .A1(n6598) );
  nand02 U3083 ( .Y(n6599), .A0(n6590), .A1(n6600) );
  nand02 U3084 ( .Y(n6601), .A0(n6590), .A1(n6602) );
  nand02 U3085 ( .Y(n6603), .A0(n6590), .A1(n6604) );
  nand02 U3086 ( .Y(n6605), .A0(n6590), .A1(n6606) );
  nand02 U3087 ( .Y(n6607), .A0(n6586), .A1(n6587) );
  inv01 U3088 ( .Y(n6592), .A(n6607) );
  nand02 U3089 ( .Y(n6608), .A0(n6586), .A1(n6587) );
  inv01 U3090 ( .Y(n6594), .A(n6608) );
  nand02 U3091 ( .Y(n6609), .A0(n6586), .A1(n6588) );
  inv01 U3092 ( .Y(n6596), .A(n6609) );
  nand02 U3093 ( .Y(n6610), .A0(n6586), .A1(n5965) );
  inv01 U3094 ( .Y(n6598), .A(n6610) );
  nand02 U3095 ( .Y(n6611), .A0(n6587), .A1(n6588) );
  inv01 U3096 ( .Y(n6600), .A(n6611) );
  nand02 U3097 ( .Y(n6612), .A0(n6587), .A1(n5965) );
  inv01 U3098 ( .Y(n6602), .A(n6612) );
  nand02 U3099 ( .Y(n6613), .A0(n6588), .A1(n6589) );
  inv01 U3100 ( .Y(n6604), .A(n6613) );
  nand02 U3101 ( .Y(n6614), .A0(n5965), .A1(n6589) );
  inv01 U3102 ( .Y(n6606), .A(n6614) );
  nand02 U3103 ( .Y(n6615), .A0(n6591), .A1(n6593) );
  inv01 U3104 ( .Y(n6616), .A(n6615) );
  nand02 U3105 ( .Y(n6617), .A0(n6595), .A1(n6597) );
  inv01 U3106 ( .Y(n6618), .A(n6617) );
  nand02 U3107 ( .Y(n6619), .A0(n6616), .A1(n6618) );
  inv01 U3108 ( .Y(n6584), .A(n6619) );
  nand02 U3109 ( .Y(n6620), .A0(n6599), .A1(n6601) );
  inv01 U3110 ( .Y(n6621), .A(n6620) );
  nand02 U3111 ( .Y(n6622), .A0(n6603), .A1(n6605) );
  inv01 U3112 ( .Y(n6623), .A(n6622) );
  nand02 U3113 ( .Y(n6624), .A0(n6621), .A1(n6623) );
  inv01 U3114 ( .Y(n6585), .A(n6624) );
  inv02 U3115 ( .Y(n8620), .A(n8032) );
  or04 U3116 ( .Y(n6625), .A0(n8830), .A1(n8831), .A2(n8832), .A3(n8833) );
  inv01 U3117 ( .Y(n6626), .A(n6625) );
  or04 U3118 ( .Y(n6627), .A0(n8838), .A1(n8839), .A2(n8840), .A3(n8841) );
  inv01 U3119 ( .Y(n6628), .A(n6627) );
  nand02 U3120 ( .Y(n8675), .A0(n6629), .A1(n6630) );
  inv01 U3121 ( .Y(n6631), .A(n8678) );
  inv01 U3122 ( .Y(n6632), .A(n8329) );
  inv01 U3123 ( .Y(n6633), .A(n5607) );
  inv02 U3124 ( .Y(n6634), .A(n8606) );
  inv02 U3125 ( .Y(n6635), .A(n8605) );
  nand02 U3126 ( .Y(n6636), .A0(n6631), .A1(n6632) );
  nand02 U3127 ( .Y(n6637), .A0(n6631), .A1(n6504) );
  nand02 U3128 ( .Y(n6638), .A0(n6631), .A1(n6633) );
  nand02 U3129 ( .Y(n6639), .A0(n6632), .A1(n6634) );
  nand02 U3130 ( .Y(n6640), .A0(n6864), .A1(n6634) );
  nand02 U3131 ( .Y(n6641), .A0(n6633), .A1(n6634) );
  nand02 U3132 ( .Y(n6642), .A0(n6632), .A1(n6635) );
  nand02 U3133 ( .Y(n6643), .A0(n5490), .A1(n6635) );
  nand02 U3134 ( .Y(n6644), .A0(n6633), .A1(n6635) );
  nand02 U3135 ( .Y(n6645), .A0(n6636), .A1(n6637) );
  inv01 U3136 ( .Y(n6646), .A(n6645) );
  nand02 U3137 ( .Y(n6647), .A0(n6638), .A1(n6646) );
  inv01 U3138 ( .Y(n6648), .A(n6647) );
  nand02 U3139 ( .Y(n6649), .A0(n6639), .A1(n6640) );
  inv01 U3140 ( .Y(n6650), .A(n6649) );
  nand02 U3141 ( .Y(n6651), .A0(n6648), .A1(n6650) );
  inv01 U3142 ( .Y(n6629), .A(n6651) );
  nand02 U3143 ( .Y(n6652), .A0(n6641), .A1(n6642) );
  inv01 U3144 ( .Y(n6653), .A(n6652) );
  nand02 U3145 ( .Y(n6654), .A0(n6643), .A1(n6644) );
  inv01 U3146 ( .Y(n6655), .A(n6654) );
  nand02 U3147 ( .Y(n6656), .A0(n6653), .A1(n6655) );
  inv01 U3148 ( .Y(n6630), .A(n6656) );
  nand02 U3149 ( .Y(n8736), .A0(n6657), .A1(n6658) );
  inv02 U3150 ( .Y(n6659), .A(n5607) );
  inv02 U3151 ( .Y(n6660), .A(n8163) );
  inv02 U3152 ( .Y(n6661), .A(n8320) );
  inv02 U3153 ( .Y(n6662), .A(n8677) );
  inv02 U3154 ( .Y(n6663), .A(n8609) );
  inv02 U3155 ( .Y(n6664), .A(n8603) );
  nand02 U3156 ( .Y(n6665), .A0(n6661), .A1(n6666) );
  nand02 U3157 ( .Y(n6667), .A0(n6662), .A1(n6668) );
  nand02 U3158 ( .Y(n6669), .A0(n6663), .A1(n6670) );
  nand02 U3159 ( .Y(n6671), .A0(n6663), .A1(n6672) );
  nand02 U3160 ( .Y(n6673), .A0(n6664), .A1(n6674) );
  nand02 U3161 ( .Y(n6675), .A0(n6664), .A1(n6676) );
  nand02 U3162 ( .Y(n6677), .A0(n6664), .A1(n6678) );
  nand02 U3163 ( .Y(n6679), .A0(n6664), .A1(n6680) );
  nand02 U3164 ( .Y(n6681), .A0(n6659), .A1(n6660) );
  inv01 U3165 ( .Y(n6666), .A(n6681) );
  nand02 U3166 ( .Y(n6682), .A0(n6659), .A1(n6660) );
  inv01 U3167 ( .Y(n6668), .A(n6682) );
  nand02 U3168 ( .Y(n6683), .A0(n6659), .A1(n6661) );
  inv01 U3169 ( .Y(n6670), .A(n6683) );
  nand02 U3170 ( .Y(n6684), .A0(n6659), .A1(n6662) );
  inv01 U3171 ( .Y(n6672), .A(n6684) );
  nand02 U3172 ( .Y(n6685), .A0(n6660), .A1(n6661) );
  inv01 U3173 ( .Y(n6674), .A(n6685) );
  nand02 U3174 ( .Y(n6686), .A0(n6660), .A1(n6662) );
  inv01 U3175 ( .Y(n6676), .A(n6686) );
  nand02 U3176 ( .Y(n6687), .A0(n6661), .A1(n6663) );
  inv01 U3177 ( .Y(n6678), .A(n6687) );
  nand02 U3178 ( .Y(n6688), .A0(n6662), .A1(n6663) );
  inv01 U3179 ( .Y(n6680), .A(n6688) );
  nand02 U3180 ( .Y(n6689), .A0(n6665), .A1(n6667) );
  inv01 U3181 ( .Y(n6690), .A(n6689) );
  nand02 U3182 ( .Y(n6691), .A0(n6669), .A1(n6671) );
  inv01 U3183 ( .Y(n6692), .A(n6691) );
  nand02 U3184 ( .Y(n6693), .A0(n6690), .A1(n6692) );
  inv01 U3185 ( .Y(n6657), .A(n6693) );
  nand02 U3186 ( .Y(n6694), .A0(n6673), .A1(n6675) );
  inv01 U3187 ( .Y(n6695), .A(n6694) );
  nand02 U3188 ( .Y(n6696), .A0(n6677), .A1(n6679) );
  inv01 U3189 ( .Y(n6697), .A(n6696) );
  nand02 U3190 ( .Y(n6698), .A0(n6695), .A1(n6697) );
  inv01 U3191 ( .Y(n6658), .A(n6698) );
  nand02 U3192 ( .Y(n8711), .A0(n6699), .A1(n6700) );
  inv02 U3193 ( .Y(n6701), .A(n8665) );
  inv02 U3194 ( .Y(n6702), .A(n8171) );
  inv02 U3195 ( .Y(n6703), .A(n8664) );
  inv02 U3196 ( .Y(n6704), .A(n8337) );
  inv02 U3197 ( .Y(n6705), .A(n8281) );
  inv02 U3198 ( .Y(n6706), .A(n8363) );
  nand02 U3199 ( .Y(n6707), .A0(n6703), .A1(n6708) );
  nand02 U3200 ( .Y(n6709), .A0(n6704), .A1(n6710) );
  nand02 U3201 ( .Y(n6711), .A0(n6705), .A1(n6712) );
  nand02 U3202 ( .Y(n6713), .A0(n6705), .A1(n6714) );
  nand02 U3203 ( .Y(n6715), .A0(n6706), .A1(n6716) );
  nand02 U3204 ( .Y(n6717), .A0(n6706), .A1(n6718) );
  nand02 U3205 ( .Y(n6719), .A0(n6706), .A1(n6720) );
  nand02 U3206 ( .Y(n6721), .A0(n6706), .A1(n6722) );
  nand02 U3207 ( .Y(n6723), .A0(n6701), .A1(n6702) );
  inv01 U3208 ( .Y(n6708), .A(n6723) );
  nand02 U3209 ( .Y(n6724), .A0(n6701), .A1(n6702) );
  inv01 U3210 ( .Y(n6710), .A(n6724) );
  nand02 U3211 ( .Y(n6725), .A0(n6701), .A1(n6703) );
  inv01 U3212 ( .Y(n6712), .A(n6725) );
  nand02 U3213 ( .Y(n6726), .A0(n6701), .A1(n6704) );
  inv01 U3214 ( .Y(n6714), .A(n6726) );
  nand02 U3215 ( .Y(n6727), .A0(n6702), .A1(n6703) );
  inv01 U3216 ( .Y(n6716), .A(n6727) );
  nand02 U3217 ( .Y(n6728), .A0(n6702), .A1(n6704) );
  inv01 U3218 ( .Y(n6718), .A(n6728) );
  nand02 U3219 ( .Y(n6729), .A0(n6703), .A1(n6705) );
  inv01 U3220 ( .Y(n6720), .A(n6729) );
  nand02 U3221 ( .Y(n6730), .A0(n6704), .A1(n6705) );
  inv01 U3222 ( .Y(n6722), .A(n6730) );
  nand02 U3223 ( .Y(n6731), .A0(n6707), .A1(n6709) );
  inv01 U3224 ( .Y(n6732), .A(n6731) );
  nand02 U3225 ( .Y(n6733), .A0(n6711), .A1(n6713) );
  inv01 U3226 ( .Y(n6734), .A(n6733) );
  nand02 U3227 ( .Y(n6735), .A0(n6732), .A1(n6734) );
  inv01 U3228 ( .Y(n6699), .A(n6735) );
  nand02 U3229 ( .Y(n6736), .A0(n6715), .A1(n6717) );
  inv01 U3230 ( .Y(n6737), .A(n6736) );
  nand02 U3231 ( .Y(n6738), .A0(n6719), .A1(n6721) );
  inv01 U3232 ( .Y(n6739), .A(n6738) );
  nand02 U3233 ( .Y(n6740), .A0(n6737), .A1(n6739) );
  inv01 U3234 ( .Y(n6700), .A(n6740) );
  nand02 U3235 ( .Y(n8667), .A0(n6741), .A1(n6742) );
  inv02 U3236 ( .Y(n6743), .A(n8674) );
  inv02 U3237 ( .Y(n6744), .A(n8673) );
  inv02 U3238 ( .Y(n6745), .A(n8595) );
  inv02 U3239 ( .Y(n6746), .A(n8345) );
  inv02 U3240 ( .Y(n6747), .A(n8338) );
  inv02 U3241 ( .Y(n6748), .A(n8337) );
  nand02 U3242 ( .Y(n6749), .A0(n6745), .A1(n6750) );
  nand02 U3243 ( .Y(n6751), .A0(n6746), .A1(n6752) );
  nand02 U3244 ( .Y(n6753), .A0(n6747), .A1(n6754) );
  nand02 U3245 ( .Y(n6755), .A0(n6747), .A1(n6756) );
  nand02 U3246 ( .Y(n6757), .A0(n6748), .A1(n6758) );
  nand02 U3247 ( .Y(n6759), .A0(n6748), .A1(n6760) );
  nand02 U3248 ( .Y(n6761), .A0(n6748), .A1(n6762) );
  nand02 U3249 ( .Y(n6763), .A0(n6748), .A1(n6764) );
  nand02 U3250 ( .Y(n6765), .A0(n6743), .A1(n6744) );
  inv01 U3251 ( .Y(n6750), .A(n6765) );
  nand02 U3252 ( .Y(n6766), .A0(n6743), .A1(n6744) );
  inv01 U3253 ( .Y(n6752), .A(n6766) );
  nand02 U3254 ( .Y(n6767), .A0(n6743), .A1(n6745) );
  inv01 U3255 ( .Y(n6754), .A(n6767) );
  nand02 U3256 ( .Y(n6768), .A0(n6743), .A1(n6746) );
  inv01 U3257 ( .Y(n6756), .A(n6768) );
  nand02 U3258 ( .Y(n6769), .A0(n6744), .A1(n6745) );
  inv01 U3259 ( .Y(n6758), .A(n6769) );
  nand02 U3260 ( .Y(n6770), .A0(n6744), .A1(n6746) );
  inv01 U3261 ( .Y(n6760), .A(n6770) );
  nand02 U3262 ( .Y(n6771), .A0(n6745), .A1(n6747) );
  inv01 U3263 ( .Y(n6762), .A(n6771) );
  nand02 U3264 ( .Y(n6772), .A0(n6746), .A1(n6747) );
  inv01 U3265 ( .Y(n6764), .A(n6772) );
  nand02 U3266 ( .Y(n6773), .A0(n6749), .A1(n6751) );
  inv01 U3267 ( .Y(n6774), .A(n6773) );
  nand02 U3268 ( .Y(n6775), .A0(n6753), .A1(n6755) );
  inv01 U3269 ( .Y(n6776), .A(n6775) );
  nand02 U3270 ( .Y(n6777), .A0(n6774), .A1(n6776) );
  inv01 U3271 ( .Y(n6741), .A(n6777) );
  nand02 U3272 ( .Y(n6778), .A0(n6757), .A1(n6759) );
  inv01 U3273 ( .Y(n6779), .A(n6778) );
  nand02 U3274 ( .Y(n6780), .A0(n6761), .A1(n6763) );
  inv01 U3275 ( .Y(n6781), .A(n6780) );
  nand02 U3276 ( .Y(n6782), .A0(n6779), .A1(n6781) );
  inv01 U3277 ( .Y(n6742), .A(n6782) );
  inv04 U3278 ( .Y(n8345), .A(n8342) );
  inv01 U3279 ( .Y(n8583), .A(n6783) );
  nor02 U3280 ( .Y(n6784), .A0(n8586), .A1(n6785) );
  nor02 U3281 ( .Y(n6786), .A0(n8586), .A1(n6787) );
  nor02 U3282 ( .Y(n6788), .A0(n8586), .A1(n6789) );
  nor02 U3283 ( .Y(n6790), .A0(n8586), .A1(n6791) );
  nor02 U3284 ( .Y(n6792), .A0(n8345), .A1(n6793) );
  nor02 U3285 ( .Y(n6794), .A0(n8345), .A1(n6795) );
  nor02 U3286 ( .Y(n6796), .A0(n8345), .A1(n6797) );
  nor02 U3287 ( .Y(n6798), .A0(n8345), .A1(n6799) );
  nor02 U3288 ( .Y(n6783), .A0(n6800), .A1(n6801) );
  nor02 U3289 ( .Y(n6802), .A0(n8584), .A1(n8585) );
  inv01 U3290 ( .Y(n6785), .A(n6802) );
  nor02 U3291 ( .Y(n6803), .A0(n8350), .A1(n8585) );
  inv01 U3292 ( .Y(n6787), .A(n6803) );
  nor02 U3293 ( .Y(n6804), .A0(n8584), .A1(n8335) );
  inv01 U3294 ( .Y(n6789), .A(n6804) );
  nor02 U3295 ( .Y(n6805), .A0(n8350), .A1(n8335) );
  inv01 U3296 ( .Y(n6791), .A(n6805) );
  nor02 U3297 ( .Y(n6806), .A0(n8584), .A1(n8585) );
  inv01 U3298 ( .Y(n6793), .A(n6806) );
  nor02 U3299 ( .Y(n6807), .A0(n8350), .A1(n8585) );
  inv01 U3300 ( .Y(n6795), .A(n6807) );
  inv01 U3301 ( .Y(n6797), .A(n6804) );
  nor02 U3302 ( .Y(n6808), .A0(n8350), .A1(n8335) );
  inv01 U3303 ( .Y(n6799), .A(n6808) );
  nor02 U3304 ( .Y(n6809), .A0(n6784), .A1(n6786) );
  inv01 U3305 ( .Y(n6810), .A(n6809) );
  nor02 U3306 ( .Y(n6811), .A0(n6788), .A1(n6790) );
  inv01 U3307 ( .Y(n6812), .A(n6811) );
  nor02 U3308 ( .Y(n6813), .A0(n6810), .A1(n6812) );
  inv01 U3309 ( .Y(n6800), .A(n6813) );
  nor02 U3310 ( .Y(n6814), .A0(n6792), .A1(n6794) );
  inv01 U3311 ( .Y(n6815), .A(n6814) );
  nor02 U3312 ( .Y(n6816), .A0(n6796), .A1(n6798) );
  inv01 U3313 ( .Y(n6817), .A(n6816) );
  nor02 U3314 ( .Y(n6818), .A0(n6815), .A1(n6817) );
  inv01 U3315 ( .Y(n6801), .A(n6818) );
  nand02 U3316 ( .Y(n8591), .A0(n6819), .A1(n6820) );
  inv02 U3317 ( .Y(n6821), .A(n8594) );
  inv02 U3318 ( .Y(n6822), .A(n8593) );
  inv02 U3319 ( .Y(n6823), .A(n8592) );
  inv02 U3320 ( .Y(n6824), .A(n8348) );
  inv02 U3321 ( .Y(n6825), .A(n8344) );
  inv02 U3322 ( .Y(n6826), .A(n8336) );
  nand02 U3323 ( .Y(n6827), .A0(n6823), .A1(n6828) );
  nand02 U3324 ( .Y(n6829), .A0(n6824), .A1(n6830) );
  nand02 U3325 ( .Y(n6831), .A0(n6825), .A1(n6832) );
  nand02 U3326 ( .Y(n6833), .A0(n6825), .A1(n6834) );
  nand02 U3327 ( .Y(n6835), .A0(n6826), .A1(n6836) );
  nand02 U3328 ( .Y(n6837), .A0(n6826), .A1(n6838) );
  nand02 U3329 ( .Y(n6839), .A0(n6826), .A1(n6840) );
  nand02 U3330 ( .Y(n6841), .A0(n6826), .A1(n6842) );
  nand02 U3331 ( .Y(n6843), .A0(n6821), .A1(n6822) );
  inv01 U3332 ( .Y(n6828), .A(n6843) );
  nand02 U3333 ( .Y(n6844), .A0(n6821), .A1(n6822) );
  inv01 U3334 ( .Y(n6830), .A(n6844) );
  nand02 U3335 ( .Y(n6845), .A0(n6821), .A1(n6823) );
  inv01 U3336 ( .Y(n6832), .A(n6845) );
  nand02 U3337 ( .Y(n6846), .A0(n6821), .A1(n6824) );
  inv01 U3338 ( .Y(n6834), .A(n6846) );
  nand02 U3339 ( .Y(n6847), .A0(n6822), .A1(n6823) );
  inv01 U3340 ( .Y(n6836), .A(n6847) );
  nand02 U3341 ( .Y(n6848), .A0(n6822), .A1(n6824) );
  inv01 U3342 ( .Y(n6838), .A(n6848) );
  nand02 U3343 ( .Y(n6849), .A0(n6823), .A1(n6825) );
  inv01 U3344 ( .Y(n6840), .A(n6849) );
  nand02 U3345 ( .Y(n6850), .A0(n6824), .A1(n6825) );
  inv01 U3346 ( .Y(n6842), .A(n6850) );
  nand02 U3347 ( .Y(n6851), .A0(n6827), .A1(n6829) );
  inv01 U3348 ( .Y(n6852), .A(n6851) );
  nand02 U3349 ( .Y(n6853), .A0(n6831), .A1(n6833) );
  inv01 U3350 ( .Y(n6854), .A(n6853) );
  nand02 U3351 ( .Y(n6855), .A0(n6852), .A1(n6854) );
  inv01 U3352 ( .Y(n6819), .A(n6855) );
  nand02 U3353 ( .Y(n6856), .A0(n6835), .A1(n6837) );
  inv01 U3354 ( .Y(n6857), .A(n6856) );
  nand02 U3355 ( .Y(n6858), .A0(n6839), .A1(n6841) );
  inv01 U3356 ( .Y(n6859), .A(n6858) );
  nand02 U3357 ( .Y(n6860), .A0(n6857), .A1(n6859) );
  inv01 U3358 ( .Y(n6820), .A(n6860) );
  inv04 U3359 ( .Y(n8350), .A(n8349) );
  inv02 U3360 ( .Y(n8593), .A(n8038) );
  nand02 U3361 ( .Y(n8700), .A0(n6861), .A1(n6862) );
  inv02 U3362 ( .Y(n6863), .A(n8642) );
  inv02 U3363 ( .Y(n6864), .A(n8609) );
  inv02 U3364 ( .Y(n6865), .A(n8633) );
  inv02 U3365 ( .Y(n6866), .A(n8678) );
  inv02 U3366 ( .Y(n6867), .A(n8281) );
  inv02 U3367 ( .Y(n6868), .A(n8363) );
  nand02 U3368 ( .Y(n6869), .A0(n6865), .A1(n6870) );
  nand02 U3369 ( .Y(n6871), .A0(n6866), .A1(n6872) );
  nand02 U3370 ( .Y(n6873), .A0(n6867), .A1(n6874) );
  nand02 U3371 ( .Y(n6875), .A0(n6867), .A1(n6876) );
  nand02 U3372 ( .Y(n6877), .A0(n6868), .A1(n6878) );
  nand02 U3373 ( .Y(n6879), .A0(n6868), .A1(n6880) );
  nand02 U3374 ( .Y(n6881), .A0(n6868), .A1(n6882) );
  nand02 U3375 ( .Y(n6883), .A0(n6868), .A1(n6884) );
  nand02 U3376 ( .Y(n6885), .A0(n6863), .A1(n6864) );
  inv01 U3377 ( .Y(n6870), .A(n6885) );
  nand02 U3378 ( .Y(n6886), .A0(n6863), .A1(n6864) );
  inv01 U3379 ( .Y(n6872), .A(n6886) );
  nand02 U3380 ( .Y(n6887), .A0(n6863), .A1(n6865) );
  inv01 U3381 ( .Y(n6874), .A(n6887) );
  nand02 U3382 ( .Y(n6888), .A0(n6863), .A1(n6866) );
  inv01 U3383 ( .Y(n6876), .A(n6888) );
  nand02 U3384 ( .Y(n6889), .A0(n6864), .A1(n6865) );
  inv01 U3385 ( .Y(n6878), .A(n6889) );
  nand02 U3386 ( .Y(n6890), .A0(n6864), .A1(n6866) );
  inv01 U3387 ( .Y(n6880), .A(n6890) );
  nand02 U3388 ( .Y(n6891), .A0(n6865), .A1(n6867) );
  inv01 U3389 ( .Y(n6882), .A(n6891) );
  nand02 U3390 ( .Y(n6892), .A0(n6866), .A1(n6867) );
  inv01 U3391 ( .Y(n6884), .A(n6892) );
  nand02 U3392 ( .Y(n6893), .A0(n6869), .A1(n6871) );
  inv01 U3393 ( .Y(n6894), .A(n6893) );
  nand02 U3394 ( .Y(n6895), .A0(n6873), .A1(n6875) );
  inv01 U3395 ( .Y(n6896), .A(n6895) );
  nand02 U3396 ( .Y(n6897), .A0(n6894), .A1(n6896) );
  inv01 U3397 ( .Y(n6861), .A(n6897) );
  nand02 U3398 ( .Y(n6898), .A0(n6877), .A1(n6879) );
  inv01 U3399 ( .Y(n6899), .A(n6898) );
  nand02 U3400 ( .Y(n6900), .A0(n6881), .A1(n6883) );
  inv01 U3401 ( .Y(n6901), .A(n6900) );
  nand02 U3402 ( .Y(n6902), .A0(n6899), .A1(n6901) );
  inv01 U3403 ( .Y(n6862), .A(n6902) );
  nand02 U3404 ( .Y(n8623), .A0(n6903), .A1(n6904) );
  inv02 U3405 ( .Y(n6905), .A(n8625) );
  inv02 U3406 ( .Y(n6906), .A(n8624) );
  inv02 U3407 ( .Y(n6907), .A(n8593) );
  inv02 U3408 ( .Y(n6908), .A(n8350) );
  inv02 U3409 ( .Y(n6909), .A(n8327) );
  inv02 U3410 ( .Y(n6910), .A(n8005) );
  nand02 U3411 ( .Y(n6911), .A0(n6907), .A1(n6912) );
  nand02 U3412 ( .Y(n6913), .A0(n6908), .A1(n6914) );
  nand02 U3413 ( .Y(n6915), .A0(n6909), .A1(n6916) );
  nand02 U3414 ( .Y(n6917), .A0(n6909), .A1(n6918) );
  nand02 U3415 ( .Y(n6919), .A0(n6910), .A1(n6920) );
  nand02 U3416 ( .Y(n6921), .A0(n6910), .A1(n6922) );
  nand02 U3417 ( .Y(n6923), .A0(n6910), .A1(n6924) );
  nand02 U3418 ( .Y(n6925), .A0(n6910), .A1(n6926) );
  nand02 U3419 ( .Y(n6927), .A0(n6905), .A1(n6906) );
  inv01 U3420 ( .Y(n6912), .A(n6927) );
  nand02 U3421 ( .Y(n6928), .A0(n6905), .A1(n6906) );
  inv01 U3422 ( .Y(n6914), .A(n6928) );
  nand02 U3423 ( .Y(n6929), .A0(n6905), .A1(n6907) );
  inv01 U3424 ( .Y(n6916), .A(n6929) );
  nand02 U3425 ( .Y(n6930), .A0(n6905), .A1(n6908) );
  inv01 U3426 ( .Y(n6918), .A(n6930) );
  nand02 U3427 ( .Y(n6931), .A0(n6906), .A1(n6907) );
  inv01 U3428 ( .Y(n6920), .A(n6931) );
  nand02 U3429 ( .Y(n6932), .A0(n6906), .A1(n6908) );
  inv01 U3430 ( .Y(n6922), .A(n6932) );
  nand02 U3431 ( .Y(n6933), .A0(n6907), .A1(n6909) );
  inv01 U3432 ( .Y(n6924), .A(n6933) );
  nand02 U3433 ( .Y(n6934), .A0(n6908), .A1(n6909) );
  inv01 U3434 ( .Y(n6926), .A(n6934) );
  nand02 U3435 ( .Y(n6935), .A0(n6911), .A1(n6913) );
  inv01 U3436 ( .Y(n6936), .A(n6935) );
  nand02 U3437 ( .Y(n6937), .A0(n6915), .A1(n6917) );
  inv01 U3438 ( .Y(n6938), .A(n6937) );
  nand02 U3439 ( .Y(n6939), .A0(n6936), .A1(n6938) );
  inv01 U3440 ( .Y(n6903), .A(n6939) );
  nand02 U3441 ( .Y(n6940), .A0(n6919), .A1(n6921) );
  inv01 U3442 ( .Y(n6941), .A(n6940) );
  nand02 U3443 ( .Y(n6942), .A0(n6923), .A1(n6925) );
  inv01 U3444 ( .Y(n6943), .A(n6942) );
  nand02 U3445 ( .Y(n6944), .A0(n6941), .A1(n6943) );
  inv01 U3446 ( .Y(n6904), .A(n6944) );
  nand02 U3447 ( .Y(n8632), .A0(n6945), .A1(n6946) );
  inv02 U3448 ( .Y(n6947), .A(n8634) );
  inv02 U3449 ( .Y(n6948), .A(n8633) );
  inv02 U3450 ( .Y(n6949), .A(n8607) );
  inv02 U3451 ( .Y(n6950), .A(n8350) );
  inv02 U3452 ( .Y(n6951), .A(n8327) );
  inv02 U3453 ( .Y(n6952), .A(n8005) );
  nand02 U3454 ( .Y(n6953), .A0(n6949), .A1(n6954) );
  nand02 U3455 ( .Y(n6955), .A0(n6950), .A1(n6956) );
  nand02 U3456 ( .Y(n6957), .A0(n6951), .A1(n6958) );
  nand02 U3457 ( .Y(n6959), .A0(n6951), .A1(n6960) );
  nand02 U3458 ( .Y(n6961), .A0(n6952), .A1(n6962) );
  nand02 U3459 ( .Y(n6963), .A0(n6952), .A1(n6964) );
  nand02 U3460 ( .Y(n6965), .A0(n6952), .A1(n6966) );
  nand02 U3461 ( .Y(n6967), .A0(n6952), .A1(n6968) );
  nand02 U3462 ( .Y(n6969), .A0(n6947), .A1(n6948) );
  inv01 U3463 ( .Y(n6954), .A(n6969) );
  nand02 U3464 ( .Y(n6970), .A0(n6947), .A1(n6948) );
  inv01 U3465 ( .Y(n6956), .A(n6970) );
  nand02 U3466 ( .Y(n6971), .A0(n6947), .A1(n6949) );
  inv01 U3467 ( .Y(n6958), .A(n6971) );
  nand02 U3468 ( .Y(n6972), .A0(n6947), .A1(n6950) );
  inv01 U3469 ( .Y(n6960), .A(n6972) );
  nand02 U3470 ( .Y(n6973), .A0(n6948), .A1(n6949) );
  inv01 U3471 ( .Y(n6962), .A(n6973) );
  nand02 U3472 ( .Y(n6974), .A0(n6948), .A1(n6950) );
  inv01 U3473 ( .Y(n6964), .A(n6974) );
  nand02 U3474 ( .Y(n6975), .A0(n6949), .A1(n6951) );
  inv01 U3475 ( .Y(n6966), .A(n6975) );
  nand02 U3476 ( .Y(n6976), .A0(n6950), .A1(n6951) );
  inv01 U3477 ( .Y(n6968), .A(n6976) );
  nand02 U3478 ( .Y(n6977), .A0(n6953), .A1(n6955) );
  inv01 U3479 ( .Y(n6978), .A(n6977) );
  nand02 U3480 ( .Y(n6979), .A0(n6957), .A1(n6959) );
  inv01 U3481 ( .Y(n6980), .A(n6979) );
  nand02 U3482 ( .Y(n6981), .A0(n6978), .A1(n6980) );
  inv01 U3483 ( .Y(n6945), .A(n6981) );
  nand02 U3484 ( .Y(n6982), .A0(n6961), .A1(n6963) );
  inv01 U3485 ( .Y(n6983), .A(n6982) );
  nand02 U3486 ( .Y(n6984), .A0(n6965), .A1(n6967) );
  inv01 U3487 ( .Y(n6985), .A(n6984) );
  nand02 U3488 ( .Y(n6986), .A0(n6983), .A1(n6985) );
  inv01 U3489 ( .Y(n6946), .A(n6986) );
  nand02 U3490 ( .Y(n8696), .A0(n6987), .A1(n6988) );
  inv02 U3491 ( .Y(n6989), .A(n8669) );
  inv02 U3492 ( .Y(n6990), .A(n8630) );
  inv02 U3493 ( .Y(n6991), .A(n8678) );
  inv02 U3494 ( .Y(n6992), .A(n8281) );
  inv02 U3495 ( .Y(n6993), .A(n8363) );
  nand02 U3496 ( .Y(n6994), .A0(n6906), .A1(n6995) );
  nand02 U3497 ( .Y(n6996), .A0(n6991), .A1(n6997) );
  nand02 U3498 ( .Y(n6998), .A0(n6992), .A1(n6999) );
  nand02 U3499 ( .Y(n7000), .A0(n6992), .A1(n7001) );
  nand02 U3500 ( .Y(n7002), .A0(n6993), .A1(n7003) );
  nand02 U3501 ( .Y(n7004), .A0(n6993), .A1(n7005) );
  nand02 U3502 ( .Y(n7006), .A0(n6993), .A1(n7007) );
  nand02 U3503 ( .Y(n7008), .A0(n6993), .A1(n7009) );
  nand02 U3504 ( .Y(n7010), .A0(n6989), .A1(n6990) );
  inv01 U3505 ( .Y(n6995), .A(n7010) );
  nand02 U3506 ( .Y(n7011), .A0(n6989), .A1(n6990) );
  inv01 U3507 ( .Y(n6997), .A(n7011) );
  nand02 U3508 ( .Y(n7012), .A0(n6989), .A1(n6906) );
  inv01 U3509 ( .Y(n6999), .A(n7012) );
  nand02 U3510 ( .Y(n7013), .A0(n6989), .A1(n6991) );
  inv01 U3511 ( .Y(n7001), .A(n7013) );
  nand02 U3512 ( .Y(n7014), .A0(n6990), .A1(n6906) );
  inv01 U3513 ( .Y(n7003), .A(n7014) );
  nand02 U3514 ( .Y(n7015), .A0(n6990), .A1(n6991) );
  inv01 U3515 ( .Y(n7005), .A(n7015) );
  nand02 U3516 ( .Y(n7016), .A0(n6906), .A1(n6992) );
  inv01 U3517 ( .Y(n7007), .A(n7016) );
  nand02 U3518 ( .Y(n7017), .A0(n6991), .A1(n6992) );
  inv01 U3519 ( .Y(n7009), .A(n7017) );
  nand02 U3520 ( .Y(n7018), .A0(n6994), .A1(n6996) );
  inv01 U3521 ( .Y(n7019), .A(n7018) );
  nand02 U3522 ( .Y(n7020), .A0(n6998), .A1(n7000) );
  inv01 U3523 ( .Y(n7021), .A(n7020) );
  nand02 U3524 ( .Y(n7022), .A0(n7019), .A1(n7021) );
  inv01 U3525 ( .Y(n6987), .A(n7022) );
  nand02 U3526 ( .Y(n7023), .A0(n7002), .A1(n7004) );
  inv01 U3527 ( .Y(n7024), .A(n7023) );
  nand02 U3528 ( .Y(n7025), .A0(n7006), .A1(n7008) );
  inv01 U3529 ( .Y(n7026), .A(n7025) );
  nand02 U3530 ( .Y(n7027), .A0(n7024), .A1(n7026) );
  inv01 U3531 ( .Y(n6988), .A(n7027) );
  nand02 U3532 ( .Y(n8707), .A0(n7028), .A1(n7029) );
  inv02 U3533 ( .Y(n7030), .A(n8657) );
  inv02 U3534 ( .Y(n7031), .A(n8307) );
  inv02 U3535 ( .Y(n7032), .A(n8692) );
  inv02 U3536 ( .Y(n7033), .A(n8678) );
  inv02 U3537 ( .Y(n7034), .A(n8281) );
  inv02 U3538 ( .Y(n7035), .A(n8363) );
  nand02 U3539 ( .Y(n7036), .A0(n7032), .A1(n7037) );
  nand02 U3540 ( .Y(n7038), .A0(n7033), .A1(n7039) );
  nand02 U3541 ( .Y(n7040), .A0(n7034), .A1(n7041) );
  nand02 U3542 ( .Y(n7042), .A0(n7034), .A1(n7043) );
  nand02 U3543 ( .Y(n7044), .A0(n7035), .A1(n7045) );
  nand02 U3544 ( .Y(n7046), .A0(n7035), .A1(n7047) );
  nand02 U3545 ( .Y(n7048), .A0(n7035), .A1(n7049) );
  nand02 U3546 ( .Y(n7050), .A0(n7035), .A1(n7051) );
  nand02 U3547 ( .Y(n7052), .A0(n7030), .A1(n7031) );
  inv01 U3548 ( .Y(n7037), .A(n7052) );
  nand02 U3549 ( .Y(n7053), .A0(n7030), .A1(n7031) );
  inv01 U3550 ( .Y(n7039), .A(n7053) );
  nand02 U3551 ( .Y(n7054), .A0(n7030), .A1(n7032) );
  inv01 U3552 ( .Y(n7041), .A(n7054) );
  nand02 U3553 ( .Y(n7055), .A0(n7030), .A1(n7033) );
  inv01 U3554 ( .Y(n7043), .A(n7055) );
  nand02 U3555 ( .Y(n7056), .A0(n7031), .A1(n7032) );
  inv01 U3556 ( .Y(n7045), .A(n7056) );
  nand02 U3557 ( .Y(n7057), .A0(n7031), .A1(n7033) );
  inv01 U3558 ( .Y(n7047), .A(n7057) );
  nand02 U3559 ( .Y(n7058), .A0(n7032), .A1(n7034) );
  inv01 U3560 ( .Y(n7049), .A(n7058) );
  nand02 U3561 ( .Y(n7059), .A0(n7033), .A1(n7034) );
  inv01 U3562 ( .Y(n7051), .A(n7059) );
  nand02 U3563 ( .Y(n7060), .A0(n7036), .A1(n7038) );
  inv01 U3564 ( .Y(n7061), .A(n7060) );
  nand02 U3565 ( .Y(n7062), .A0(n7040), .A1(n7042) );
  inv01 U3566 ( .Y(n7063), .A(n7062) );
  nand02 U3567 ( .Y(n7064), .A0(n7061), .A1(n7063) );
  inv01 U3568 ( .Y(n7028), .A(n7064) );
  nand02 U3569 ( .Y(n7065), .A0(n7044), .A1(n7046) );
  inv01 U3570 ( .Y(n7066), .A(n7065) );
  nand02 U3571 ( .Y(n7067), .A0(n7048), .A1(n7050) );
  inv01 U3572 ( .Y(n7068), .A(n7067) );
  nand02 U3573 ( .Y(n7069), .A0(n7066), .A1(n7068) );
  inv01 U3574 ( .Y(n7029), .A(n7069) );
  inv02 U3575 ( .Y(n8669), .A(n8044) );
  nand02 U3576 ( .Y(n8734), .A0(n7070), .A1(n7071) );
  inv02 U3577 ( .Y(n7072), .A(n8610) );
  inv02 U3578 ( .Y(n7073), .A(n8069) );
  inv02 U3579 ( .Y(n7074), .A(n8635) );
  inv02 U3580 ( .Y(n7075), .A(n8335) );
  inv02 U3581 ( .Y(n7076), .A(n8735) );
  inv02 U3582 ( .Y(n7077), .A(n8344) );
  nand02 U3583 ( .Y(n7078), .A0(n7074), .A1(n7079) );
  nand02 U3584 ( .Y(n7080), .A0(n7075), .A1(n7081) );
  nand02 U3585 ( .Y(n7082), .A0(n7076), .A1(n7083) );
  nand02 U3586 ( .Y(n7084), .A0(n7076), .A1(n7085) );
  nand02 U3587 ( .Y(n7086), .A0(n7077), .A1(n7087) );
  nand02 U3588 ( .Y(n7088), .A0(n7077), .A1(n7089) );
  nand02 U3589 ( .Y(n7090), .A0(n7077), .A1(n7091) );
  nand02 U3590 ( .Y(n7092), .A0(n7077), .A1(n7093) );
  nand02 U3591 ( .Y(n7094), .A0(n7072), .A1(n7073) );
  inv01 U3592 ( .Y(n7079), .A(n7094) );
  nand02 U3593 ( .Y(n7095), .A0(n7072), .A1(n7073) );
  inv01 U3594 ( .Y(n7081), .A(n7095) );
  nand02 U3595 ( .Y(n7096), .A0(n7072), .A1(n7074) );
  inv01 U3596 ( .Y(n7083), .A(n7096) );
  nand02 U3597 ( .Y(n7097), .A0(n7072), .A1(n7075) );
  inv01 U3598 ( .Y(n7085), .A(n7097) );
  nand02 U3599 ( .Y(n7098), .A0(n7073), .A1(n7074) );
  inv01 U3600 ( .Y(n7087), .A(n7098) );
  nand02 U3601 ( .Y(n7099), .A0(n7073), .A1(n7075) );
  inv01 U3602 ( .Y(n7089), .A(n7099) );
  nand02 U3603 ( .Y(n7100), .A0(n7074), .A1(n7076) );
  inv01 U3604 ( .Y(n7091), .A(n7100) );
  nand02 U3605 ( .Y(n7101), .A0(n7075), .A1(n7076) );
  inv01 U3606 ( .Y(n7093), .A(n7101) );
  nand02 U3607 ( .Y(n7102), .A0(n7078), .A1(n7080) );
  inv01 U3608 ( .Y(n7103), .A(n7102) );
  nand02 U3609 ( .Y(n7104), .A0(n7082), .A1(n7084) );
  inv01 U3610 ( .Y(n7105), .A(n7104) );
  nand02 U3611 ( .Y(n7106), .A0(n7103), .A1(n7105) );
  inv01 U3612 ( .Y(n7070), .A(n7106) );
  nand02 U3613 ( .Y(n7107), .A0(n7086), .A1(n7088) );
  inv01 U3614 ( .Y(n7108), .A(n7107) );
  nand02 U3615 ( .Y(n7109), .A0(n7090), .A1(n7092) );
  inv01 U3616 ( .Y(n7110), .A(n7109) );
  nand02 U3617 ( .Y(n7111), .A0(n7108), .A1(n7110) );
  inv01 U3618 ( .Y(n7071), .A(n7111) );
  inv01 U3619 ( .Y(n8570), .A(n7112) );
  nor02 U3620 ( .Y(n7113), .A0(n8576), .A1(n7114) );
  nor02 U3621 ( .Y(n7115), .A0(n8576), .A1(n7116) );
  nor02 U3622 ( .Y(n7117), .A0(n8576), .A1(n7118) );
  nor02 U3623 ( .Y(n7119), .A0(n8576), .A1(n7120) );
  nor02 U3624 ( .Y(n7121), .A0(n8344), .A1(n7122) );
  nor02 U3625 ( .Y(n7123), .A0(n8344), .A1(n7124) );
  nor02 U3626 ( .Y(n7125), .A0(n8344), .A1(n7126) );
  nor02 U3627 ( .Y(n7127), .A0(n8344), .A1(n7128) );
  nor02 U3628 ( .Y(n7112), .A0(n7129), .A1(n7130) );
  nor02 U3629 ( .Y(n7131), .A0(n8572), .A1(n8574) );
  inv01 U3630 ( .Y(n7114), .A(n7131) );
  nor02 U3631 ( .Y(n7132), .A0(n8571), .A1(n8574) );
  inv01 U3632 ( .Y(n7116), .A(n7132) );
  nor02 U3633 ( .Y(n7133), .A0(n8572), .A1(n8333) );
  inv01 U3634 ( .Y(n7118), .A(n7133) );
  nor02 U3635 ( .Y(n7134), .A0(n8571), .A1(n8333) );
  inv01 U3636 ( .Y(n7120), .A(n7134) );
  nor02 U3637 ( .Y(n7135), .A0(n8572), .A1(n8574) );
  inv01 U3638 ( .Y(n7122), .A(n7135) );
  nor02 U3639 ( .Y(n7136), .A0(n8571), .A1(n8574) );
  inv01 U3640 ( .Y(n7124), .A(n7136) );
  nor02 U3641 ( .Y(n7137), .A0(n8572), .A1(n8333) );
  inv01 U3642 ( .Y(n7126), .A(n7137) );
  nor02 U3643 ( .Y(n7138), .A0(n8571), .A1(n8333) );
  inv01 U3644 ( .Y(n7128), .A(n7138) );
  nor02 U3645 ( .Y(n7139), .A0(n7113), .A1(n7115) );
  inv01 U3646 ( .Y(n7140), .A(n7139) );
  nor02 U3647 ( .Y(n7141), .A0(n7117), .A1(n7119) );
  inv01 U3648 ( .Y(n7142), .A(n7141) );
  nor02 U3649 ( .Y(n7143), .A0(n7140), .A1(n7142) );
  inv01 U3650 ( .Y(n7129), .A(n7143) );
  nor02 U3651 ( .Y(n7144), .A0(n7121), .A1(n7123) );
  inv01 U3652 ( .Y(n7145), .A(n7144) );
  nor02 U3653 ( .Y(n7146), .A0(n7125), .A1(n7127) );
  inv01 U3654 ( .Y(n7147), .A(n7146) );
  nor02 U3655 ( .Y(n7148), .A0(n7145), .A1(n7147) );
  inv01 U3656 ( .Y(n7130), .A(n7148) );
  inv02 U3657 ( .Y(n8333), .A(n8332) );
  inv04 U3658 ( .Y(n8344), .A(n8342) );
  nand02 U3659 ( .Y(n8691), .A0(n7149), .A1(n7150) );
  inv02 U3660 ( .Y(n7151), .A(n8693) );
  inv02 U3661 ( .Y(n7152), .A(n8692) );
  inv02 U3662 ( .Y(n7153), .A(n8614) );
  inv02 U3663 ( .Y(n7154), .A(n8352) );
  inv02 U3664 ( .Y(n7155), .A(n8327) );
  inv02 U3665 ( .Y(n7156), .A(n8005) );
  nand02 U3666 ( .Y(n7157), .A0(n7153), .A1(n7158) );
  nand02 U3667 ( .Y(n7159), .A0(n7154), .A1(n7160) );
  nand02 U3668 ( .Y(n7161), .A0(n7155), .A1(n7162) );
  nand02 U3669 ( .Y(n7163), .A0(n7155), .A1(n7164) );
  nand02 U3670 ( .Y(n7165), .A0(n7156), .A1(n7166) );
  nand02 U3671 ( .Y(n7167), .A0(n7156), .A1(n7168) );
  nand02 U3672 ( .Y(n7169), .A0(n7156), .A1(n7170) );
  nand02 U3673 ( .Y(n7171), .A0(n7156), .A1(n7172) );
  nand02 U3674 ( .Y(n7173), .A0(n7151), .A1(n7152) );
  inv01 U3675 ( .Y(n7158), .A(n7173) );
  nand02 U3676 ( .Y(n7174), .A0(n7151), .A1(n7152) );
  inv01 U3677 ( .Y(n7160), .A(n7174) );
  nand02 U3678 ( .Y(n7175), .A0(n7151), .A1(n7153) );
  inv01 U3679 ( .Y(n7162), .A(n7175) );
  nand02 U3680 ( .Y(n7176), .A0(n7151), .A1(n7154) );
  inv01 U3681 ( .Y(n7164), .A(n7176) );
  nand02 U3682 ( .Y(n7177), .A0(n7152), .A1(n7153) );
  inv01 U3683 ( .Y(n7166), .A(n7177) );
  nand02 U3684 ( .Y(n7178), .A0(n7152), .A1(n7154) );
  inv01 U3685 ( .Y(n7168), .A(n7178) );
  nand02 U3686 ( .Y(n7179), .A0(n7153), .A1(n7155) );
  inv01 U3687 ( .Y(n7170), .A(n7179) );
  nand02 U3688 ( .Y(n7180), .A0(n7154), .A1(n7155) );
  inv01 U3689 ( .Y(n7172), .A(n7180) );
  nand02 U3690 ( .Y(n7181), .A0(n7157), .A1(n7159) );
  inv01 U3691 ( .Y(n7182), .A(n7181) );
  nand02 U3692 ( .Y(n7183), .A0(n7161), .A1(n7163) );
  inv01 U3693 ( .Y(n7184), .A(n7183) );
  nand02 U3694 ( .Y(n7185), .A0(n7182), .A1(n7184) );
  inv01 U3695 ( .Y(n7149), .A(n7185) );
  nand02 U3696 ( .Y(n7186), .A0(n7165), .A1(n7167) );
  inv01 U3697 ( .Y(n7187), .A(n7186) );
  nand02 U3698 ( .Y(n7188), .A0(n7169), .A1(n7171) );
  inv01 U3699 ( .Y(n7189), .A(n7188) );
  nand02 U3700 ( .Y(n7190), .A0(n7187), .A1(n7189) );
  inv01 U3701 ( .Y(n7150), .A(n7190) );
  nand02 U3702 ( .Y(n8652), .A0(n7191), .A1(n7192) );
  inv02 U3703 ( .Y(n7193), .A(n8320) );
  inv02 U3704 ( .Y(n7194), .A(n5607) );
  inv02 U3705 ( .Y(n7195), .A(n8163) );
  inv02 U3706 ( .Y(n7196), .A(n8307) );
  inv02 U3707 ( .Y(n7197), .A(n8615) );
  inv02 U3708 ( .Y(n7198), .A(n8654) );
  nand02 U3709 ( .Y(n7199), .A0(n7195), .A1(n7200) );
  nand02 U3710 ( .Y(n7201), .A0(n7196), .A1(n7202) );
  nand02 U3711 ( .Y(n7203), .A0(n7197), .A1(n7204) );
  nand02 U3712 ( .Y(n7205), .A0(n7197), .A1(n7206) );
  nand02 U3713 ( .Y(n7207), .A0(n7198), .A1(n7208) );
  nand02 U3714 ( .Y(n7209), .A0(n7198), .A1(n7210) );
  nand02 U3715 ( .Y(n7211), .A0(n7198), .A1(n7212) );
  nand02 U3716 ( .Y(n7213), .A0(n7198), .A1(n7214) );
  nand02 U3717 ( .Y(n7215), .A0(n7193), .A1(n7194) );
  inv01 U3718 ( .Y(n7200), .A(n7215) );
  nand02 U3719 ( .Y(n7216), .A0(n7193), .A1(n7194) );
  inv01 U3720 ( .Y(n7202), .A(n7216) );
  nand02 U3721 ( .Y(n7217), .A0(n7193), .A1(n7195) );
  inv01 U3722 ( .Y(n7204), .A(n7217) );
  nand02 U3723 ( .Y(n7218), .A0(n7193), .A1(n7196) );
  inv01 U3724 ( .Y(n7206), .A(n7218) );
  nand02 U3725 ( .Y(n7219), .A0(n7194), .A1(n7195) );
  inv01 U3726 ( .Y(n7208), .A(n7219) );
  nand02 U3727 ( .Y(n7220), .A0(n7194), .A1(n7196) );
  inv01 U3728 ( .Y(n7210), .A(n7220) );
  nand02 U3729 ( .Y(n7221), .A0(n7195), .A1(n7197) );
  inv01 U3730 ( .Y(n7212), .A(n7221) );
  nand02 U3731 ( .Y(n7222), .A0(n7196), .A1(n7197) );
  inv01 U3732 ( .Y(n7214), .A(n7222) );
  nand02 U3733 ( .Y(n7223), .A0(n7199), .A1(n7201) );
  inv01 U3734 ( .Y(n7224), .A(n7223) );
  nand02 U3735 ( .Y(n7225), .A0(n7203), .A1(n7205) );
  inv01 U3736 ( .Y(n7226), .A(n7225) );
  nand02 U3737 ( .Y(n7227), .A0(n7224), .A1(n7226) );
  inv01 U3738 ( .Y(n7191), .A(n7227) );
  nand02 U3739 ( .Y(n7228), .A0(n7207), .A1(n7209) );
  inv01 U3740 ( .Y(n7229), .A(n7228) );
  nand02 U3741 ( .Y(n7230), .A0(n7211), .A1(n7213) );
  inv01 U3742 ( .Y(n7231), .A(n7230) );
  nand02 U3743 ( .Y(n7232), .A0(n7229), .A1(n7231) );
  inv01 U3744 ( .Y(n7192), .A(n7232) );
  nand02 U3745 ( .Y(n8662), .A0(n7233), .A1(n7234) );
  inv02 U3746 ( .Y(n7235), .A(n5607) );
  inv02 U3747 ( .Y(n7236), .A(n8171) );
  inv02 U3748 ( .Y(n7237), .A(n8321) );
  inv02 U3749 ( .Y(n7238), .A(n8663) );
  inv02 U3750 ( .Y(n7239), .A(n8163) );
  inv02 U3751 ( .Y(n7240), .A(n8664) );
  nand02 U3752 ( .Y(n7241), .A0(n7237), .A1(n7242) );
  nand02 U3753 ( .Y(n7243), .A0(n7238), .A1(n7244) );
  nand02 U3754 ( .Y(n7245), .A0(n7239), .A1(n7246) );
  nand02 U3755 ( .Y(n7247), .A0(n7239), .A1(n7248) );
  nand02 U3756 ( .Y(n7249), .A0(n7240), .A1(n7250) );
  nand02 U3757 ( .Y(n7251), .A0(n7240), .A1(n7252) );
  nand02 U3758 ( .Y(n7253), .A0(n7240), .A1(n7254) );
  nand02 U3759 ( .Y(n7255), .A0(n7240), .A1(n7256) );
  nand02 U3760 ( .Y(n7257), .A0(n7235), .A1(n7236) );
  inv01 U3761 ( .Y(n7242), .A(n7257) );
  nand02 U3762 ( .Y(n7258), .A0(n7235), .A1(n7236) );
  inv01 U3763 ( .Y(n7244), .A(n7258) );
  nand02 U3764 ( .Y(n7259), .A0(n7235), .A1(n7237) );
  inv01 U3765 ( .Y(n7246), .A(n7259) );
  nand02 U3766 ( .Y(n7260), .A0(n7235), .A1(n7238) );
  inv01 U3767 ( .Y(n7248), .A(n7260) );
  nand02 U3768 ( .Y(n7261), .A0(n7236), .A1(n7237) );
  inv01 U3769 ( .Y(n7250), .A(n7261) );
  nand02 U3770 ( .Y(n7262), .A0(n7236), .A1(n7238) );
  inv01 U3771 ( .Y(n7252), .A(n7262) );
  nand02 U3772 ( .Y(n7263), .A0(n7237), .A1(n7239) );
  inv01 U3773 ( .Y(n7254), .A(n7263) );
  nand02 U3774 ( .Y(n7264), .A0(n7238), .A1(n7239) );
  inv01 U3775 ( .Y(n7256), .A(n7264) );
  nand02 U3776 ( .Y(n7265), .A0(n7241), .A1(n7243) );
  inv01 U3777 ( .Y(n7266), .A(n7265) );
  nand02 U3778 ( .Y(n7267), .A0(n7245), .A1(n7247) );
  inv01 U3779 ( .Y(n7268), .A(n7267) );
  nand02 U3780 ( .Y(n7269), .A0(n7266), .A1(n7268) );
  inv01 U3781 ( .Y(n7233), .A(n7269) );
  nand02 U3782 ( .Y(n7270), .A0(n7249), .A1(n7251) );
  inv01 U3783 ( .Y(n7271), .A(n7270) );
  nand02 U3784 ( .Y(n7272), .A0(n7253), .A1(n7255) );
  inv01 U3785 ( .Y(n7273), .A(n7272) );
  nand02 U3786 ( .Y(n7274), .A0(n7271), .A1(n7273) );
  inv01 U3787 ( .Y(n7234), .A(n7274) );
  nand02 U3788 ( .Y(n8668), .A0(n7275), .A1(n7276) );
  inv02 U3789 ( .Y(n7277), .A(n8670) );
  inv02 U3790 ( .Y(n7278), .A(n8669) );
  inv02 U3791 ( .Y(n7279), .A(n8359) );
  inv02 U3792 ( .Y(n7280), .A(n8329) );
  inv02 U3793 ( .Y(n7281), .A(n8363) );
  nand02 U3794 ( .Y(n7282), .A0(n7278), .A1(n7283) );
  nand02 U3795 ( .Y(n7284), .A0(n7279), .A1(n7285) );
  nand02 U3796 ( .Y(n7286), .A0(n7280), .A1(n7287) );
  nand02 U3797 ( .Y(n7288), .A0(n7280), .A1(n7289) );
  nand02 U3798 ( .Y(n7290), .A0(n7281), .A1(n7291) );
  nand02 U3799 ( .Y(n7292), .A0(n7281), .A1(n7293) );
  nand02 U3800 ( .Y(n7294), .A0(n7281), .A1(n7295) );
  nand02 U3801 ( .Y(n7296), .A0(n7281), .A1(n7297) );
  nand02 U3802 ( .Y(n7298), .A0(n7277), .A1(n6821) );
  inv01 U3803 ( .Y(n7283), .A(n7298) );
  nand02 U3804 ( .Y(n7299), .A0(n7277), .A1(n6821) );
  inv01 U3805 ( .Y(n7285), .A(n7299) );
  nand02 U3806 ( .Y(n7300), .A0(n7277), .A1(n7278) );
  inv01 U3807 ( .Y(n7287), .A(n7300) );
  nand02 U3808 ( .Y(n7301), .A0(n7277), .A1(n7279) );
  inv01 U3809 ( .Y(n7289), .A(n7301) );
  nand02 U3810 ( .Y(n7302), .A0(n6821), .A1(n7278) );
  inv01 U3811 ( .Y(n7291), .A(n7302) );
  nand02 U3812 ( .Y(n7303), .A0(n6821), .A1(n7279) );
  inv01 U3813 ( .Y(n7293), .A(n7303) );
  nand02 U3814 ( .Y(n7304), .A0(n7278), .A1(n7280) );
  inv01 U3815 ( .Y(n7295), .A(n7304) );
  nand02 U3816 ( .Y(n7305), .A0(n7279), .A1(n7280) );
  inv01 U3817 ( .Y(n7297), .A(n7305) );
  nand02 U3818 ( .Y(n7306), .A0(n7282), .A1(n7284) );
  inv01 U3819 ( .Y(n7307), .A(n7306) );
  nand02 U3820 ( .Y(n7308), .A0(n7286), .A1(n7288) );
  inv01 U3821 ( .Y(n7309), .A(n7308) );
  nand02 U3822 ( .Y(n7310), .A0(n7307), .A1(n7309) );
  inv01 U3823 ( .Y(n7275), .A(n7310) );
  nand02 U3824 ( .Y(n7311), .A0(n7290), .A1(n7292) );
  inv01 U3825 ( .Y(n7312), .A(n7311) );
  nand02 U3826 ( .Y(n7313), .A0(n7294), .A1(n7296) );
  inv01 U3827 ( .Y(n7314), .A(n7313) );
  nand02 U3828 ( .Y(n7315), .A0(n7312), .A1(n7314) );
  inv01 U3829 ( .Y(n7276), .A(n7315) );
  nand02 U3830 ( .Y(n8649), .A0(n7316), .A1(n7317) );
  inv02 U3831 ( .Y(n7318), .A(n8574) );
  inv02 U3832 ( .Y(n7319), .A(n8651) );
  inv02 U3833 ( .Y(n7320), .A(n8650) );
  inv02 U3834 ( .Y(n7321), .A(n8359) );
  inv02 U3835 ( .Y(n7322), .A(n8363) );
  inv02 U3836 ( .Y(n7323), .A(n8329) );
  nand02 U3837 ( .Y(n7324), .A0(n7320), .A1(n7325) );
  nand02 U3838 ( .Y(n7326), .A0(n7321), .A1(n7327) );
  nand02 U3839 ( .Y(n7328), .A0(n7322), .A1(n7329) );
  nand02 U3840 ( .Y(n7330), .A0(n7322), .A1(n7331) );
  nand02 U3841 ( .Y(n7332), .A0(n7323), .A1(n7333) );
  nand02 U3842 ( .Y(n7334), .A0(n7323), .A1(n7335) );
  nand02 U3843 ( .Y(n7336), .A0(n7323), .A1(n7337) );
  nand02 U3844 ( .Y(n7338), .A0(n7323), .A1(n7339) );
  nand02 U3845 ( .Y(n7340), .A0(n7318), .A1(n7319) );
  inv01 U3846 ( .Y(n7325), .A(n7340) );
  nand02 U3847 ( .Y(n7341), .A0(n7318), .A1(n7319) );
  inv01 U3848 ( .Y(n7327), .A(n7341) );
  nand02 U3849 ( .Y(n7342), .A0(n7318), .A1(n7320) );
  inv01 U3850 ( .Y(n7329), .A(n7342) );
  nand02 U3851 ( .Y(n7343), .A0(n7318), .A1(n7321) );
  inv01 U3852 ( .Y(n7331), .A(n7343) );
  nand02 U3853 ( .Y(n7344), .A0(n7319), .A1(n7320) );
  inv01 U3854 ( .Y(n7333), .A(n7344) );
  nand02 U3855 ( .Y(n7345), .A0(n7319), .A1(n7321) );
  inv01 U3856 ( .Y(n7335), .A(n7345) );
  nand02 U3857 ( .Y(n7346), .A0(n7320), .A1(n7322) );
  inv01 U3858 ( .Y(n7337), .A(n7346) );
  nand02 U3859 ( .Y(n7347), .A0(n7321), .A1(n7322) );
  inv01 U3860 ( .Y(n7339), .A(n7347) );
  nand02 U3861 ( .Y(n7348), .A0(n7324), .A1(n7326) );
  inv01 U3862 ( .Y(n7349), .A(n7348) );
  nand02 U3863 ( .Y(n7350), .A0(n7328), .A1(n7330) );
  inv01 U3864 ( .Y(n7351), .A(n7350) );
  nand02 U3865 ( .Y(n7352), .A0(n7349), .A1(n7351) );
  inv01 U3866 ( .Y(n7316), .A(n7352) );
  nand02 U3867 ( .Y(n7353), .A0(n7332), .A1(n7334) );
  inv01 U3868 ( .Y(n7354), .A(n7353) );
  nand02 U3869 ( .Y(n7355), .A0(n7336), .A1(n7338) );
  inv01 U3870 ( .Y(n7356), .A(n7355) );
  nand02 U3871 ( .Y(n7357), .A0(n7354), .A1(n7356) );
  inv01 U3872 ( .Y(n7317), .A(n7357) );
  nand02 U3873 ( .Y(n8659), .A0(n7358), .A1(n7359) );
  inv02 U3874 ( .Y(n7360), .A(n8585) );
  inv02 U3875 ( .Y(n7361), .A(n8661) );
  inv02 U3876 ( .Y(n7362), .A(n8660) );
  inv02 U3877 ( .Y(n7363), .A(n8359) );
  inv02 U3878 ( .Y(n7364), .A(n8363) );
  inv02 U3879 ( .Y(n7365), .A(n8329) );
  nand02 U3880 ( .Y(n7366), .A0(n7362), .A1(n7367) );
  nand02 U3881 ( .Y(n7368), .A0(n7363), .A1(n7369) );
  nand02 U3882 ( .Y(n7370), .A0(n7364), .A1(n7371) );
  nand02 U3883 ( .Y(n7372), .A0(n7364), .A1(n7373) );
  nand02 U3884 ( .Y(n7374), .A0(n7365), .A1(n7375) );
  nand02 U3885 ( .Y(n7376), .A0(n7365), .A1(n7377) );
  nand02 U3886 ( .Y(n7378), .A0(n7365), .A1(n7379) );
  nand02 U3887 ( .Y(n7380), .A0(n7365), .A1(n7381) );
  nand02 U3888 ( .Y(n7382), .A0(n7360), .A1(n7361) );
  inv01 U3889 ( .Y(n7367), .A(n7382) );
  nand02 U3890 ( .Y(n7383), .A0(n7360), .A1(n7361) );
  inv01 U3891 ( .Y(n7369), .A(n7383) );
  nand02 U3892 ( .Y(n7384), .A0(n7360), .A1(n7362) );
  inv01 U3893 ( .Y(n7371), .A(n7384) );
  nand02 U3894 ( .Y(n7385), .A0(n7360), .A1(n7363) );
  inv01 U3895 ( .Y(n7373), .A(n7385) );
  nand02 U3896 ( .Y(n7386), .A0(n7361), .A1(n7362) );
  inv01 U3897 ( .Y(n7375), .A(n7386) );
  nand02 U3898 ( .Y(n7387), .A0(n7361), .A1(n7363) );
  inv01 U3899 ( .Y(n7377), .A(n7387) );
  nand02 U3900 ( .Y(n7388), .A0(n7362), .A1(n7364) );
  inv01 U3901 ( .Y(n7379), .A(n7388) );
  nand02 U3902 ( .Y(n7389), .A0(n7363), .A1(n7364) );
  inv01 U3903 ( .Y(n7381), .A(n7389) );
  nand02 U3904 ( .Y(n7390), .A0(n7366), .A1(n7368) );
  inv01 U3905 ( .Y(n7391), .A(n7390) );
  nand02 U3906 ( .Y(n7392), .A0(n7370), .A1(n7372) );
  inv01 U3907 ( .Y(n7393), .A(n7392) );
  nand02 U3908 ( .Y(n7394), .A0(n7391), .A1(n7393) );
  inv01 U3909 ( .Y(n7358), .A(n7394) );
  nand02 U3910 ( .Y(n7395), .A0(n7374), .A1(n7376) );
  inv01 U3911 ( .Y(n7396), .A(n7395) );
  nand02 U3912 ( .Y(n7397), .A0(n7378), .A1(n7380) );
  inv01 U3913 ( .Y(n7398), .A(n7397) );
  nand02 U3914 ( .Y(n7399), .A0(n7396), .A1(n7398) );
  inv01 U3915 ( .Y(n7359), .A(n7399) );
  inv02 U3916 ( .Y(n8574), .A(n8652) );
  inv02 U3917 ( .Y(n8660), .A(n8050) );
  inv02 U3918 ( .Y(n8585), .A(n8662) );
  nand02 U3919 ( .Y(n8740), .A0(n7400), .A1(n7401) );
  inv02 U3920 ( .Y(n7402), .A(n8714) );
  inv02 U3921 ( .Y(n7403), .A(n8171) );
  inv02 U3922 ( .Y(n7404), .A(n8741) );
  inv02 U3923 ( .Y(n7405), .A(n8005) );
  inv02 U3924 ( .Y(n7406), .A(n8363) );
  inv02 U3925 ( .Y(n7407), .A(n8327) );
  nand02 U3926 ( .Y(n7408), .A0(n7404), .A1(n7409) );
  nand02 U3927 ( .Y(n7410), .A0(n7405), .A1(n7411) );
  nand02 U3928 ( .Y(n7412), .A0(n7406), .A1(n7413) );
  nand02 U3929 ( .Y(n7414), .A0(n7406), .A1(n7415) );
  nand02 U3930 ( .Y(n7416), .A0(n7407), .A1(n7417) );
  nand02 U3931 ( .Y(n7418), .A0(n7407), .A1(n7419) );
  nand02 U3932 ( .Y(n7420), .A0(n7407), .A1(n7421) );
  nand02 U3933 ( .Y(n7422), .A0(n7407), .A1(n7423) );
  nand02 U3934 ( .Y(n7424), .A0(n7402), .A1(n7403) );
  inv01 U3935 ( .Y(n7409), .A(n7424) );
  nand02 U3936 ( .Y(n7425), .A0(n7402), .A1(n7403) );
  inv01 U3937 ( .Y(n7411), .A(n7425) );
  nand02 U3938 ( .Y(n7426), .A0(n7402), .A1(n7404) );
  inv01 U3939 ( .Y(n7413), .A(n7426) );
  nand02 U3940 ( .Y(n7427), .A0(n7402), .A1(n7405) );
  inv01 U3941 ( .Y(n7415), .A(n7427) );
  nand02 U3942 ( .Y(n7428), .A0(n7403), .A1(n7404) );
  inv01 U3943 ( .Y(n7417), .A(n7428) );
  nand02 U3944 ( .Y(n7429), .A0(n7403), .A1(n7405) );
  inv01 U3945 ( .Y(n7419), .A(n7429) );
  nand02 U3946 ( .Y(n7430), .A0(n7404), .A1(n7406) );
  inv01 U3947 ( .Y(n7421), .A(n7430) );
  nand02 U3948 ( .Y(n7431), .A0(n7405), .A1(n7406) );
  inv01 U3949 ( .Y(n7423), .A(n7431) );
  nand02 U3950 ( .Y(n7432), .A0(n7408), .A1(n7410) );
  inv01 U3951 ( .Y(n7433), .A(n7432) );
  nand02 U3952 ( .Y(n7434), .A0(n7412), .A1(n7414) );
  inv01 U3953 ( .Y(n7435), .A(n7434) );
  nand02 U3954 ( .Y(n7436), .A0(n7433), .A1(n7435) );
  inv01 U3955 ( .Y(n7400), .A(n7436) );
  nand02 U3956 ( .Y(n7437), .A0(n7416), .A1(n7418) );
  inv01 U3957 ( .Y(n7438), .A(n7437) );
  nand02 U3958 ( .Y(n7439), .A0(n7420), .A1(n7422) );
  inv01 U3959 ( .Y(n7440), .A(n7439) );
  nand02 U3960 ( .Y(n7441), .A0(n7438), .A1(n7440) );
  inv01 U3961 ( .Y(n7401), .A(n7441) );
  inv01 U3962 ( .Y(n7442), .A(n8410) );
  or04 U3963 ( .Y(n7443), .A0(n8842), .A1(n8843), .A2(n8844), .A3(n8845) );
  inv01 U3964 ( .Y(n7444), .A(n7443) );
  or04 U3965 ( .Y(n7445), .A0(n8834), .A1(n8835), .A2(n8836), .A3(n8837) );
  inv01 U3966 ( .Y(n7446), .A(n7445) );
  nand02 U3967 ( .Y(n8715), .A0(n7447), .A1(n7448) );
  inv02 U3968 ( .Y(n7449), .A(n8597) );
  inv02 U3969 ( .Y(n7450), .A(n8672) );
  inv02 U3970 ( .Y(n7451), .A(n8595) );
  inv02 U3971 ( .Y(n7452), .A(n8348) );
  inv02 U3972 ( .Y(n7453), .A(n8338) );
  inv02 U3973 ( .Y(n7454), .A(n8352) );
  nand02 U3974 ( .Y(n7455), .A0(n7451), .A1(n7456) );
  nand02 U3975 ( .Y(n7457), .A0(n7452), .A1(n7458) );
  nand02 U3976 ( .Y(n7459), .A0(n7453), .A1(n7460) );
  nand02 U3977 ( .Y(n7461), .A0(n7453), .A1(n7462) );
  nand02 U3978 ( .Y(n7463), .A0(n7454), .A1(n7464) );
  nand02 U3979 ( .Y(n7465), .A0(n7454), .A1(n7466) );
  nand02 U3980 ( .Y(n7467), .A0(n7454), .A1(n7468) );
  nand02 U3981 ( .Y(n7469), .A0(n7454), .A1(n7470) );
  nand02 U3982 ( .Y(n7471), .A0(n7449), .A1(n7450) );
  inv01 U3983 ( .Y(n7456), .A(n7471) );
  nand02 U3984 ( .Y(n7472), .A0(n7449), .A1(n7450) );
  inv01 U3985 ( .Y(n7458), .A(n7472) );
  nand02 U3986 ( .Y(n7473), .A0(n7449), .A1(n7451) );
  inv01 U3987 ( .Y(n7460), .A(n7473) );
  nand02 U3988 ( .Y(n7474), .A0(n7449), .A1(n7452) );
  inv01 U3989 ( .Y(n7462), .A(n7474) );
  nand02 U3990 ( .Y(n7475), .A0(n7450), .A1(n7451) );
  inv01 U3991 ( .Y(n7464), .A(n7475) );
  nand02 U3992 ( .Y(n7476), .A0(n7450), .A1(n7452) );
  inv01 U3993 ( .Y(n7466), .A(n7476) );
  nand02 U3994 ( .Y(n7477), .A0(n7451), .A1(n7453) );
  inv01 U3995 ( .Y(n7468), .A(n7477) );
  nand02 U3996 ( .Y(n7478), .A0(n7452), .A1(n7453) );
  inv01 U3997 ( .Y(n7470), .A(n7478) );
  nand02 U3998 ( .Y(n7479), .A0(n7455), .A1(n7457) );
  inv01 U3999 ( .Y(n7480), .A(n7479) );
  nand02 U4000 ( .Y(n7481), .A0(n7459), .A1(n7461) );
  inv01 U4001 ( .Y(n7482), .A(n7481) );
  nand02 U4002 ( .Y(n7483), .A0(n7480), .A1(n7482) );
  inv01 U4003 ( .Y(n7447), .A(n7483) );
  nand02 U4004 ( .Y(n7484), .A0(n7463), .A1(n7465) );
  inv01 U4005 ( .Y(n7485), .A(n7484) );
  nand02 U4006 ( .Y(n7486), .A0(n7467), .A1(n7469) );
  inv01 U4007 ( .Y(n7487), .A(n7486) );
  nand02 U4008 ( .Y(n7488), .A0(n7485), .A1(n7487) );
  inv01 U4009 ( .Y(n7448), .A(n7488) );
  inv01 U4010 ( .Y(n8680), .A(n7489) );
  nor02 U4011 ( .Y(n7490), .A0(n5559), .A1(n7491) );
  nor02 U4012 ( .Y(n7492), .A0(n5559), .A1(n7493) );
  nor02 U4013 ( .Y(n7494), .A0(n5559), .A1(n7495) );
  nor02 U4014 ( .Y(n7496), .A0(n5559), .A1(n7497) );
  nor02 U4015 ( .Y(n7498), .A0(n8337), .A1(n7499) );
  nor02 U4016 ( .Y(n7500), .A0(n8337), .A1(n7501) );
  nor02 U4017 ( .Y(n7502), .A0(n8638), .A1(n7503) );
  nor02 U4018 ( .Y(n7504), .A0(n8337), .A1(n7505) );
  nor02 U4019 ( .Y(n7489), .A0(n7506), .A1(n7507) );
  nor02 U4020 ( .Y(n7508), .A0(n5554), .A1(n8657) );
  inv01 U4021 ( .Y(n7491), .A(n7508) );
  nor02 U4022 ( .Y(n7509), .A0(n8338), .A1(n8657) );
  inv01 U4023 ( .Y(n7493), .A(n7509) );
  nor02 U4024 ( .Y(n7510), .A0(n5555), .A1(n8359) );
  inv01 U4025 ( .Y(n7495), .A(n7510) );
  nor02 U4026 ( .Y(n7511), .A0(n8338), .A1(n8359) );
  inv01 U4027 ( .Y(n7497), .A(n7511) );
  nor02 U4028 ( .Y(n7512), .A0(n5554), .A1(n8657) );
  inv01 U4029 ( .Y(n7499), .A(n7512) );
  nor02 U4030 ( .Y(n7513), .A0(n8338), .A1(n8657) );
  inv01 U4031 ( .Y(n7501), .A(n7513) );
  nor02 U4032 ( .Y(n7514), .A0(n5553), .A1(n8359) );
  inv01 U4033 ( .Y(n7503), .A(n7514) );
  nor02 U4034 ( .Y(n7515), .A0(n8338), .A1(n8359) );
  inv01 U4035 ( .Y(n7505), .A(n7515) );
  nor02 U4036 ( .Y(n7516), .A0(n7490), .A1(n7492) );
  inv01 U4037 ( .Y(n7517), .A(n7516) );
  nor02 U4038 ( .Y(n7518), .A0(n7494), .A1(n7496) );
  inv01 U4039 ( .Y(n7519), .A(n7518) );
  nor02 U4040 ( .Y(n7520), .A0(n7517), .A1(n7519) );
  inv01 U4041 ( .Y(n7506), .A(n7520) );
  nor02 U4042 ( .Y(n7521), .A0(n7498), .A1(n7500) );
  inv01 U4043 ( .Y(n7522), .A(n7521) );
  nor02 U4044 ( .Y(n7523), .A0(n7502), .A1(n7504) );
  inv01 U4045 ( .Y(n7524), .A(n7523) );
  nor02 U4046 ( .Y(n7525), .A0(n7522), .A1(n7524) );
  inv01 U4047 ( .Y(n7507), .A(n7525) );
  inv04 U4048 ( .Y(n8348), .A(n8346) );
  inv02 U4049 ( .Y(n8654), .A(n8215) );
  nand02 U4050 ( .Y(n8726), .A0(n7526), .A1(n7527) );
  inv02 U4051 ( .Y(n7528), .A(n8589) );
  inv02 U4052 ( .Y(n7529), .A(n8588) );
  inv02 U4053 ( .Y(n7530), .A(n8587) );
  inv02 U4054 ( .Y(n7531), .A(n8351) );
  inv02 U4055 ( .Y(n7532), .A(n8347) );
  nand02 U4056 ( .Y(n7533), .A0(n7530), .A1(n7534) );
  nand02 U4057 ( .Y(n7535), .A0(n5965), .A1(n7536) );
  nand02 U4058 ( .Y(n7537), .A0(n7531), .A1(n7538) );
  nand02 U4059 ( .Y(n7539), .A0(n7531), .A1(n7540) );
  nand02 U4060 ( .Y(n7541), .A0(n7532), .A1(n7542) );
  nand02 U4061 ( .Y(n7543), .A0(n7532), .A1(n7544) );
  nand02 U4062 ( .Y(n7545), .A0(n7532), .A1(n7546) );
  nand02 U4063 ( .Y(n7547), .A0(n7532), .A1(n7548) );
  nand02 U4064 ( .Y(n7549), .A0(n7528), .A1(n7529) );
  inv01 U4065 ( .Y(n7534), .A(n7549) );
  nand02 U4066 ( .Y(n7550), .A0(n7528), .A1(n7529) );
  inv01 U4067 ( .Y(n7536), .A(n7550) );
  nand02 U4068 ( .Y(n7551), .A0(n7528), .A1(n7530) );
  inv01 U4069 ( .Y(n7538), .A(n7551) );
  nand02 U4070 ( .Y(n7552), .A0(n7528), .A1(n5965) );
  inv01 U4071 ( .Y(n7540), .A(n7552) );
  nand02 U4072 ( .Y(n7553), .A0(n7529), .A1(n7530) );
  inv01 U4073 ( .Y(n7542), .A(n7553) );
  nand02 U4074 ( .Y(n7554), .A0(n7529), .A1(n5965) );
  inv01 U4075 ( .Y(n7544), .A(n7554) );
  nand02 U4076 ( .Y(n7555), .A0(n7530), .A1(n7531) );
  inv01 U4077 ( .Y(n7546), .A(n7555) );
  nand02 U4078 ( .Y(n7556), .A0(n5965), .A1(n7531) );
  inv01 U4079 ( .Y(n7548), .A(n7556) );
  nand02 U4080 ( .Y(n7557), .A0(n7533), .A1(n7535) );
  inv01 U4081 ( .Y(n7558), .A(n7557) );
  nand02 U4082 ( .Y(n7559), .A0(n7537), .A1(n7539) );
  inv01 U4083 ( .Y(n7560), .A(n7559) );
  nand02 U4084 ( .Y(n7561), .A0(n7558), .A1(n7560) );
  inv01 U4085 ( .Y(n7526), .A(n7561) );
  nand02 U4086 ( .Y(n7562), .A0(n7541), .A1(n7543) );
  inv01 U4087 ( .Y(n7563), .A(n7562) );
  nand02 U4088 ( .Y(n7564), .A0(n7545), .A1(n7547) );
  inv01 U4089 ( .Y(n7565), .A(n7564) );
  nand02 U4090 ( .Y(n7566), .A0(n7563), .A1(n7565) );
  inv01 U4091 ( .Y(n7527), .A(n7566) );
  nand02 U4092 ( .Y(n8730), .A0(n7567), .A1(n7568) );
  inv02 U4093 ( .Y(n7569), .A(n8630) );
  inv02 U4094 ( .Y(n7570), .A(n8597) );
  inv02 U4095 ( .Y(n7571), .A(n8595) );
  inv02 U4096 ( .Y(n7572), .A(n8347) );
  inv02 U4097 ( .Y(n7573), .A(n8338) );
  nand02 U4098 ( .Y(n7574), .A0(n7571), .A1(n7575) );
  nand02 U4099 ( .Y(n7576), .A0(n5965), .A1(n7577) );
  nand02 U4100 ( .Y(n7578), .A0(n7572), .A1(n7579) );
  nand02 U4101 ( .Y(n7580), .A0(n7572), .A1(n7581) );
  nand02 U4102 ( .Y(n7582), .A0(n7573), .A1(n7583) );
  nand02 U4103 ( .Y(n7584), .A0(n7573), .A1(n7585) );
  nand02 U4104 ( .Y(n7586), .A0(n7573), .A1(n7587) );
  nand02 U4105 ( .Y(n7588), .A0(n7573), .A1(n7589) );
  nand02 U4106 ( .Y(n7590), .A0(n7569), .A1(n7570) );
  inv01 U4107 ( .Y(n7575), .A(n7590) );
  nand02 U4108 ( .Y(n7591), .A0(n7569), .A1(n7570) );
  inv01 U4109 ( .Y(n7577), .A(n7591) );
  nand02 U4110 ( .Y(n7592), .A0(n7569), .A1(n7571) );
  inv01 U4111 ( .Y(n7579), .A(n7592) );
  nand02 U4112 ( .Y(n7593), .A0(n7569), .A1(n5965) );
  inv01 U4113 ( .Y(n7581), .A(n7593) );
  nand02 U4114 ( .Y(n7594), .A0(n7570), .A1(n7571) );
  inv01 U4115 ( .Y(n7583), .A(n7594) );
  nand02 U4116 ( .Y(n7595), .A0(n7570), .A1(n5965) );
  inv01 U4117 ( .Y(n7585), .A(n7595) );
  nand02 U4118 ( .Y(n7596), .A0(n7571), .A1(n7572) );
  inv01 U4119 ( .Y(n7587), .A(n7596) );
  nand02 U4120 ( .Y(n7597), .A0(n5965), .A1(n7572) );
  inv01 U4121 ( .Y(n7589), .A(n7597) );
  nand02 U4122 ( .Y(n7598), .A0(n7574), .A1(n7576) );
  inv01 U4123 ( .Y(n7599), .A(n7598) );
  nand02 U4124 ( .Y(n7600), .A0(n7578), .A1(n7580) );
  inv01 U4125 ( .Y(n7601), .A(n7600) );
  nand02 U4126 ( .Y(n7602), .A0(n7599), .A1(n7601) );
  inv01 U4127 ( .Y(n7567), .A(n7602) );
  nand02 U4128 ( .Y(n7603), .A0(n7582), .A1(n7584) );
  inv01 U4129 ( .Y(n7604), .A(n7603) );
  nand02 U4130 ( .Y(n7605), .A0(n7586), .A1(n7588) );
  inv01 U4131 ( .Y(n7606), .A(n7605) );
  nand02 U4132 ( .Y(n7607), .A0(n7604), .A1(n7606) );
  inv01 U4133 ( .Y(n7568), .A(n7607) );
  nand02 U4134 ( .Y(n8600), .A0(n7608), .A1(n7609) );
  inv02 U4135 ( .Y(n7610), .A(n8604) );
  inv02 U4136 ( .Y(n7611), .A(n8603) );
  inv02 U4137 ( .Y(n7612), .A(n8601) );
  inv02 U4138 ( .Y(n7613), .A(n8363) );
  inv02 U4139 ( .Y(n7614), .A(n8347) );
  nand02 U4140 ( .Y(n7615), .A0(n7612), .A1(n7616) );
  nand02 U4141 ( .Y(n7617), .A0(n5965), .A1(n7618) );
  nand02 U4142 ( .Y(n7619), .A0(n7613), .A1(n7620) );
  nand02 U4143 ( .Y(n7621), .A0(n7613), .A1(n7622) );
  nand02 U4144 ( .Y(n7623), .A0(n7614), .A1(n7624) );
  nand02 U4145 ( .Y(n7625), .A0(n7614), .A1(n7626) );
  nand02 U4146 ( .Y(n7627), .A0(n7614), .A1(n7628) );
  nand02 U4147 ( .Y(n7629), .A0(n7614), .A1(n7630) );
  nand02 U4148 ( .Y(n7631), .A0(n7610), .A1(n7611) );
  inv01 U4149 ( .Y(n7616), .A(n7631) );
  nand02 U4150 ( .Y(n7632), .A0(n7610), .A1(n7611) );
  inv01 U4151 ( .Y(n7618), .A(n7632) );
  nand02 U4152 ( .Y(n7633), .A0(n7610), .A1(n7612) );
  inv01 U4153 ( .Y(n7620), .A(n7633) );
  nand02 U4154 ( .Y(n7634), .A0(n7610), .A1(n5965) );
  inv01 U4155 ( .Y(n7622), .A(n7634) );
  nand02 U4156 ( .Y(n7635), .A0(n7611), .A1(n7612) );
  inv01 U4157 ( .Y(n7624), .A(n7635) );
  nand02 U4158 ( .Y(n7636), .A0(n7611), .A1(n5965) );
  inv01 U4159 ( .Y(n7626), .A(n7636) );
  nand02 U4160 ( .Y(n7637), .A0(n7612), .A1(n7613) );
  inv01 U4161 ( .Y(n7628), .A(n7637) );
  nand02 U4162 ( .Y(n7638), .A0(n5965), .A1(n7613) );
  inv01 U4163 ( .Y(n7630), .A(n7638) );
  nand02 U4164 ( .Y(n7639), .A0(n7615), .A1(n7617) );
  inv01 U4165 ( .Y(n7640), .A(n7639) );
  nand02 U4166 ( .Y(n7641), .A0(n7619), .A1(n7621) );
  inv01 U4167 ( .Y(n7642), .A(n7641) );
  nand02 U4168 ( .Y(n7643), .A0(n7640), .A1(n7642) );
  inv01 U4169 ( .Y(n7608), .A(n7643) );
  nand02 U4170 ( .Y(n7644), .A0(n7623), .A1(n7625) );
  inv01 U4171 ( .Y(n7645), .A(n7644) );
  nand02 U4172 ( .Y(n7646), .A0(n7627), .A1(n7629) );
  inv01 U4173 ( .Y(n7647), .A(n7646) );
  nand02 U4174 ( .Y(n7648), .A0(n7645), .A1(n7647) );
  inv01 U4175 ( .Y(n7609), .A(n7648) );
  nand02 U4176 ( .Y(n8611), .A0(n7649), .A1(n7650) );
  inv02 U4177 ( .Y(n7651), .A(n8581) );
  inv02 U4178 ( .Y(n7652), .A(n8307) );
  inv02 U4179 ( .Y(n7653), .A(n8578) );
  inv02 U4180 ( .Y(n7654), .A(n8359) );
  inv02 U4181 ( .Y(n7655), .A(n8347) );
  nand02 U4182 ( .Y(n7656), .A0(n7653), .A1(n7657) );
  nand02 U4183 ( .Y(n7658), .A0(n5965), .A1(n7659) );
  nand02 U4184 ( .Y(n7660), .A0(n7654), .A1(n7661) );
  nand02 U4185 ( .Y(n7662), .A0(n7654), .A1(n7663) );
  nand02 U4186 ( .Y(n7664), .A0(n7655), .A1(n7665) );
  nand02 U4187 ( .Y(n7666), .A0(n7655), .A1(n7667) );
  nand02 U4188 ( .Y(n7668), .A0(n7655), .A1(n7669) );
  nand02 U4189 ( .Y(n7670), .A0(n7655), .A1(n7671) );
  nand02 U4190 ( .Y(n7672), .A0(n7651), .A1(n7652) );
  inv01 U4191 ( .Y(n7657), .A(n7672) );
  nand02 U4192 ( .Y(n7673), .A0(n7651), .A1(n7652) );
  inv01 U4193 ( .Y(n7659), .A(n7673) );
  nand02 U4194 ( .Y(n7674), .A0(n7651), .A1(n7653) );
  inv01 U4195 ( .Y(n7661), .A(n7674) );
  nand02 U4196 ( .Y(n7675), .A0(n7651), .A1(n5965) );
  inv01 U4197 ( .Y(n7663), .A(n7675) );
  nand02 U4198 ( .Y(n7676), .A0(n7652), .A1(n7653) );
  inv01 U4199 ( .Y(n7665), .A(n7676) );
  nand02 U4200 ( .Y(n7677), .A0(n7652), .A1(n5965) );
  inv01 U4201 ( .Y(n7667), .A(n7677) );
  nand02 U4202 ( .Y(n7678), .A0(n7653), .A1(n7654) );
  inv01 U4203 ( .Y(n7669), .A(n7678) );
  nand02 U4204 ( .Y(n7679), .A0(n5965), .A1(n7654) );
  inv01 U4205 ( .Y(n7671), .A(n7679) );
  nand02 U4206 ( .Y(n7680), .A0(n7656), .A1(n7658) );
  inv01 U4207 ( .Y(n7681), .A(n7680) );
  nand02 U4208 ( .Y(n7682), .A0(n7660), .A1(n7662) );
  inv01 U4209 ( .Y(n7683), .A(n7682) );
  nand02 U4210 ( .Y(n7684), .A0(n7681), .A1(n7683) );
  inv01 U4211 ( .Y(n7649), .A(n7684) );
  nand02 U4212 ( .Y(n7685), .A0(n7664), .A1(n7666) );
  inv01 U4213 ( .Y(n7686), .A(n7685) );
  nand02 U4214 ( .Y(n7687), .A0(n7668), .A1(n7670) );
  inv01 U4215 ( .Y(n7688), .A(n7687) );
  nand02 U4216 ( .Y(n7689), .A0(n7686), .A1(n7688) );
  inv01 U4217 ( .Y(n7650), .A(n7689) );
  inv04 U4218 ( .Y(n8347), .A(n8346) );
  inv02 U4219 ( .Y(n8581), .A(n8257) );
  nand02 U4220 ( .Y(n8716), .A0(n7690), .A1(n7691) );
  inv02 U4221 ( .Y(n7692), .A(n8604) );
  inv02 U4222 ( .Y(n7693), .A(n8603) );
  inv02 U4223 ( .Y(n7694), .A(n8601) );
  inv02 U4224 ( .Y(n7695), .A(n8352) );
  inv02 U4225 ( .Y(n7696), .A(n8338) );
  inv02 U4226 ( .Y(n7697), .A(n8344) );
  nand02 U4227 ( .Y(n7698), .A0(n7694), .A1(n7699) );
  nand02 U4228 ( .Y(n7700), .A0(n7695), .A1(n7701) );
  nand02 U4229 ( .Y(n7702), .A0(n7696), .A1(n7703) );
  nand02 U4230 ( .Y(n7704), .A0(n7696), .A1(n7705) );
  nand02 U4231 ( .Y(n7706), .A0(n7697), .A1(n7707) );
  nand02 U4232 ( .Y(n7708), .A0(n7697), .A1(n7709) );
  nand02 U4233 ( .Y(n7710), .A0(n7697), .A1(n7711) );
  nand02 U4234 ( .Y(n7712), .A0(n7697), .A1(n7713) );
  nand02 U4235 ( .Y(n7714), .A0(n7692), .A1(n7693) );
  inv01 U4236 ( .Y(n7699), .A(n7714) );
  nand02 U4237 ( .Y(n7715), .A0(n7692), .A1(n7693) );
  inv01 U4238 ( .Y(n7701), .A(n7715) );
  nand02 U4239 ( .Y(n7716), .A0(n7692), .A1(n7694) );
  inv01 U4240 ( .Y(n7703), .A(n7716) );
  nand02 U4241 ( .Y(n7717), .A0(n7692), .A1(n7695) );
  inv01 U4242 ( .Y(n7705), .A(n7717) );
  nand02 U4243 ( .Y(n7718), .A0(n7693), .A1(n7694) );
  inv01 U4244 ( .Y(n7707), .A(n7718) );
  nand02 U4245 ( .Y(n7719), .A0(n7693), .A1(n7695) );
  inv01 U4246 ( .Y(n7709), .A(n7719) );
  nand02 U4247 ( .Y(n7720), .A0(n7694), .A1(n7696) );
  inv01 U4248 ( .Y(n7711), .A(n7720) );
  nand02 U4249 ( .Y(n7721), .A0(n7695), .A1(n7696) );
  inv01 U4250 ( .Y(n7713), .A(n7721) );
  nand02 U4251 ( .Y(n7722), .A0(n7698), .A1(n7700) );
  inv01 U4252 ( .Y(n7723), .A(n7722) );
  nand02 U4253 ( .Y(n7724), .A0(n7702), .A1(n7704) );
  inv01 U4254 ( .Y(n7725), .A(n7724) );
  nand02 U4255 ( .Y(n7726), .A0(n7723), .A1(n7725) );
  inv01 U4256 ( .Y(n7690), .A(n7726) );
  nand02 U4257 ( .Y(n7727), .A0(n7706), .A1(n7708) );
  inv01 U4258 ( .Y(n7728), .A(n7727) );
  nand02 U4259 ( .Y(n7729), .A0(n7710), .A1(n7712) );
  inv01 U4260 ( .Y(n7730), .A(n7729) );
  nand02 U4261 ( .Y(n7731), .A0(n7728), .A1(n7730) );
  inv01 U4262 ( .Y(n7691), .A(n7731) );
  inv02 U4263 ( .Y(n8603), .A(n8300) );
  buf02 U4264 ( .Y(n7732), .A(n8757) );
  inv01 U4265 ( .Y(n8676), .A(n7733) );
  nor02 U4266 ( .Y(n7734), .A0(n8637), .A1(n7735) );
  nor02 U4267 ( .Y(n7736), .A0(n8637), .A1(n7737) );
  nor02 U4268 ( .Y(n7738), .A0(n8637), .A1(n7739) );
  nor02 U4269 ( .Y(n7740), .A0(n8637), .A1(n7741) );
  nor02 U4270 ( .Y(n7742), .A0(n8338), .A1(n7743) );
  nor02 U4271 ( .Y(n7744), .A0(n8338), .A1(n7745) );
  nor02 U4272 ( .Y(n7746), .A0(n8338), .A1(n7747) );
  nor02 U4273 ( .Y(n7748), .A0(n8338), .A1(n7749) );
  nor02 U4274 ( .Y(n7733), .A0(n7750), .A1(n7751) );
  nor02 U4275 ( .Y(n7752), .A0(n8677), .A1(n8642) );
  inv01 U4276 ( .Y(n7735), .A(n7752) );
  nor02 U4277 ( .Y(n7753), .A0(n8337), .A1(n8642) );
  inv01 U4278 ( .Y(n7737), .A(n7753) );
  nor02 U4279 ( .Y(n7754), .A0(n8677), .A1(n8359) );
  inv01 U4280 ( .Y(n7739), .A(n7754) );
  nor02 U4281 ( .Y(n7755), .A0(n8337), .A1(n8359) );
  inv01 U4282 ( .Y(n7741), .A(n7755) );
  nor02 U4283 ( .Y(n7756), .A0(n8677), .A1(n8642) );
  inv01 U4284 ( .Y(n7743), .A(n7756) );
  nor02 U4285 ( .Y(n7757), .A0(n8337), .A1(n8642) );
  inv01 U4286 ( .Y(n7745), .A(n7757) );
  inv01 U4287 ( .Y(n7747), .A(n7754) );
  nor02 U4288 ( .Y(n7758), .A0(n8337), .A1(n8359) );
  inv01 U4289 ( .Y(n7749), .A(n7758) );
  nor02 U4290 ( .Y(n7759), .A0(n7734), .A1(n7736) );
  inv01 U4291 ( .Y(n7760), .A(n7759) );
  nor02 U4292 ( .Y(n7761), .A0(n7738), .A1(n7740) );
  inv01 U4293 ( .Y(n7762), .A(n7761) );
  nor02 U4294 ( .Y(n7763), .A0(n7760), .A1(n7762) );
  inv01 U4295 ( .Y(n7750), .A(n7763) );
  nor02 U4296 ( .Y(n7764), .A0(n7742), .A1(n7744) );
  inv01 U4297 ( .Y(n7765), .A(n7764) );
  nor02 U4298 ( .Y(n7766), .A0(n7746), .A1(n7748) );
  inv01 U4299 ( .Y(n7767), .A(n7766) );
  nor02 U4300 ( .Y(n7768), .A0(n7765), .A1(n7767) );
  inv01 U4301 ( .Y(n7751), .A(n7768) );
  buf08 U4302 ( .Y(n8359), .A(n8608) );
  buf08 U4303 ( .Y(n8338), .A(n8641) );
  xor2 U4304 ( .Y(n7769), .A0(s_shr1_4_), .A1(n5597) );
  inv02 U4305 ( .Y(n7770), .A(n7769) );
  inv02 U4306 ( .Y(n8746), .A(s_shr1_5_) );
  buf02 U4307 ( .Y(n7771), .A(n8621) );
  inv02 U4308 ( .Y(n8473), .A(n7772) );
  nand02 U4309 ( .Y(n7772), .A0(n5507), .A1(n7773) );
  nand02 U4310 ( .Y(n7774), .A0(n8489), .A1(n8506) );
  inv01 U4311 ( .Y(n7773), .A(n7774) );
  inv02 U4312 ( .Y(n8477), .A(n7775) );
  nand02 U4313 ( .Y(n7775), .A0(n5530), .A1(n7776) );
  nand02 U4314 ( .Y(n7777), .A0(n8499), .A1(n8504) );
  inv01 U4315 ( .Y(n7776), .A(n7777) );
  inv01 U4316 ( .Y(n8484), .A(n7778) );
  inv01 U4317 ( .Y(n7779), .A(n5513) );
  inv01 U4318 ( .Y(n7780), .A(n8419) );
  inv01 U4319 ( .Y(n7781), .A(n8418) );
  inv01 U4320 ( .Y(n7782), .A(n8485) );
  nand02 U4321 ( .Y(n7778), .A0(n7783), .A1(n7784) );
  nand02 U4322 ( .Y(n7785), .A0(n7779), .A1(n7780) );
  inv01 U4323 ( .Y(n7783), .A(n7785) );
  nand02 U4324 ( .Y(n7786), .A0(n7781), .A1(n7782) );
  inv01 U4325 ( .Y(n7784), .A(n7786) );
  inv02 U4326 ( .Y(n8738), .A(s_shl1_0_) );
  xor2 U4327 ( .Y(n7787), .A0(n8168), .A1(n8717) );
  inv02 U4328 ( .Y(n7788), .A(n7787) );
  or04 U4329 ( .Y(n7789), .A0(s_opa_i_11_), .A1(n8527), .A2(s_opa_i_10_), .A3(
        s_opa_i_0_) );
  inv01 U4330 ( .Y(n7790), .A(n7789) );
  or04 U4331 ( .Y(n7791), .A0(s_opb_i_11_), .A1(n8538), .A2(s_opb_i_10_), .A3(
        s_opb_i_0_) );
  inv01 U4332 ( .Y(n7792), .A(n7791) );
  or04 U4333 ( .Y(n7793), .A0(n8794), .A1(s_fraco1_0_), .A2(s_rmndr_i_10_), 
        .A3(s_rmndr_i_0_) );
  inv01 U4334 ( .Y(n7794), .A(n7793) );
  nand02 U4335 ( .Y(n8617), .A0(n7795), .A1(n7796) );
  inv02 U4336 ( .Y(n7797), .A(n7771) );
  inv02 U4337 ( .Y(n7798), .A(n8620) );
  inv02 U4338 ( .Y(n7799), .A(n8334) );
  inv02 U4339 ( .Y(n7800), .A(n8619) );
  inv02 U4340 ( .Y(n7801), .A(n8618) );
  inv02 U4341 ( .Y(n7802), .A(n8343) );
  inv02 U4342 ( .Y(n7803), .A(n8327) );
  nand02 U4343 ( .Y(n7804), .A0(n7799), .A1(n7805) );
  nand02 U4344 ( .Y(n7806), .A0(n7800), .A1(n7807) );
  nand02 U4345 ( .Y(n7808), .A0(n7801), .A1(n7809) );
  nand02 U4346 ( .Y(n7810), .A0(n7802), .A1(n7811) );
  nand02 U4347 ( .Y(n7812), .A0(n7802), .A1(n7813) );
  nand02 U4348 ( .Y(n7814), .A0(n7802), .A1(n7815) );
  nand02 U4349 ( .Y(n7816), .A0(n7803), .A1(n7817) );
  nand02 U4350 ( .Y(n7818), .A0(n7803), .A1(n7819) );
  nand02 U4351 ( .Y(n7820), .A0(n7803), .A1(n7821) );
  nand02 U4352 ( .Y(n7822), .A0(n7803), .A1(n7823) );
  nand02 U4353 ( .Y(n7824), .A0(n7803), .A1(n7825) );
  nand02 U4354 ( .Y(n7826), .A0(n7803), .A1(n7827) );
  nand02 U4355 ( .Y(n7828), .A0(n7797), .A1(n7798) );
  inv01 U4356 ( .Y(n7805), .A(n7828) );
  nand02 U4357 ( .Y(n7829), .A0(n7797), .A1(n7798) );
  inv01 U4358 ( .Y(n7807), .A(n7829) );
  nand02 U4359 ( .Y(n7830), .A0(n7797), .A1(n7798) );
  inv01 U4360 ( .Y(n7809), .A(n7830) );
  nand02 U4361 ( .Y(n7831), .A0(n7797), .A1(n7799) );
  inv01 U4362 ( .Y(n7811), .A(n7831) );
  nand02 U4363 ( .Y(n7832), .A0(n7797), .A1(n7800) );
  inv01 U4364 ( .Y(n7813), .A(n7832) );
  nand02 U4365 ( .Y(n7833), .A0(n7797), .A1(n7801) );
  inv01 U4366 ( .Y(n7815), .A(n7833) );
  nand02 U4367 ( .Y(n7834), .A0(n7798), .A1(n7799) );
  inv01 U4368 ( .Y(n7817), .A(n7834) );
  nand02 U4369 ( .Y(n7835), .A0(n7798), .A1(n7800) );
  inv01 U4370 ( .Y(n7819), .A(n7835) );
  nand02 U4371 ( .Y(n7836), .A0(n7798), .A1(n7801) );
  inv01 U4372 ( .Y(n7821), .A(n7836) );
  nand02 U4373 ( .Y(n7837), .A0(n7799), .A1(n7802) );
  inv01 U4374 ( .Y(n7823), .A(n7837) );
  nand02 U4375 ( .Y(n7838), .A0(n7800), .A1(n7802) );
  inv01 U4376 ( .Y(n7825), .A(n7838) );
  nand02 U4377 ( .Y(n7839), .A0(n7801), .A1(n7802) );
  inv01 U4378 ( .Y(n7827), .A(n7839) );
  nand02 U4379 ( .Y(n7840), .A0(n7804), .A1(n7806) );
  inv01 U4380 ( .Y(n7841), .A(n7840) );
  nand02 U4381 ( .Y(n7842), .A0(n7808), .A1(n7841) );
  inv01 U4382 ( .Y(n7843), .A(n7842) );
  nand02 U4383 ( .Y(n7844), .A0(n7810), .A1(n7812) );
  inv01 U4384 ( .Y(n7845), .A(n7844) );
  nand02 U4385 ( .Y(n7846), .A0(n7814), .A1(n7845) );
  inv01 U4386 ( .Y(n7847), .A(n7846) );
  nand02 U4387 ( .Y(n7848), .A0(n7843), .A1(n7847) );
  inv01 U4388 ( .Y(n7795), .A(n7848) );
  nand02 U4389 ( .Y(n7849), .A0(n7816), .A1(n7818) );
  inv01 U4390 ( .Y(n7850), .A(n7849) );
  nand02 U4391 ( .Y(n7851), .A0(n7820), .A1(n7850) );
  inv01 U4392 ( .Y(n7852), .A(n7851) );
  nand02 U4393 ( .Y(n7853), .A0(n7822), .A1(n7824) );
  inv01 U4394 ( .Y(n7854), .A(n7853) );
  nand02 U4395 ( .Y(n7855), .A0(n7826), .A1(n7854) );
  inv01 U4396 ( .Y(n7856), .A(n7855) );
  nand02 U4397 ( .Y(n7857), .A0(n7852), .A1(n7856) );
  inv01 U4398 ( .Y(n7796), .A(n7857) );
  nand02 U4399 ( .Y(n8687), .A0(n7858), .A1(n7859) );
  inv02 U4400 ( .Y(n7860), .A(n8660) );
  inv02 U4401 ( .Y(n7861), .A(n7771) );
  inv02 U4402 ( .Y(n7862), .A(n8329) );
  inv02 U4403 ( .Y(n7863), .A(n8619) );
  inv02 U4404 ( .Y(n7864), .A(n8618) );
  inv02 U4405 ( .Y(n7865), .A(n8678) );
  inv02 U4406 ( .Y(n7866), .A(n8363) );
  nand02 U4407 ( .Y(n7867), .A0(n7862), .A1(n7868) );
  nand02 U4408 ( .Y(n7869), .A0(n7863), .A1(n7870) );
  nand02 U4409 ( .Y(n7871), .A0(n7864), .A1(n7872) );
  nand02 U4410 ( .Y(n7873), .A0(n7865), .A1(n7874) );
  nand02 U4411 ( .Y(n7875), .A0(n7865), .A1(n7876) );
  nand02 U4412 ( .Y(n7877), .A0(n7865), .A1(n7878) );
  nand02 U4413 ( .Y(n7879), .A0(n7866), .A1(n7880) );
  nand02 U4414 ( .Y(n7881), .A0(n7866), .A1(n7882) );
  nand02 U4415 ( .Y(n7883), .A0(n7866), .A1(n7884) );
  nand02 U4416 ( .Y(n7885), .A0(n7866), .A1(n7886) );
  nand02 U4417 ( .Y(n7887), .A0(n7866), .A1(n7888) );
  nand02 U4418 ( .Y(n7889), .A0(n7866), .A1(n7890) );
  nand02 U4419 ( .Y(n7891), .A0(n7860), .A1(n7861) );
  inv01 U4420 ( .Y(n7868), .A(n7891) );
  nand02 U4421 ( .Y(n7892), .A0(n7860), .A1(n7861) );
  inv01 U4422 ( .Y(n7870), .A(n7892) );
  nand02 U4423 ( .Y(n7893), .A0(n7860), .A1(n7861) );
  inv01 U4424 ( .Y(n7872), .A(n7893) );
  nand02 U4425 ( .Y(n7894), .A0(n7860), .A1(n7862) );
  inv01 U4426 ( .Y(n7874), .A(n7894) );
  nand02 U4427 ( .Y(n7895), .A0(n7860), .A1(n7863) );
  inv01 U4428 ( .Y(n7876), .A(n7895) );
  nand02 U4429 ( .Y(n7896), .A0(n7860), .A1(n7864) );
  inv01 U4430 ( .Y(n7878), .A(n7896) );
  nand02 U4431 ( .Y(n7897), .A0(n7861), .A1(n7862) );
  inv01 U4432 ( .Y(n7880), .A(n7897) );
  nand02 U4433 ( .Y(n7898), .A0(n7861), .A1(n7863) );
  inv01 U4434 ( .Y(n7882), .A(n7898) );
  nand02 U4435 ( .Y(n7899), .A0(n7861), .A1(n7864) );
  inv01 U4436 ( .Y(n7884), .A(n7899) );
  nand02 U4437 ( .Y(n7900), .A0(n7862), .A1(n7865) );
  inv01 U4438 ( .Y(n7886), .A(n7900) );
  nand02 U4439 ( .Y(n7901), .A0(n7863), .A1(n7865) );
  inv01 U4440 ( .Y(n7888), .A(n7901) );
  nand02 U4441 ( .Y(n7902), .A0(n7864), .A1(n7865) );
  inv01 U4442 ( .Y(n7890), .A(n7902) );
  nand02 U4443 ( .Y(n7903), .A0(n7867), .A1(n7869) );
  inv01 U4444 ( .Y(n7904), .A(n7903) );
  nand02 U4445 ( .Y(n7905), .A0(n7871), .A1(n7904) );
  inv01 U4446 ( .Y(n7906), .A(n7905) );
  nand02 U4447 ( .Y(n7907), .A0(n7873), .A1(n7875) );
  inv01 U4448 ( .Y(n7908), .A(n7907) );
  nand02 U4449 ( .Y(n7909), .A0(n7877), .A1(n7908) );
  inv01 U4450 ( .Y(n7910), .A(n7909) );
  nand02 U4451 ( .Y(n7911), .A0(n7906), .A1(n7910) );
  inv01 U4452 ( .Y(n7858), .A(n7911) );
  nand02 U4453 ( .Y(n7912), .A0(n7879), .A1(n7881) );
  inv01 U4454 ( .Y(n7913), .A(n7912) );
  nand02 U4455 ( .Y(n7914), .A0(n7883), .A1(n7913) );
  inv01 U4456 ( .Y(n7915), .A(n7914) );
  nand02 U4457 ( .Y(n7916), .A0(n7885), .A1(n7887) );
  inv01 U4458 ( .Y(n7917), .A(n7916) );
  nand02 U4459 ( .Y(n7918), .A0(n7889), .A1(n7917) );
  inv01 U4460 ( .Y(n7919), .A(n7918) );
  nand02 U4461 ( .Y(n7920), .A0(n7915), .A1(n7919) );
  inv01 U4462 ( .Y(n7859), .A(n7920) );
  or04 U4463 ( .Y(n7921), .A0(n8526), .A1(s_opa_i_14_), .A2(s_opa_i_16_), .A3(
        s_opa_i_15_) );
  inv01 U4464 ( .Y(n7922), .A(n7921) );
  or04 U4465 ( .Y(n7923), .A0(n8537), .A1(s_opb_i_14_), .A2(s_opb_i_16_), .A3(
        s_opb_i_15_) );
  inv01 U4466 ( .Y(n7924), .A(n7923) );
  inv02 U4467 ( .Y(n8618), .A(n5470) );
  inv02 U4468 ( .Y(n8619), .A(s_shl1_3_) );
  or04 U4469 ( .Y(n7925), .A0(n8793), .A1(s_rmndr_i_15_), .A2(s_rmndr_i_17_), 
        .A3(s_rmndr_i_16_) );
  inv01 U4470 ( .Y(n7926), .A(n7925) );
  or04 U4471 ( .Y(n7927), .A0(n8525), .A1(s_opa_i_1_), .A2(s_opa_i_21_), .A3(
        s_opa_i_20_) );
  inv01 U4472 ( .Y(n7928), .A(n7927) );
  or04 U4473 ( .Y(n7929), .A0(n8536), .A1(s_opb_i_1_), .A2(s_opb_i_21_), .A3(
        s_opb_i_20_) );
  inv01 U4474 ( .Y(n7930), .A(n7929) );
  or04 U4475 ( .Y(n7931), .A0(n8792), .A1(s_rmndr_i_21_), .A2(s_rmndr_i_23_), 
        .A3(s_rmndr_i_22_) );
  inv01 U4476 ( .Y(n7932), .A(n7931) );
  inv01 U4477 ( .Y(n8534), .A(n7933) );
  inv01 U4478 ( .Y(n7934), .A(n8518) );
  inv01 U4479 ( .Y(n7935), .A(s_opb_i_23_) );
  inv01 U4480 ( .Y(n7936), .A(s_opb_i_24_) );
  inv01 U4481 ( .Y(n7937), .A(s_opb_i_25_) );
  nand02 U4482 ( .Y(n7933), .A0(n7938), .A1(n7939) );
  nand02 U4483 ( .Y(n7940), .A0(n7934), .A1(n7935) );
  inv01 U4484 ( .Y(n7938), .A(n7940) );
  nand02 U4485 ( .Y(n7941), .A0(n7936), .A1(n7937) );
  inv01 U4486 ( .Y(n7939), .A(n7941) );
  or04 U4487 ( .Y(n7942), .A0(n8535), .A1(s_opb_i_4_), .A2(s_opb_i_6_), .A3(
        s_opb_i_5_) );
  inv01 U4488 ( .Y(n7943), .A(n7942) );
  or04 U4489 ( .Y(n7944), .A0(n8524), .A1(s_opa_i_4_), .A2(s_opa_i_6_), .A3(
        s_opa_i_5_) );
  inv01 U4490 ( .Y(n7945), .A(n7944) );
  inv01 U4491 ( .Y(n8523), .A(n7946) );
  inv01 U4492 ( .Y(n7947), .A(n8522) );
  inv01 U4493 ( .Y(n7948), .A(s_opa_i_23_) );
  inv01 U4494 ( .Y(n7949), .A(s_opa_i_24_) );
  inv01 U4495 ( .Y(n7950), .A(s_opa_i_25_) );
  nand02 U4496 ( .Y(n7946), .A0(n7951), .A1(n7952) );
  nand02 U4497 ( .Y(n7953), .A0(n7947), .A1(n7948) );
  inv01 U4498 ( .Y(n7951), .A(n7953) );
  nand02 U4499 ( .Y(n7954), .A0(n7949), .A1(n7950) );
  inv01 U4500 ( .Y(n7952), .A(n7954) );
  or04 U4501 ( .Y(n7955), .A0(n8791), .A1(s_rmndr_i_3_), .A2(s_rmndr_i_5_), 
        .A3(s_rmndr_i_4_) );
  inv01 U4502 ( .Y(n7956), .A(n7955) );
  inv01 U4503 ( .Y(n8539), .A(n7957) );
  inv01 U4504 ( .Y(n7958), .A(n5538) );
  inv01 U4505 ( .Y(n7959), .A(s_round) );
  inv01 U4506 ( .Y(n7960), .A(n8883) );
  nand02 U4507 ( .Y(n7957), .A0(n7960), .A1(n7961) );
  nand02 U4508 ( .Y(n7962), .A0(n7958), .A1(n7959) );
  inv01 U4509 ( .Y(n7961), .A(n7962) );
  inv02 U4510 ( .Y(n7963), .A(n8394) );
  inv08 U4511 ( .Y(n7964), .A(n7963) );
  inv01 U4512 ( .Y(n7965), .A(n7963) );
  inv02 U4513 ( .Y(n8422), .A(n7966) );
  nand02 U4514 ( .Y(n7966), .A0(s_qutnt_i[15]), .A1(n7967) );
  nand02 U4515 ( .Y(n7968), .A0(n5530), .A1(n8499) );
  inv01 U4516 ( .Y(n7967), .A(n7968) );
  inv02 U4517 ( .Y(n8395), .A(n8759) );
  or02 U4518 ( .Y(n7969), .A0(s_qutnt_i[26]), .A1(n8416) );
  inv02 U4519 ( .Y(n7970), .A(n7969) );
  nand02 U4520 ( .Y(n8714), .A0(n7971), .A1(n7972) );
  inv01 U4521 ( .Y(n7973), .A(n8323) );
  inv01 U4522 ( .Y(n7974), .A(n8688) );
  inv01 U4523 ( .Y(n7975), .A(n8275) );
  inv01 U4524 ( .Y(n7976), .A(n8689) );
  inv01 U4525 ( .Y(n7977), .A(n8328) );
  inv01 U4526 ( .Y(n7978), .A(n8742) );
  nand02 U4527 ( .Y(n7979), .A0(n7973), .A1(n7974) );
  nand02 U4528 ( .Y(n7980), .A0(n7975), .A1(n7976) );
  nand02 U4529 ( .Y(n7971), .A0(n7977), .A1(n7978) );
  nand02 U4530 ( .Y(n7981), .A0(n7979), .A1(n7980) );
  inv01 U4531 ( .Y(n7972), .A(n7981) );
  nand02 U4532 ( .Y(n8633), .A0(n7982), .A1(n7983) );
  inv01 U4533 ( .Y(n7984), .A(n8322) );
  inv01 U4534 ( .Y(n7985), .A(n8705) );
  inv01 U4535 ( .Y(n7986), .A(n8704) );
  inv01 U4536 ( .Y(n7987), .A(n8275) );
  inv01 U4537 ( .Y(n7988), .A(n8328) );
  inv01 U4538 ( .Y(n7989), .A(n8702) );
  nand02 U4539 ( .Y(n7990), .A0(n7984), .A1(n7985) );
  nand02 U4540 ( .Y(n7991), .A0(n7986), .A1(n7987) );
  nand02 U4541 ( .Y(n7982), .A0(n7988), .A1(n7989) );
  nand02 U4542 ( .Y(n7992), .A0(n7990), .A1(n7991) );
  inv01 U4543 ( .Y(n7983), .A(n7992) );
  nand02 U4544 ( .Y(n8692), .A0(n7993), .A1(n7994) );
  inv01 U4545 ( .Y(n7995), .A(n8328) );
  inv01 U4546 ( .Y(n7996), .A(n8709) );
  inv01 U4547 ( .Y(n7997), .A(n8322) );
  inv01 U4548 ( .Y(n7998), .A(n8683) );
  inv01 U4549 ( .Y(n7999), .A(n8275) );
  inv01 U4550 ( .Y(n8000), .A(n8681) );
  nand02 U4551 ( .Y(n8001), .A0(n7995), .A1(n7996) );
  nand02 U4552 ( .Y(n8002), .A0(n7997), .A1(n7998) );
  nand02 U4553 ( .Y(n7993), .A0(n7999), .A1(n8000) );
  nand02 U4554 ( .Y(n8003), .A0(n8001), .A1(n8002) );
  inv01 U4555 ( .Y(n7994), .A(n8003) );
  buf02 U4556 ( .Y(n8275), .A(n8703) );
  nand02 U4557 ( .Y(n8004), .A0(n8744), .A1(n8031) );
  inv02 U4558 ( .Y(n8005), .A(n8004) );
  inv01 U4559 ( .Y(n8650), .A(n8006) );
  nor02 U4560 ( .Y(n8007), .A0(n8478), .A1(n8377) );
  nor02 U4561 ( .Y(n8008), .A0(n8500), .A1(n8386) );
  inv01 U4562 ( .Y(n8009), .A(n8685) );
  nor02 U4563 ( .Y(n8006), .A0(n8009), .A1(n8010) );
  nor02 U4564 ( .Y(n8011), .A0(n8007), .A1(n8008) );
  inv01 U4565 ( .Y(n8010), .A(n8011) );
  inv01 U4566 ( .Y(n8614), .A(n8012) );
  nor02 U4567 ( .Y(n8013), .A0(n8508), .A1(n8376) );
  nor02 U4568 ( .Y(n8014), .A0(n8474), .A1(n8379) );
  inv01 U4569 ( .Y(n8015), .A(n8694) );
  nor02 U4570 ( .Y(n8012), .A0(n8015), .A1(n8016) );
  nor02 U4571 ( .Y(n8017), .A0(n8013), .A1(n8014) );
  inv01 U4572 ( .Y(n8016), .A(n8017) );
  inv01 U4573 ( .Y(n8644), .A(n8018) );
  nor02 U4574 ( .Y(n8019), .A0(n8500), .A1(n8377) );
  nor02 U4575 ( .Y(n8020), .A0(n8498), .A1(n8387) );
  inv01 U4576 ( .Y(n8021), .A(n5382) );
  nor02 U4577 ( .Y(n8018), .A0(n8021), .A1(n8022) );
  nor02 U4578 ( .Y(n8023), .A0(n8019), .A1(n8020) );
  inv01 U4579 ( .Y(n8022), .A(n8023) );
  inv01 U4580 ( .Y(n8607), .A(n8024) );
  nor02 U4581 ( .Y(n8025), .A0(n8507), .A1(n8376) );
  nor02 U4582 ( .Y(n8026), .A0(n8508), .A1(n8380) );
  inv01 U4583 ( .Y(n8027), .A(n5462) );
  nor02 U4584 ( .Y(n8024), .A0(n8027), .A1(n8028) );
  nor02 U4585 ( .Y(n8029), .A0(n8025), .A1(n8026) );
  inv01 U4586 ( .Y(n8028), .A(n8029) );
  buf02 U4587 ( .Y(n8030), .A(n8745) );
  buf02 U4588 ( .Y(n8031), .A(n8745) );
  nor02 U4589 ( .Y(n8033), .A0(n8474), .A1(n8376) );
  nor02 U4590 ( .Y(n8034), .A0(n8509), .A1(n8379) );
  inv01 U4591 ( .Y(n8035), .A(n5213) );
  nor02 U4592 ( .Y(n8032), .A0(n8035), .A1(n8036) );
  nor02 U4593 ( .Y(n8037), .A0(n8033), .A1(n8034) );
  inv01 U4594 ( .Y(n8036), .A(n8037) );
  buf04 U4595 ( .Y(n8379), .A(n8626) );
  inv02 U4596 ( .Y(n8474), .A(s_qutnt_i[7]) );
  nor02 U4597 ( .Y(n8039), .A0(n8489), .A1(n8376) );
  nor02 U4598 ( .Y(n8040), .A0(n8507), .A1(n8379) );
  inv01 U4599 ( .Y(n8041), .A(n5323) );
  nor02 U4600 ( .Y(n8038), .A0(n8041), .A1(n8042) );
  nor02 U4601 ( .Y(n8043), .A0(n8039), .A1(n8040) );
  inv01 U4602 ( .Y(n8042), .A(n8043) );
  nor02 U4603 ( .Y(n8045), .A0(n8503), .A1(n8377) );
  nor02 U4604 ( .Y(n8046), .A0(n8501), .A1(n8387) );
  inv01 U4605 ( .Y(n8047), .A(n5307) );
  nor02 U4606 ( .Y(n8044), .A0(n8047), .A1(n8048) );
  nor02 U4607 ( .Y(n8049), .A0(n8045), .A1(n8046) );
  inv01 U4608 ( .Y(n8048), .A(n8049) );
  nor02 U4609 ( .Y(n8051), .A0(n8501), .A1(n8377) );
  nor02 U4610 ( .Y(n8052), .A0(n8478), .A1(n8385) );
  inv01 U4611 ( .Y(n8053), .A(n5444) );
  nor02 U4612 ( .Y(n8050), .A0(n8053), .A1(n8054) );
  nor02 U4613 ( .Y(n8055), .A0(n8051), .A1(n8052) );
  inv01 U4614 ( .Y(n8054), .A(n8055) );
  inv02 U4615 ( .Y(n8478), .A(s_qutnt_i[19]) );
  inv02 U4616 ( .Y(n8421), .A(n8056) );
  nand02 U4617 ( .Y(n8056), .A0(s_qutnt_i[23]), .A1(n8057) );
  nand02 U4618 ( .Y(n8058), .A0(n5594), .A1(n8495) );
  inv01 U4619 ( .Y(n8057), .A(n8058) );
  inv02 U4620 ( .Y(n8424), .A(n8059) );
  nand02 U4621 ( .Y(n8059), .A0(n5595), .A1(n8060) );
  nand02 U4622 ( .Y(n8061), .A0(n8479), .A1(n8306) );
  inv01 U4623 ( .Y(n8060), .A(n8061) );
  inv02 U4624 ( .Y(n8718), .A(n8062) );
  nor02 U4625 ( .Y(n8063), .A0(n8479), .A1(n8376) );
  nor02 U4626 ( .Y(n8064), .A0(n8494), .A1(n8379) );
  inv01 U4627 ( .Y(n8065), .A(n5341) );
  nor02 U4628 ( .Y(n8062), .A0(n8065), .A1(n8066) );
  nor02 U4629 ( .Y(n8067), .A0(n8063), .A1(n8064) );
  inv01 U4630 ( .Y(n8066), .A(n8067) );
  inv02 U4631 ( .Y(n8494), .A(s_qutnt_i[24]) );
  inv02 U4632 ( .Y(n8479), .A(s_qutnt_i[25]) );
  nand02 U4633 ( .Y(n8068), .A0(n8327), .A1(n8698) );
  inv02 U4634 ( .Y(n8069), .A(n8068) );
  xor2 U4635 ( .Y(n8070), .A0(n8089), .A1(s_exp_10_i_8_) );
  inv02 U4636 ( .Y(n8071), .A(n8070) );
  nand02 U4637 ( .Y(n8605), .A0(n8072), .A1(n8073) );
  inv01 U4638 ( .Y(n8074), .A(s_shr1_2_) );
  inv08 U4639 ( .Y(n8075), .A(n8717) );
  inv01 U4640 ( .Y(n8076), .A(n8705) );
  inv01 U4641 ( .Y(n8077), .A(n8704) );
  nand02 U4642 ( .Y(n8078), .A0(n8074), .A1(n8075) );
  nand02 U4643 ( .Y(n8079), .A0(n8074), .A1(n8076) );
  nand02 U4644 ( .Y(n8080), .A0(n8075), .A1(n8077) );
  nand02 U4645 ( .Y(n8081), .A0(n8076), .A1(n8077) );
  nand02 U4646 ( .Y(n8082), .A0(n8078), .A1(n8079) );
  inv02 U4647 ( .Y(n8072), .A(n8082) );
  nand02 U4648 ( .Y(n8083), .A0(n8080), .A1(n8081) );
  inv02 U4649 ( .Y(n8073), .A(n8083) );
  inv02 U4650 ( .Y(n8705), .A(n8718) );
  nand02 U4651 ( .Y(n8744), .A0(n8084), .A1(n8085) );
  inv01 U4652 ( .Y(n8086), .A(s_shr1_5_) );
  inv01 U4653 ( .Y(n8087), .A(n8030) );
  inv01 U4654 ( .Y(n8088), .A(n8370) );
  nand02 U4655 ( .Y(n8084), .A0(n8086), .A1(n8087) );
  nand02 U4656 ( .Y(n8085), .A0(n8086), .A1(n8088) );
  buf02 U4657 ( .Y(n8089), .A(n8766) );
  buf02 U4658 ( .Y(n8090), .A(n8766) );
  inv02 U4659 ( .Y(n8572), .A(n8091) );
  nor02 U4660 ( .Y(n8092), .A0(n8494), .A1(n8376) );
  nor02 U4661 ( .Y(n8093), .A0(n8496), .A1(n8379) );
  inv01 U4662 ( .Y(n8094), .A(n5279) );
  nor02 U4663 ( .Y(n8091), .A0(n8094), .A1(n8095) );
  nor02 U4664 ( .Y(n8096), .A0(n8092), .A1(n8093) );
  inv01 U4665 ( .Y(n8095), .A(n8096) );
  inv02 U4666 ( .Y(n8683), .A(n8572) );
  inv02 U4667 ( .Y(n8589), .A(n8097) );
  nor02 U4668 ( .Y(n8098), .A0(n8496), .A1(n8376) );
  nor02 U4669 ( .Y(n8099), .A0(n8495), .A1(n8380) );
  inv01 U4670 ( .Y(n8100), .A(n5436) );
  nor02 U4671 ( .Y(n8097), .A0(n8100), .A1(n8101) );
  nor02 U4672 ( .Y(n8102), .A0(n8098), .A1(n8099) );
  inv01 U4673 ( .Y(n8101), .A(n8102) );
  inv02 U4674 ( .Y(n8688), .A(n8589) );
  inv02 U4675 ( .Y(n8496), .A(s_qutnt_i[23]) );
  inv02 U4676 ( .Y(n8673), .A(n8103) );
  nor02 U4677 ( .Y(n8104), .A0(n8505), .A1(n8377) );
  nor02 U4678 ( .Y(n8105), .A0(n8499), .A1(n8386) );
  inv01 U4679 ( .Y(n8106), .A(n5327) );
  nor02 U4680 ( .Y(n8103), .A0(n8106), .A1(n8107) );
  nor02 U4681 ( .Y(n8108), .A0(n8104), .A1(n8105) );
  inv01 U4682 ( .Y(n8107), .A(n8108) );
  inv02 U4683 ( .Y(n8596), .A(n8109) );
  nor02 U4684 ( .Y(n8110), .A0(n8499), .A1(n8376) );
  nor02 U4685 ( .Y(n8111), .A0(n8505), .A1(n8379) );
  inv01 U4686 ( .Y(n8112), .A(n5402) );
  nor02 U4687 ( .Y(n8109), .A0(n8112), .A1(n8113) );
  nor02 U4688 ( .Y(n8114), .A0(n8110), .A1(n8111) );
  inv01 U4689 ( .Y(n8113), .A(n8114) );
  inv02 U4690 ( .Y(n8576), .A(n8115) );
  nor02 U4691 ( .Y(n8116), .A0(n8486), .A1(n8376) );
  nor02 U4692 ( .Y(n8117), .A0(n8506), .A1(n8380) );
  inv01 U4693 ( .Y(n8118), .A(n5261) );
  nor02 U4694 ( .Y(n8115), .A0(n8118), .A1(n8119) );
  nor02 U4695 ( .Y(n8120), .A0(n8116), .A1(n8117) );
  inv01 U4696 ( .Y(n8119), .A(n8120) );
  buf04 U4697 ( .Y(n8380), .A(n8378) );
  inv02 U4698 ( .Y(n8610), .A(n8121) );
  nor02 U4699 ( .Y(n8122), .A0(n8505), .A1(n8376) );
  nor02 U4700 ( .Y(n8123), .A0(n8486), .A1(n8380) );
  inv01 U4701 ( .Y(n8124), .A(n5380) );
  nor02 U4702 ( .Y(n8121), .A0(n8124), .A1(n8125) );
  nor02 U4703 ( .Y(n8126), .A0(n8122), .A1(n8123) );
  inv01 U4704 ( .Y(n8125), .A(n8126) );
  inv02 U4705 ( .Y(n8486), .A(s_qutnt_i[12]) );
  inv02 U4706 ( .Y(n8505), .A(s_qutnt_i[13]) );
  inv02 U4707 ( .Y(n8586), .A(n8127) );
  nor02 U4708 ( .Y(n8128), .A0(n8506), .A1(n8376) );
  nor02 U4709 ( .Y(n8129), .A0(n8489), .A1(n8380) );
  inv01 U4710 ( .Y(n8130), .A(n5440) );
  nor02 U4711 ( .Y(n8127), .A0(n8130), .A1(n8131) );
  nor02 U4712 ( .Y(n8132), .A0(n8128), .A1(n8129) );
  inv01 U4713 ( .Y(n8131), .A(n8132) );
  inv02 U4714 ( .Y(n8489), .A(s_qutnt_i[10]) );
  inv02 U4715 ( .Y(n8665), .A(n8133) );
  nor02 U4716 ( .Y(n8134), .A0(n8499), .A1(n8377) );
  nor02 U4717 ( .Y(n8135), .A0(n8504), .A1(n8387) );
  inv01 U4718 ( .Y(n8136), .A(n5416) );
  nor02 U4719 ( .Y(n8133), .A0(n8136), .A1(n8137) );
  nor02 U4720 ( .Y(n8138), .A0(n8134), .A1(n8135) );
  inv01 U4721 ( .Y(n8137), .A(n8138) );
  inv02 U4722 ( .Y(n8657), .A(n8139) );
  nor02 U4723 ( .Y(n8140), .A0(n8504), .A1(n8377) );
  nor02 U4724 ( .Y(n8141), .A0(n8502), .A1(n8385) );
  inv01 U4725 ( .Y(n8142), .A(n8708) );
  nor02 U4726 ( .Y(n8139), .A0(n8142), .A1(n8143) );
  nor02 U4727 ( .Y(n8144), .A0(n8140), .A1(n8141) );
  inv01 U4728 ( .Y(n8143), .A(n8144) );
  inv02 U4729 ( .Y(n8642), .A(n8145) );
  nor02 U4730 ( .Y(n8146), .A0(n8502), .A1(n8377) );
  nor02 U4731 ( .Y(n8147), .A0(n8503), .A1(n8386) );
  inv01 U4732 ( .Y(n8148), .A(n8701) );
  nor02 U4733 ( .Y(n8145), .A0(n8148), .A1(n8149) );
  nor02 U4734 ( .Y(n8150), .A0(n8146), .A1(n8147) );
  inv01 U4735 ( .Y(n8149), .A(n8150) );
  inv02 U4736 ( .Y(n8499), .A(s_qutnt_i[14]) );
  inv02 U4737 ( .Y(n8502), .A(s_qutnt_i[16]) );
  inv02 U4738 ( .Y(n8664), .A(n8151) );
  nor02 U4739 ( .Y(n8152), .A0(n8377), .A1(n8492) );
  nor02 U4740 ( .Y(n8153), .A0(n8387), .A1(n8510) );
  inv01 U4741 ( .Y(n8154), .A(n8728) );
  nor02 U4742 ( .Y(n8151), .A0(n8154), .A1(n8155) );
  nor02 U4743 ( .Y(n8156), .A0(n8152), .A1(n8153) );
  inv01 U4744 ( .Y(n8155), .A(n8156) );
  inv02 U4745 ( .Y(n8579), .A(n8157) );
  nor02 U4746 ( .Y(n8158), .A0(n8479), .A1(n8722) );
  nor02 U4747 ( .Y(n8159), .A0(n8306), .A1(n8360) );
  nor02 U4748 ( .Y(n8157), .A0(n8158), .A1(n8159) );
  or02 U4749 ( .Y(n8160), .A0(n8400), .A1(n8760) );
  inv02 U4750 ( .Y(n8161), .A(n8160) );
  inv02 U4751 ( .Y(s_expo2[0]), .A(n5467) );
  or02 U4752 ( .Y(n8162), .A0(n8619), .A1(s_shl1_2_) );
  inv02 U4753 ( .Y(n8163), .A(n8162) );
  ao21 U4754 ( .Y(n8164), .A0(s_exp_10_i_3_), .A1(n8771), .B0(n5159) );
  inv01 U4755 ( .Y(n8165), .A(n8164) );
  inv01 U4756 ( .Y(n8167), .A(n8164) );
  inv01 U4757 ( .Y(n8166), .A(n8164) );
  buf02 U4758 ( .Y(n8168), .A(n8783) );
  buf02 U4759 ( .Y(n8169), .A(n8783) );
  or02 U4760 ( .Y(n8170), .A0(n8461), .A1(n8721) );
  inv02 U4761 ( .Y(n8171), .A(n8170) );
  buf02 U4762 ( .Y(n8172), .A(n8719) );
  inv02 U4763 ( .Y(n8410), .A(n8406) );
  inv02 U4764 ( .Y(n8578), .A(n8173) );
  nor02 U4765 ( .Y(n8174), .A0(n8500), .A1(n8376) );
  nor02 U4766 ( .Y(n8175), .A0(n8478), .A1(n8379) );
  inv01 U4767 ( .Y(n8176), .A(n5442) );
  nor02 U4768 ( .Y(n8173), .A0(n8176), .A1(n8177) );
  nor02 U4769 ( .Y(n8178), .A0(n8174), .A1(n8175) );
  inv01 U4770 ( .Y(n8177), .A(n8178) );
  inv02 U4771 ( .Y(n8672), .A(n8179) );
  nor02 U4772 ( .Y(n8180), .A0(n8511), .A1(n8377) );
  nor02 U4773 ( .Y(n8181), .A0(n8509), .A1(n8385) );
  inv01 U4774 ( .Y(n8182), .A(n5167) );
  nor02 U4775 ( .Y(n8179), .A0(n8182), .A1(n8183) );
  nor02 U4776 ( .Y(n8184), .A0(n8180), .A1(n8181) );
  inv01 U4777 ( .Y(n8183), .A(n8184) );
  inv02 U4778 ( .Y(n8601), .A(n8185) );
  nor02 U4779 ( .Y(n8186), .A0(n8498), .A1(n8376) );
  nor02 U4780 ( .Y(n8187), .A0(n8500), .A1(n8379) );
  inv01 U4781 ( .Y(n8188), .A(n5195) );
  nor02 U4782 ( .Y(n8185), .A0(n8188), .A1(n8189) );
  nor02 U4783 ( .Y(n8190), .A0(n8186), .A1(n8187) );
  inv01 U4784 ( .Y(n8189), .A(n8190) );
  inv02 U4785 ( .Y(n8588), .A(n8191) );
  nor02 U4786 ( .Y(n8192), .A0(n8478), .A1(n8376) );
  nor02 U4787 ( .Y(n8193), .A0(n8501), .A1(n8379) );
  inv01 U4788 ( .Y(n8194), .A(n8743) );
  nor02 U4789 ( .Y(n8191), .A0(n8194), .A1(n8195) );
  nor02 U4790 ( .Y(n8196), .A0(n8192), .A1(n8193) );
  inv01 U4791 ( .Y(n8195), .A(n8196) );
  inv02 U4792 ( .Y(n8500), .A(s_qutnt_i[20]) );
  inv02 U4793 ( .Y(n8498), .A(s_qutnt_i[21]) );
  inv02 U4794 ( .Y(n8677), .A(n8197) );
  nor02 U4795 ( .Y(n8198), .A0(n8508), .A1(n8377) );
  nor02 U4796 ( .Y(n8199), .A0(n8507), .A1(n8386) );
  inv01 U4797 ( .Y(n8200), .A(n8737) );
  nor02 U4798 ( .Y(n8197), .A0(n8200), .A1(n8201) );
  nor02 U4799 ( .Y(n8202), .A0(n8198), .A1(n8199) );
  inv01 U4800 ( .Y(n8201), .A(n8202) );
  inv02 U4801 ( .Y(n8637), .A(n8203) );
  nor02 U4802 ( .Y(n8204), .A0(n8486), .A1(n8377) );
  nor02 U4803 ( .Y(n8205), .A0(n8505), .A1(n8385) );
  inv01 U4804 ( .Y(n8206), .A(n5418) );
  nor02 U4805 ( .Y(n8203), .A0(n8206), .A1(n8207) );
  nor02 U4806 ( .Y(n8208), .A0(n8204), .A1(n8205) );
  inv01 U4807 ( .Y(n8207), .A(n8208) );
  inv02 U4808 ( .Y(n8597), .A(n8209) );
  nor02 U4809 ( .Y(n8210), .A0(n8495), .A1(n8376) );
  nor02 U4810 ( .Y(n8211), .A0(n8498), .A1(n8380) );
  inv01 U4811 ( .Y(n8212), .A(n5384) );
  nor02 U4812 ( .Y(n8209), .A0(n8212), .A1(n8213) );
  nor02 U4813 ( .Y(n8214), .A0(n8210), .A1(n8211) );
  inv01 U4814 ( .Y(n8213), .A(n8214) );
  nor02 U4815 ( .Y(n8216), .A0(n8474), .A1(n8377) );
  nor02 U4816 ( .Y(n8217), .A0(n8508), .A1(n8386) );
  inv01 U4817 ( .Y(n8218), .A(n8725) );
  nor02 U4818 ( .Y(n8215), .A0(n8218), .A1(n8219) );
  nor02 U4819 ( .Y(n8220), .A0(n8216), .A1(n8217) );
  inv02 U4820 ( .Y(n8219), .A(n8220) );
  inv02 U4821 ( .Y(n8663), .A(n8221) );
  nor02 U4822 ( .Y(n8222), .A0(n8509), .A1(n8377) );
  nor02 U4823 ( .Y(n8223), .A0(n8474), .A1(n8385) );
  inv01 U4824 ( .Y(n8224), .A(n5398) );
  nor02 U4825 ( .Y(n8221), .A0(n8224), .A1(n8225) );
  nor02 U4826 ( .Y(n8226), .A0(n8222), .A1(n8223) );
  inv01 U4827 ( .Y(n8225), .A(n8226) );
  inv02 U4828 ( .Y(n8674), .A(n8227) );
  nor02 U4829 ( .Y(n8228), .A0(n8507), .A1(n8377) );
  nor02 U4830 ( .Y(n8229), .A0(n8489), .A1(n8386) );
  inv01 U4831 ( .Y(n8230), .A(n5446) );
  nor02 U4832 ( .Y(n8227), .A0(n8230), .A1(n8231) );
  nor02 U4833 ( .Y(n8232), .A0(n8228), .A1(n8229) );
  inv01 U4834 ( .Y(n8231), .A(n8232) );
  inv02 U4835 ( .Y(n8508), .A(s_qutnt_i[8]) );
  inv02 U4836 ( .Y(n8507), .A(s_qutnt_i[9]) );
  inv02 U4837 ( .Y(n8592), .A(n8233) );
  nor02 U4838 ( .Y(n8234), .A0(n8501), .A1(n8376) );
  nor02 U4839 ( .Y(n8235), .A0(n8503), .A1(n8380) );
  inv01 U4840 ( .Y(n8236), .A(n5293) );
  nor02 U4841 ( .Y(n8233), .A0(n8236), .A1(n8237) );
  nor02 U4842 ( .Y(n8238), .A0(n8234), .A1(n8235) );
  inv01 U4843 ( .Y(n8237), .A(n8238) );
  inv02 U4844 ( .Y(n8501), .A(s_qutnt_i[18]) );
  inv02 U4845 ( .Y(n8587), .A(n8239) );
  nor02 U4846 ( .Y(n8240), .A0(n8306), .A1(n8380) );
  nor02 U4847 ( .Y(n8241), .A0(n8494), .A1(n8722) );
  nor02 U4848 ( .Y(n8242), .A0(n8479), .A1(n8360) );
  nor02 U4849 ( .Y(n8239), .A0(n8242), .A1(n8243) );
  nor02 U4850 ( .Y(n8244), .A0(n8240), .A1(n8241) );
  inv01 U4851 ( .Y(n8243), .A(n8244) );
  inv02 U4852 ( .Y(n8689), .A(n8587) );
  buf04 U4853 ( .Y(n8360), .A(n8627) );
  inv02 U4854 ( .Y(n8666), .A(n8245) );
  nor02 U4855 ( .Y(n8246), .A0(n8489), .A1(n8377) );
  nor02 U4856 ( .Y(n8247), .A0(n8506), .A1(n8387) );
  inv01 U4857 ( .Y(n8248), .A(n8729) );
  nor02 U4858 ( .Y(n8245), .A0(n8248), .A1(n8249) );
  nor02 U4859 ( .Y(n8250), .A0(n8246), .A1(n8247) );
  inv01 U4860 ( .Y(n8249), .A(n8250) );
  inv02 U4861 ( .Y(n8656), .A(n8251) );
  nor02 U4862 ( .Y(n8252), .A0(n8506), .A1(n8377) );
  nor02 U4863 ( .Y(n8253), .A0(n8486), .A1(n8387) );
  inv01 U4864 ( .Y(n8254), .A(n8724) );
  nor02 U4865 ( .Y(n8251), .A0(n8254), .A1(n8255) );
  nor02 U4866 ( .Y(n8256), .A0(n8252), .A1(n8253) );
  inv01 U4867 ( .Y(n8255), .A(n8256) );
  inv02 U4868 ( .Y(n8506), .A(s_qutnt_i[11]) );
  nor02 U4869 ( .Y(n8258), .A0(n8502), .A1(n8376) );
  nor02 U4870 ( .Y(n8259), .A0(n8504), .A1(n8380) );
  inv01 U4871 ( .Y(n8260), .A(n8723) );
  nor02 U4872 ( .Y(n8257), .A0(n8260), .A1(n8261) );
  nor02 U4873 ( .Y(n8262), .A0(n8258), .A1(n8259) );
  inv02 U4874 ( .Y(n8261), .A(n8262) );
  inv02 U4875 ( .Y(n8584), .A(n8263) );
  nor02 U4876 ( .Y(n8264), .A0(n8504), .A1(n8376) );
  nor02 U4877 ( .Y(n8265), .A0(n8499), .A1(n8380) );
  inv01 U4878 ( .Y(n8266), .A(n5309) );
  nor02 U4879 ( .Y(n8263), .A0(n8266), .A1(n8267) );
  nor02 U4880 ( .Y(n8268), .A0(n8264), .A1(n8265) );
  inv01 U4881 ( .Y(n8267), .A(n8268) );
  inv02 U4882 ( .Y(n8504), .A(s_qutnt_i[15]) );
  inv02 U4883 ( .Y(n8604), .A(n8269) );
  nor02 U4884 ( .Y(n8270), .A0(n8503), .A1(n8376) );
  nor02 U4885 ( .Y(n8271), .A0(n8502), .A1(n8380) );
  inv01 U4886 ( .Y(n8272), .A(n5277) );
  nor02 U4887 ( .Y(n8269), .A0(n8272), .A1(n8273) );
  nor02 U4888 ( .Y(n8274), .A0(n8270), .A1(n8271) );
  inv01 U4889 ( .Y(n8273), .A(n8274) );
  inv02 U4890 ( .Y(n8503), .A(s_qutnt_i[17]) );
  nand02 U4891 ( .Y(n8276), .A0(n5165), .A1(n8340) );
  inv02 U4892 ( .Y(n8277), .A(n8276) );
  or04 U4893 ( .Y(n8278), .A0(n8460), .A1(n8463), .A2(s_qutnt_i[0]), .A3(
        s_qutnt_i[1]) );
  inv02 U4894 ( .Y(n8279), .A(n8278) );
  nand02 U4895 ( .Y(n8280), .A0(n8329), .A1(n8320) );
  inv02 U4896 ( .Y(n8615), .A(n8282) );
  nor02 U4897 ( .Y(n8283), .A0(n8377), .A1(n8510) );
  nor02 U4898 ( .Y(n8284), .A0(n8385), .A1(n8493) );
  inv01 U4899 ( .Y(n8285), .A(n5366) );
  nor02 U4900 ( .Y(n8282), .A0(n8285), .A1(n8286) );
  nor02 U4901 ( .Y(n8287), .A0(n8283), .A1(n8284) );
  inv01 U4902 ( .Y(n8286), .A(n8287) );
  buf04 U4903 ( .Y(n8385), .A(n8645) );
  inv02 U4904 ( .Y(n8630), .A(n8288) );
  nor02 U4905 ( .Y(n8289), .A0(n8377), .A1(n8462) );
  nor02 U4906 ( .Y(n8290), .A0(n8386), .A1(n8492) );
  inv01 U4907 ( .Y(n8291), .A(n8731) );
  nor02 U4908 ( .Y(n8288), .A0(n8291), .A1(n8292) );
  nor02 U4909 ( .Y(n8293), .A0(n8289), .A1(n8290) );
  inv01 U4910 ( .Y(n8292), .A(n8293) );
  inv02 U4911 ( .Y(n8462), .A(s_qutnt_i[1]) );
  inv02 U4912 ( .Y(n8595), .A(n8294) );
  nor02 U4913 ( .Y(n8295), .A0(n8306), .A1(n8376) );
  nor02 U4914 ( .Y(n8296), .A0(n8479), .A1(n8379) );
  inv01 U4915 ( .Y(n8297), .A(n8732) );
  nor02 U4916 ( .Y(n8294), .A0(n8297), .A1(n8298) );
  nor02 U4917 ( .Y(n8299), .A0(n8295), .A1(n8296) );
  inv01 U4918 ( .Y(n8298), .A(n8299) );
  buf02 U4919 ( .Y(n8306), .A(n8392) );
  nor02 U4920 ( .Y(n8301), .A0(n8493), .A1(n8377) );
  nor02 U4921 ( .Y(n8302), .A0(n8511), .A1(n8387) );
  inv01 U4922 ( .Y(n8303), .A(n5177) );
  nor02 U4923 ( .Y(n8300), .A0(n8303), .A1(n8304) );
  nor02 U4924 ( .Y(n8305), .A0(n8301), .A1(n8302) );
  inv02 U4925 ( .Y(n8304), .A(n8305) );
  inv02 U4926 ( .Y(n8511), .A(s_qutnt_i[5]) );
  inv02 U4927 ( .Y(n8509), .A(s_qutnt_i[6]) );
  nor02 U4928 ( .Y(n8310), .A0(n8492), .A1(n8721) );
  nor02 U4929 ( .Y(n8311), .A0(n8386), .A1(n8462) );
  nor02 U4930 ( .Y(n8312), .A0(n8377), .A1(n8461) );
  nor02 U4931 ( .Y(n8309), .A0(n8312), .A1(n8313) );
  nor02 U4932 ( .Y(n8314), .A0(n8310), .A1(n8311) );
  inv01 U4933 ( .Y(n8313), .A(n8314) );
  inv02 U4934 ( .Y(n8461), .A(s_qutnt_i[0]) );
  buf04 U4935 ( .Y(n8386), .A(n8383) );
  inv02 U4936 ( .Y(n8721), .A(n8374) );
  inv04 U4937 ( .Y(n8515), .A(n5575) );
  inv01 U4938 ( .Y(n8315), .A(n5699) );
  inv01 U4939 ( .Y(n8316), .A(n8521) );
  inv01 U4940 ( .Y(n8317), .A(n8520) );
  nor02 U4941 ( .Y(n8319), .A0(n8315), .A1(n8316) );
  inv02 U4942 ( .Y(n8318), .A(n8319) );
  buf02 U4943 ( .Y(n8320), .A(n8655) );
  buf02 U4944 ( .Y(n8321), .A(n8655) );
  buf02 U4945 ( .Y(n8322), .A(n8682) );
  buf02 U4946 ( .Y(n8323), .A(n8682) );
  inv04 U4947 ( .Y(n8325), .A(n8324) );
  nand02 U4948 ( .Y(n8326), .A0(s_shr1_4_), .A1(n8744) );
  inv04 U4949 ( .Y(n8327), .A(n8326) );
  inv04 U4950 ( .Y(n8678), .A(n8172) );
  buf04 U4951 ( .Y(n8329), .A(n8636) );
  inv04 U4952 ( .Y(n8331), .A(n8330) );
  inv02 U4953 ( .Y(n8332), .A(n8573) );
  inv02 U4954 ( .Y(n8336), .A(n8332) );
  inv02 U4955 ( .Y(n8334), .A(n8332) );
  inv02 U4956 ( .Y(n8335), .A(n8332) );
  buf02 U4957 ( .Y(n8339), .A(n8393) );
  buf02 U4958 ( .Y(n8341), .A(n8393) );
  buf02 U4959 ( .Y(n8340), .A(n8393) );
  inv02 U4960 ( .Y(n8342), .A(n8575) );
  inv02 U4961 ( .Y(n8343), .A(n8342) );
  inv02 U4962 ( .Y(n8346), .A(n8577) );
  inv02 U4963 ( .Y(n8349), .A(n8580) );
  inv02 U4964 ( .Y(n8352), .A(n8349) );
  inv02 U4965 ( .Y(n8351), .A(n8349) );
  inv01 U4966 ( .Y(n8354), .A(n8606) );
  inv01 U4967 ( .Y(n8355), .A(n8172) );
  inv04 U4968 ( .Y(n8356), .A(n8717) );
  nand02 U4969 ( .Y(n8353), .A0(n8356), .A1(n8357) );
  nand02 U4970 ( .Y(n8358), .A0(n8354), .A1(n8355) );
  inv04 U4971 ( .Y(n8357), .A(n8358) );
  inv04 U4972 ( .Y(n8717), .A(s_shr1_2_) );
  inv02 U4973 ( .Y(n8606), .A(s_shr1_3_) );
  inv08 U4974 ( .Y(n8361), .A(n8360) );
  buf12 U4975 ( .Y(n8362), .A(n8512) );
  buf16 U4976 ( .Y(n8363), .A(n8602) );
  inv04 U4977 ( .Y(n8364), .A(n5161) );
  inv02 U4978 ( .Y(n8365), .A(n8364) );
  inv02 U4979 ( .Y(n8367), .A(n8364) );
  inv02 U4980 ( .Y(n8368), .A(n8629) );
  inv04 U4981 ( .Y(n8369), .A(n8368) );
  inv04 U4982 ( .Y(n8370), .A(n8368) );
  inv02 U4983 ( .Y(n8371), .A(n8647) );
  inv02 U4984 ( .Y(n8372), .A(n8371) );
  inv04 U4985 ( .Y(n8374), .A(n8371) );
  inv02 U4986 ( .Y(n8373), .A(n8371) );
  buf16 U4987 ( .Y(n8375), .A(n8542) );
  buf16 U4988 ( .Y(n8376), .A(n8628) );
  buf16 U4989 ( .Y(n8377), .A(n8646) );
  or02 U4990 ( .Y(n8378), .A0(n8785), .A1(s_shr1_0_) );
  buf16 U4991 ( .Y(n8382), .A(n8540) );
  or02 U4992 ( .Y(n8383), .A0(n8738), .A1(s_shl1_1_) );
  or02 U4993 ( .Y(n8384), .A0(n8738), .A1(s_shl1_1_) );
  inv04 U4994 ( .Y(n8553), .A(n8382) );
  nor02 U4995 ( .Y(n8468), .A0(n8422), .A1(n8419) );
  nor02 U4996 ( .Y(n8467), .A0(n8424), .A1(n8421) );
  nand02 U4997 ( .Y(n8466), .A0(s_qutnt_i[6]), .A1(n8279) );
  and02 U4998 ( .Y(n8388), .A0(n8462), .A1(n8463) );
  inv01 U4999 ( .Y(n8472), .A(n8426) );
  inv01 U5000 ( .Y(n8471), .A(n8433) );
  nor02 U5001 ( .Y(n8470), .A0(n8432), .A1(n5515) );
  nor02 U5002 ( .Y(n8455), .A0(n5513), .A1(n8418) );
  inv01 U5003 ( .Y(n8454), .A(n8422) );
  nor02 U5004 ( .Y(n8453), .A0(n8423), .A1(n8421) );
  nand02 U5005 ( .Y(n8452), .A0(s_qutnt_i[6]), .A1(n8279) );
  nand03 U5006 ( .Y(n8450), .A0(n8457), .A1(n8458), .A2(n8456) );
  and04 U5007 ( .Y(n8389), .A0(n8459), .A1(n8460), .A2(n8461), .A3(n8462) );
  inv01 U5008 ( .Y(n8457), .A(n8434) );
  inv01 U5009 ( .Y(n8456), .A(n8432) );
  nand03 U5010 ( .Y(n8437), .A0(n8439), .A1(n8440), .A2(n8438) );
  nor02 U5011 ( .Y(n8440), .A0(n8419), .A1(n8420) );
  nor02 U5012 ( .Y(n8439), .A0(n8421), .A1(n8423) );
  nor02 U5013 ( .Y(n8438), .A0(n8424), .A1(n8425) );
  nand03 U5014 ( .Y(n8436), .A0(n5565), .A1(n8442), .A2(n8441) );
  nor02 U5015 ( .Y(n8442), .A0(n8429), .A1(n8431) );
  inv01 U5016 ( .Y(n8441), .A(n5515) );
  nand03 U5017 ( .Y(n8444), .A0(n8446), .A1(n8447), .A2(n8445) );
  nor02 U5018 ( .Y(n8447), .A0(n5513), .A1(n8417) );
  inv01 U5019 ( .Y(n8446), .A(n8422) );
  nor02 U5020 ( .Y(n8445), .A0(n8424), .A1(n8425) );
  nand03 U5021 ( .Y(n8443), .A0(n8449), .A1(n5592), .A2(n8448) );
  nor02 U5022 ( .Y(n8449), .A0(n8430), .A1(n8431) );
  nor02 U5023 ( .Y(n8448), .A0(n5515), .A1(n8435) );
  and03 U5025 ( .Y(v_shl433_0_), .A0(n8391), .A1(n8306), .A2(n8071) );
  ao21 U5026 ( .Y(s_shr1482_5_), .A0(n5158), .A1(n8341), .B0(n8277) );
  ao21 U5027 ( .Y(s_shr1482_4_), .A0(n8396), .A1(n8339), .B0(n8277) );
  ao21 U5028 ( .Y(n8396), .A0(n5621), .A1(n8397), .B0(n7965) );
  nor02 U5029 ( .Y(n8394), .A0(n8397), .A1(n5621) );
  ao21 U5030 ( .Y(s_shr1482_3_), .A0(n8401), .A1(n8339), .B0(n8277) );
  ao21 U5031 ( .Y(n8401), .A0(n8402), .A1(n8403), .B0(n5168) );
  nor02 U5032 ( .Y(n8398), .A0(n8403), .A1(n8402) );
  inv01 U5033 ( .Y(n8403), .A(n8404) );
  xor2 U5034 ( .Y(n8402), .A0(n8166), .A1(n5561) );
  ao21 U5035 ( .Y(s_shr1482_2_), .A0(n8407), .A1(n8340), .B0(n8277) );
  ao21 U5036 ( .Y(n8407), .A0(n8408), .A1(n8409), .B0(n5169) );
  nor02 U5037 ( .Y(n8404), .A0(n8409), .A1(n8408) );
  ao21 U5038 ( .Y(s_shr1482_1_), .A0(n8412), .A1(n8340), .B0(n8277) );
  nand02 U5039 ( .Y(n8409), .A0(n7970), .A1(n8410) );
  ao21 U5040 ( .Y(s_shr1482_0_), .A0(n8413), .A1(n8341), .B0(n8277) );
  nand02 U5041 ( .Y(n8415), .A0(n8395), .A1(n8161) );
  ao21 U5042 ( .Y(n8413), .A0(n8416), .A1(s_qutnt_i[26]), .B0(n7970) );
  or02 U5043 ( .Y(s_r_zeros_4_), .A0(n8436), .A1(n8437) );
  or02 U5044 ( .Y(s_r_zeros_3_), .A0(n8443), .A1(n8444) );
  or02 U5045 ( .Y(s_r_zeros_2_), .A0(n8450), .A1(n8451) );
  nand04 U5046 ( .Y(n8451), .A0(n8455), .A1(n8453), .A2(n8454), .A3(n8452) );
  inv01 U5047 ( .Y(n8459), .A(n8463) );
  or02 U5048 ( .Y(s_r_zeros_1_), .A0(n8464), .A1(n8465) );
  nand04 U5049 ( .Y(n8465), .A0(n8466), .A1(n8467), .A2(n8468), .A3(n5163) );
  inv01 U5050 ( .Y(n8417), .A(n8469) );
  nand04 U5051 ( .Y(n8464), .A0(n8470), .A1(n8471), .A2(n8472), .A3(n5573) );
  and02 U5052 ( .Y(n8427), .A0(s_qutnt_i[14]), .A1(n5530) );
  and02 U5053 ( .Y(n8428), .A0(s_qutnt_i[12]), .A1(n8473) );
  and03 U5054 ( .Y(n8430), .A0(n5689), .A1(n8474), .A2(s_qutnt_i[8]) );
  and02 U5055 ( .Y(n8426), .A0(s_qutnt_i[10]), .A1(n5507) );
  and02 U5056 ( .Y(n8431), .A0(s_qutnt_i[24]), .A1(n8475) );
  and02 U5057 ( .Y(n8433), .A0(s_qutnt_i[18]), .A1(n8476) );
  and02 U5058 ( .Y(n8429), .A0(s_qutnt_i[16]), .A1(n8477) );
  and03 U5059 ( .Y(n8434), .A0(n5691), .A1(n8478), .A2(s_qutnt_i[20]) );
  and02 U5060 ( .Y(n8432), .A0(s_qutnt_i[22]), .A1(n5594) );
  inv01 U5061 ( .Y(n8435), .A(n8481) );
  nand03 U5062 ( .Y(s_r_zeros_0_), .A0(n8482), .A1(n8483), .A2(n8484) );
  and02 U5063 ( .Y(n8419), .A0(s_qutnt_i[19]), .A1(n5691) );
  and02 U5064 ( .Y(n8418), .A0(s_qutnt_i[7]), .A1(n5689) );
  ao21 U5065 ( .Y(n8485), .A0(n8487), .A1(n8461), .B0(n8488) );
  nand02 U5066 ( .Y(n8488), .A0(n8481), .A1(n8469) );
  nand03 U5067 ( .Y(n8469), .A0(n5507), .A1(n8489), .A2(s_qutnt_i[11]) );
  nand02 U5068 ( .Y(n8481), .A0(s_qutnt_i[9]), .A1(n8490) );
  ao21 U5069 ( .Y(n8487), .A0(n8491), .A1(n8492), .B0(s_qutnt_i[1]) );
  ao21 U5070 ( .Y(n8491), .A0(s_qutnt_i[5]), .A1(n8493), .B0(s_qutnt_i[3]) );
  and02 U5071 ( .Y(n8425), .A0(s_qutnt_i[25]), .A1(n5596) );
  and02 U5072 ( .Y(n8480), .A0(n8475), .A1(n8494) );
  and03 U5073 ( .Y(n8475), .A0(n8495), .A1(n8496), .A2(n5594) );
  and02 U5074 ( .Y(n8423), .A0(s_qutnt_i[21]), .A1(n8497) );
  and03 U5075 ( .Y(n8497), .A0(n8478), .A1(n8500), .A2(n5691) );
  and03 U5076 ( .Y(n8476), .A0(n8502), .A1(n8503), .A2(n8477) );
  and03 U5077 ( .Y(n8420), .A0(n8477), .A1(n8502), .A2(s_qutnt_i[17]) );
  and03 U5078 ( .Y(n8490), .A0(n8474), .A1(n8508), .A2(n5689) );
  nand02 U5079 ( .Y(n8463), .A0(n8510), .A1(n8492) );
  nand02 U5080 ( .Y(n8460), .A0(n8511), .A1(n8493) );
  or02 U5081 ( .Y(s_output_o_31_), .A0(n8513), .A1(s_sign_i) );
  ao21 U5082 ( .Y(s_output_o_30_), .A0(n8331), .A1(s_expo3_7_), .B0(n8515) );
  ao21 U5083 ( .Y(s_output_o_29_), .A0(n8331), .A1(s_expo3_6_), .B0(n8515) );
  ao21 U5084 ( .Y(s_output_o_28_), .A0(n8331), .A1(s_expo3_5_), .B0(n8515) );
  ao21 U5085 ( .Y(s_output_o_27_), .A0(n8331), .A1(s_expo3_4_), .B0(n8515) );
  ao21 U5086 ( .Y(s_output_o_26_), .A0(n8331), .A1(s_expo3_3_), .B0(n8515) );
  ao21 U5087 ( .Y(s_output_o_25_), .A0(n8331), .A1(s_expo3_2_), .B0(n8515) );
  ao21 U5088 ( .Y(s_output_o_24_), .A0(n8331), .A1(s_expo3_1_), .B0(n8515) );
  ao21 U5089 ( .Y(s_output_o_23_), .A0(n8331), .A1(s_expo3_0_), .B0(n8515) );
  ao21 U5090 ( .Y(s_output_o_22_), .A0(s_fraco2_22_), .A1(n8331), .B0(n8513)
         );
  ao221 U5091 ( .Y(n8513), .A0(n5537), .A1(n8517), .B0(n5531), .B1(n8519), 
        .C0(n5469) );
  inv01 U5092 ( .Y(n8512), .A(n8331) );
  nor02 U5093 ( .Y(n8514), .A0(n8515), .A1(n8516) );
  and04 U5094 ( .Y(n8516), .A0(n8828), .A1(n8829), .A2(n5609), .A3(n8523) );
  nand04 U5095 ( .Y(n8522), .A0(n7790), .A1(n7922), .A2(n7928), .A3(n7945) );
  nand03 U5096 ( .Y(n8524), .A0(n8818), .A1(n8819), .A2(n8817) );
  nand03 U5097 ( .Y(n8525), .A0(n8821), .A1(n8822), .A2(n8820) );
  nand03 U5098 ( .Y(n8526), .A0(n8824), .A1(n8825), .A2(n8823) );
  nand02 U5099 ( .Y(n8527), .A0(n8826), .A1(n8827) );
  inv01 U5100 ( .Y(n8517), .A(n8528) );
  inv01 U5101 ( .Y(n8530), .A(n8521) );
  nand02 U5102 ( .Y(n8521), .A0(n6628), .A1(n7444) );
  nand02 U5103 ( .Y(n8533), .A0(n5694), .A1(n8859) );
  nand04 U5104 ( .Y(n8528), .A0(n8857), .A1(n8858), .A2(n5611), .A3(n8534) );
  nand04 U5105 ( .Y(n8518), .A0(n7792), .A1(n7924), .A2(n7930), .A3(n7943) );
  nand03 U5106 ( .Y(n8535), .A0(n8847), .A1(n8848), .A2(n8846) );
  nand03 U5107 ( .Y(n8536), .A0(n8850), .A1(n8851), .A2(n8849) );
  nand03 U5108 ( .Y(n8537), .A0(n8853), .A1(n8854), .A2(n8852) );
  nand02 U5109 ( .Y(n8538), .A0(n8855), .A1(n8856) );
  and04 U5110 ( .Y(n8532), .A0(s_expo3_0_), .A1(s_expo3_1_), .A2(s_expo3_2_), 
        .A3(s_expo3_3_) );
  and04 U5111 ( .Y(n8531), .A0(s_expo3_4_), .A1(s_expo3_5_), .A2(s_expo3_6_), 
        .A3(s_expo3_7_) );
  inv01 U5112 ( .Y(n8519), .A(n8520) );
  nand02 U5113 ( .Y(n8520), .A0(n6626), .A1(n7446) );
  inv01 U5114 ( .Y(n8529), .A(n8539) );
  inv01 U5115 ( .Y(n8543), .A(n____return3241_9_) );
  inv01 U5116 ( .Y(n8545), .A(n____return3241_8_) );
  inv01 U5117 ( .Y(n8546), .A(n____return3241_7_) );
  inv01 U5118 ( .Y(n8547), .A(n____return3241_6_) );
  inv01 U5119 ( .Y(n8548), .A(n____return3241_5_) );
  inv01 U5120 ( .Y(n8549), .A(n____return3241_4_) );
  inv01 U5121 ( .Y(n8550), .A(n____return3241_3_) );
  inv01 U5122 ( .Y(n8554), .A(n____return3241_22_) );
  inv01 U5123 ( .Y(n8555), .A(n____return3241_21_) );
  inv01 U5124 ( .Y(n8557), .A(n____return3241_1_) );
  inv01 U5125 ( .Y(n8551), .A(n____return3241_2_) );
  inv01 U5126 ( .Y(n8556), .A(n____return3241_20_) );
  inv01 U5127 ( .Y(n8558), .A(n____return3241_19_) );
  inv01 U5128 ( .Y(n8559), .A(n____return3241_18_) );
  inv01 U5129 ( .Y(n8560), .A(n____return3241_17_) );
  inv01 U5130 ( .Y(n8562), .A(n____return3241_15_) );
  inv01 U5131 ( .Y(n8563), .A(n____return3241_14_) );
  inv01 U5132 ( .Y(n8564), .A(n____return3241_13_) );
  inv01 U5133 ( .Y(n8565), .A(n____return3241_12_) );
  inv01 U5134 ( .Y(n8541), .A(n____return3241_10_) );
  inv01 U5135 ( .Y(n8566), .A(n____return3241_11_) );
  ao21 U5136 ( .Y(s_fraco23289_0_), .A0(n5556), .A1(s_fraco1_3_), .B0(n8568)
         );
  ao22 U5137 ( .Y(n8568), .A0(n____return3241_0_), .A1(n8552), .B0(
        n____return3241_1_), .B1(n8553) );
  inv01 U5138 ( .Y(n8552), .A(n8375) );
  nand02 U5139 ( .Y(n8542), .A0(n8381), .A1(n8382) );
  nand02 U5140 ( .Y(s_fraco1812_9_), .A0(n8569), .A1(n8570) );
  nand02 U5141 ( .Y(s_fraco1812_8_), .A0(n8582), .A1(n8583) );
  nand02 U5142 ( .Y(s_fraco1812_7_), .A0(n8590), .A1(n8591) );
  nand03 U5143 ( .Y(s_fraco1812_6_), .A0(n8598), .A1(n8599), .A2(n8600) );
  nand03 U5144 ( .Y(s_fraco1812_5_), .A0(n5482), .A1(n5511), .A2(n8611) );
  nand02 U5145 ( .Y(s_fraco1812_4_), .A0(n8616), .A1(n8617) );
  nand02 U5146 ( .Y(s_fraco1812_3_), .A0(n8622), .A1(n8623) );
  nand02 U5147 ( .Y(s_fraco1812_2_), .A0(n8631), .A1(n8632) );
  ao221 U5148 ( .Y(s_fraco1812_26_), .A0(n8635), .A1(n8329), .B0(n8637), .B1(
        n8337), .C0(n8639) );
  inv01 U5149 ( .Y(n8639), .A(n8640) );
  nand02 U5150 ( .Y(s_fraco1812_25_), .A0(n8648), .A1(n8649) );
  nand02 U5151 ( .Y(s_fraco1812_24_), .A0(n8658), .A1(n8659) );
  nand02 U5152 ( .Y(s_fraco1812_23_), .A0(n8667), .A1(n8668) );
  ao22 U5153 ( .Y(n8594), .A0(n8630), .A1(n8653), .B0(n8672), .B1(n8321) );
  nand03 U5154 ( .Y(s_fraco1812_22_), .A0(n5484), .A1(n8675), .A2(n8676) );
  nand03 U5155 ( .Y(s_fraco1812_21_), .A0(n5486), .A1(n8679), .A2(n8680) );
  nand02 U5156 ( .Y(s_fraco1812_20_), .A0(n8686), .A1(n8687) );
  oai22 U5157 ( .Y(n8621), .A0(n8688), .A1(n8328), .B0(n8689), .B1(n8323) );
  nand02 U5158 ( .Y(s_fraco1812_1_), .A0(n8690), .A1(n8691) );
  nand02 U5159 ( .Y(s_fraco1812_19_), .A0(n8695), .A1(n8696) );
  ao22 U5160 ( .Y(n8624), .A0(n8595), .A1(n8697), .B0(n8597), .B1(n8698) );
  nand02 U5161 ( .Y(s_fraco1812_18_), .A0(n8699), .A1(n8700) );
  inv01 U5162 ( .Y(n8702), .A(n8601) );
  nand02 U5163 ( .Y(s_fraco1812_17_), .A0(n8706), .A1(n8707) );
  inv01 U5164 ( .Y(n8709), .A(n8578) );
  inv01 U5165 ( .Y(n8681), .A(n8579) );
  nand02 U5166 ( .Y(s_fraco1812_16_), .A0(n8710), .A1(n8711) );
  nor02 U5167 ( .Y(n8636), .A0(n8712), .A1(n5552) );
  inv01 U5168 ( .Y(n8712), .A(s_shl1_4_) );
  nand03 U5169 ( .Y(s_fraco1812_15_), .A0(n5478), .A1(n5502), .A2(n8715) );
  nand03 U5170 ( .Y(s_fraco1812_14_), .A0(n5500), .A1(n5687), .A2(n8716) );
  oai22 U5171 ( .Y(n8612), .A0(n8721), .A1(n8462), .B0(n8385), .B1(n8461) );
  and03 U5172 ( .Y(n8638), .A0(s_shl1_3_), .A1(s_shl1_2_), .A2(n8334) );
  nand03 U5173 ( .Y(s_fraco1812_12_), .A0(n5480), .A1(n5647), .A2(n8726) );
  mux21 U5174 ( .Y(n8727), .A0(n8664), .A1(n8171), .S0(s_shl1_2_) );
  nand03 U5175 ( .Y(s_fraco1812_11_), .A0(n5476), .A1(n5509), .A2(n8730) );
  and02 U5176 ( .Y(n8641), .A0(n8335), .A1(n8163) );
  and02 U5177 ( .Y(n8608), .A0(n8333), .A1(n5607) );
  nand02 U5178 ( .Y(s_fraco1812_10_), .A0(n8733), .A1(n8734) );
  nor02 U5179 ( .Y(n8575), .A0(n8172), .A1(n8328) );
  inv01 U5180 ( .Y(n8698), .A(n8328) );
  inv01 U5181 ( .Y(n8735), .A(n8704) );
  nand02 U5182 ( .Y(n8704), .A0(n8370), .A1(s_qutnt_i[26]) );
  inv01 U5183 ( .Y(n8635), .A(n8736) );
  and02 U5184 ( .Y(n8653), .A0(s_shl1_2_), .A1(n8619) );
  nand02 U5185 ( .Y(n8646), .A0(s_shl1_1_), .A1(n8738) );
  or02 U5186 ( .Y(n8645), .A0(n8738), .A1(s_shl1_1_) );
  nand02 U5187 ( .Y(s_fraco1812_0_), .A0(n8739), .A1(n8740) );
  inv01 U5188 ( .Y(n8392), .A(s_qutnt_i[26]) );
  inv01 U5189 ( .Y(n8722), .A(n8370) );
  inv01 U5190 ( .Y(n8742), .A(n8588) );
  nor02 U5191 ( .Y(n8647), .A0(s_shl1_1_), .A1(s_shl1_0_) );
  and02 U5192 ( .Y(n8602), .A0(n8336), .A1(n8321) );
  nor02 U5193 ( .Y(n8655), .A0(s_shl1_3_), .A1(s_shl1_2_) );
  nor02 U5194 ( .Y(n8573), .A0(n5552), .A1(s_shl1_4_) );
  nand04 U5195 ( .Y(n8713), .A0(n8369), .A1(n8030), .A2(n8882), .A3(n8746) );
  nor02 U5196 ( .Y(n8577), .A0(n8275), .A1(n8172) );
  nor02 U5197 ( .Y(n8580), .A0(n8323), .A1(n8172) );
  nand02 U5198 ( .Y(n8719), .A0(n8744), .A1(n8747) );
  nor02 U5199 ( .Y(n8745), .A0(n8328), .A1(s_shr1_4_) );
  nand02 U5200 ( .Y(n8684), .A0(n8606), .A1(n8717) );
  nor02 U5201 ( .Y(n8629), .A0(s_shr1_1_), .A1(s_shr1_0_) );
  ao22 U5202 ( .Y(s_expo33281_8_), .A0(n____return3316_8_), .A1(n8553), .B0(
        s_expo2[8]), .B1(n8382) );
  ao22 U5203 ( .Y(s_expo33281_7_), .A0(n3318_7_), .A1(n8553), .B0(s_expo2[7]), 
        .B1(n8382) );
  ao22 U5204 ( .Y(s_expo33281_6_), .A0(n____return3316_6_), .A1(n8553), .B0(
        s_expo2[6]), .B1(n8382) );
  ao22 U5205 ( .Y(s_expo33281_5_), .A0(n____return3316_5_), .A1(n8553), .B0(
        s_expo2[5]), .B1(n8382) );
  ao22 U5206 ( .Y(s_expo33281_4_), .A0(n____return3316_4_), .A1(n8553), .B0(
        s_expo2[4]), .B1(n8382) );
  ao22 U5207 ( .Y(s_expo33281_3_), .A0(n____return3316_3_), .A1(n8553), .B0(
        s_expo2[3]), .B1(n8382) );
  ao22 U5208 ( .Y(s_expo33281_2_), .A0(n____return3316_2_), .A1(n8553), .B0(
        s_expo2[2]), .B1(n8382) );
  ao22 U5209 ( .Y(s_expo33281_1_), .A0(n____return3316_1_), .A1(n8553), .B0(
        s_expo2[1]), .B1(n8382) );
  ao22 U5210 ( .Y(s_expo33281_0_), .A0(n____return3316_0_), .A1(n8553), .B0(
        s_expo2[0]), .B1(n8382) );
  mux21 U5211 ( .Y(n8748), .A0(n1238_8_), .A1(s_expo1[8]), .S0(n8325) );
  mux21 U5212 ( .Y(n8749), .A0(n____return1236_7_), .A1(s_expo1[7]), .S0(n8325) );
  mux21 U5213 ( .Y(n8750), .A0(n____return1236_6_), .A1(s_expo1[6]), .S0(
        s_fraco1_26_) );
  mux21 U5214 ( .Y(n8751), .A0(n____return1236_5_), .A1(s_expo1[5]), .S0(
        s_fraco1_26_) );
  mux21 U5215 ( .Y(n8752), .A0(n____return1236_4_), .A1(s_expo1[4]), .S0(
        s_fraco1_26_) );
  mux21 U5216 ( .Y(n8753), .A0(n____return1236_3_), .A1(s_expo1[3]), .S0(
        s_fraco1_26_) );
  mux21 U5217 ( .Y(n8754), .A0(n____return1236_2_), .A1(s_expo1[2]), .S0(n8325) );
  mux21 U5218 ( .Y(n8755), .A0(n____return1236_1_), .A1(s_expo1[1]), .S0(n8325) );
  mux21 U5219 ( .Y(n8756), .A0(n____return1236_0_), .A1(s_expo1[0]), .S0(n8325) );
  nand02 U5220 ( .Y(s_expo1480_0_), .A0(n8391), .A1(n8416) );
  inv01 U5221 ( .Y(n8391), .A(n8340) );
  ao21 U5222 ( .Y(n8393), .A0(n8762), .A1(n8763), .B0(n5153) );
  nor02 U5223 ( .Y(n8764), .A0(s_exp_10_i_8_), .A1(n8765) );
  inv01 U5224 ( .Y(n8765), .A(n8090) );
  and03 U5225 ( .Y(n8763), .A0(n7732), .A1(n8161), .A2(n8071) );
  ao21 U5226 ( .Y(n8760), .A0(s_exp_10_i_4_), .A1(n8767), .B0(n5156) );
  ao21 U5227 ( .Y(n8406), .A0(s_exp_10_i_1_), .A1(n8769), .B0(n5178) );
  inv01 U5228 ( .Y(n8411), .A(n8405) );
  aoi21 U5229 ( .Y(n8757), .A0(s_exp_10_i_7_), .A1(n8775), .B0(n8090) );
  nor02 U5230 ( .Y(n8766), .A0(n8775), .A1(s_exp_10_i_7_) );
  ao21 U5231 ( .Y(n8759), .A0(s_exp_10_i_5_), .A1(n8777), .B0(n5155) );
  ao21 U5232 ( .Y(n8758), .A0(s_exp_10_i_6_), .A1(n8779), .B0(n5154) );
  nor02 U5233 ( .Y(n8776), .A0(n8779), .A1(s_exp_10_i_6_) );
  inv01 U5234 ( .Y(n8779), .A(n8778) );
  nor02 U5235 ( .Y(n8778), .A0(n8777), .A1(s_exp_10_i_5_) );
  inv01 U5236 ( .Y(n8777), .A(n8768) );
  nor02 U5237 ( .Y(n8768), .A0(n8767), .A1(s_exp_10_i_4_) );
  inv01 U5238 ( .Y(n8767), .A(n8772) );
  nor02 U5239 ( .Y(n8772), .A0(n8771), .A1(s_exp_10_i_3_) );
  inv01 U5240 ( .Y(n8771), .A(n8774) );
  nor02 U5241 ( .Y(n8774), .A0(n8773), .A1(s_exp_10_i_2_) );
  inv01 U5242 ( .Y(n8773), .A(n8770) );
  nor02 U5243 ( .Y(n8770), .A0(n8769), .A1(s_exp_10_i_1_) );
  inv01 U5244 ( .Y(n8769), .A(n8780) );
  ao21 U5245 ( .Y(n8761), .A0(s_qutnt_i[26]), .A1(s_exp_10_i_0_), .B0(n5448)
         );
  nor02 U5246 ( .Y(n8780), .A0(s_qutnt_i[26]), .A1(s_exp_10_i_0_) );
  nor02 U5247 ( .Y(n8781), .A0(n8747), .A1(n5597) );
  inv01 U5248 ( .Y(n8747), .A(s_shr1_4_) );
  nand03 U5249 ( .Y(n8782), .A0(s_shr1_3_), .A1(s_shr1_2_), .A2(n8169) );
  nand02 U5250 ( .Y(n____return2878_3_), .A0(n8784), .A1(n8275) );
  nand02 U5251 ( .Y(n8703), .A0(s_shr1_3_), .A1(n8717) );
  mux21 U5252 ( .Y(n8784), .A0(s_shr1_3_), .A1(n8697), .S0(n8169) );
  inv01 U5253 ( .Y(n8697), .A(n8322) );
  nand02 U5254 ( .Y(n8682), .A0(s_shr1_2_), .A1(n8606) );
  nor02 U5255 ( .Y(n8783), .A0(n8376), .A1(n8382) );
  nand02 U5256 ( .Y(n8628), .A0(s_shr1_1_), .A1(s_shr1_0_) );
  nand02 U5257 ( .Y(n____return2878_1_), .A0(n5464), .A1(n8379) );
  or02 U5258 ( .Y(n8626), .A0(n8785), .A1(s_shr1_0_) );
  nand02 U5259 ( .Y(n8627), .A0(s_shr1_0_), .A1(n8785) );
  inv01 U5260 ( .Y(n8785), .A(s_shr1_1_) );
  nand02 U5261 ( .Y(n8540), .A0(n3243_24_), .A1(n8381) );
  inv01 U5262 ( .Y(n8544), .A(n8567) );
  mux21 U5263 ( .Y(n8567), .A0(n8786), .A1(n8787), .S0(s_rmode_i_1_) );
  nor02 U5264 ( .Y(n8787), .A0(n8539), .A1(n8788) );
  xor2 U5265 ( .Y(n8788), .A0(s_sign_i), .A1(s_rmode_i_0_) );
  nand04 U5266 ( .Y(n8789), .A0(n7794), .A1(n7926), .A2(n7932), .A3(n7956) );
  nand04 U5267 ( .Y(n8791), .A0(n8884), .A1(n8885), .A2(n8886), .A3(n8887) );
  nand04 U5268 ( .Y(n8792), .A0(n8888), .A1(n8889), .A2(n8890), .A3(n8891) );
  nand04 U5269 ( .Y(n8793), .A0(n8894), .A1(n8895), .A2(n8892), .A3(n8893) );
  nand04 U5270 ( .Y(n8794), .A0(n8896), .A1(n8897), .A2(n8898), .A3(n8899) );
  inv01 U5271 ( .Y(n8790), .A(n8883) );
  post_norm_div_DW01_inc_9_0 add_216_plus_plus ( .A(s_expo2), .SUM({
        n____return3316_8_, n3318_7_, n____return3316_6_, n____return3316_5_, 
        n____return3316_4_, n____return3316_3_, n____return3316_2_, 
        n____return3316_1_, n____return3316_0_}) );
  post_norm_div_DW01_cmp2_6_0 gt_194_gt_gt ( .A({1'b0, s_r_zeros_4_, 
        s_r_zeros_3_, s_r_zeros_2_, s_r_zeros_1_, s_r_zeros_0_}), .B({n5151, 
        n7770, n____return2878_3_, n7788, n____return2878_1_, n5619}), .LEQ(
        1'b0), .TC(1'b0), .LT_LE(n____return2916) );
  post_norm_div_DW01_inc_25_0 add_209_plus_plus ( .A({1'b0, n8325, 
        s_fraco1_25_, s_fraco1_24_, s_fraco1_23_, s_fraco1_22_, s_fraco1_21_, 
        s_fraco1_20_, s_fraco1_19_, s_fraco1_18_, s_fraco1_17_, s_fraco1_16_, 
        s_fraco1_15_, s_fraco1_14_, s_fraco1_13_, s_fraco1_12_, s_fraco1_11_, 
        s_fraco1_10_, s_fraco1_9_, s_fraco1_8_, s_fraco1_7_, s_fraco1_6_, 
        s_fraco1_5_, s_fraco1_4_, s_fraco1_3_}), .SUM({n3243_24_, 
        n____return3241_23_, n____return3241_22_, n____return3241_21_, 
        n____return3241_20_, n____return3241_19_, n____return3241_18_, 
        n____return3241_17_, n____return3241_16_, n____return3241_15_, 
        n____return3241_14_, n____return3241_13_, n____return3241_12_, 
        n____return3241_11_, n____return3241_10_, n____return3241_9_, 
        n____return3241_8_, n____return3241_7_, n____return3241_6_, 
        n____return3241_5_, n____return3241_4_, n____return3241_3_, 
        n____return3241_2_, n____return3241_1_, n____return3241_0_}) );
  post_norm_div_DW01_dec_9_0 sub_188_minus_minus ( .A(s_expo1), .SUM({n1238_8_, 
        n____return1236_7_, n____return1236_6_, n____return1236_5_, 
        n____return1236_4_, n____return1236_3_, n____return1236_2_, 
        n____return1236_1_, n____return1236_0_}) );
endmodule


module pre_norm_sqrt_DW01_sub_9_0 ( A, B, CI, DIFF, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] DIFF;
  input CI;
  output CO;
  wire   carry_8_, carry_7_, carry_5_, carry_4_, carry_3_, carry_2_, B_not_4_,
         B_not_3_, B_not_2_, B_not_1_, B_not_0_, n5, n7, n9, n10, n11, n13,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50;

  xor2 U6 ( .Y(n5), .A0(A[6]), .A1(n18) );
  inv01 U7 ( .Y(DIFF[6]), .A(n5) );
  xor2 U8 ( .Y(n7), .A0(A[8]), .A1(n10) );
  inv01 U9 ( .Y(DIFF[8]), .A(n7) );
  inv01 U10 ( .Y(n9), .A(carry_8_) );
  inv01 U11 ( .Y(n10), .A(n9) );
  xor2 U12 ( .Y(n11), .A0(A[7]), .A1(n20) );
  inv01 U13 ( .Y(DIFF[7]), .A(n11) );
  xor2 U14 ( .Y(n13), .A0(A[5]), .A1(n50) );
  inv01 U15 ( .Y(DIFF[5]), .A(n13) );
  nor02 U16 ( .Y(n15), .A0(B_not_0_), .A1(A[0]) );
  inv02 U17 ( .Y(n16), .A(n15) );
  nor02 U18 ( .Y(n17), .A0(A[5]), .A1(n50) );
  inv01 U19 ( .Y(n18), .A(n17) );
  inv01 U20 ( .Y(n19), .A(n17) );
  buf02 U21 ( .Y(n20), .A(carry_7_) );
  buf02 U22 ( .Y(n21), .A(carry_7_) );
  buf02 U23 ( .Y(n22), .A(carry_4_) );
  inv01 U24 ( .Y(DIFF[2]), .A(n23) );
  inv02 U25 ( .Y(carry_3_), .A(n24) );
  inv02 U26 ( .Y(n25), .A(B_not_2_) );
  inv02 U27 ( .Y(n26), .A(A[2]) );
  inv02 U28 ( .Y(n27), .A(n49) );
  nor02 U29 ( .Y(n28), .A0(n25), .A1(n29) );
  nor02 U30 ( .Y(n30), .A0(n26), .A1(n31) );
  nor02 U31 ( .Y(n32), .A0(n27), .A1(n33) );
  nor02 U32 ( .Y(n34), .A0(n27), .A1(n35) );
  nor02 U33 ( .Y(n23), .A0(n36), .A1(n37) );
  nor02 U34 ( .Y(n38), .A0(n26), .A1(n27) );
  nor02 U35 ( .Y(n39), .A0(n25), .A1(n27) );
  nor02 U36 ( .Y(n40), .A0(n25), .A1(n26) );
  nor02 U37 ( .Y(n24), .A0(n40), .A1(n41) );
  nor02 U38 ( .Y(n42), .A0(A[2]), .A1(n49) );
  inv01 U39 ( .Y(n29), .A(n42) );
  nor02 U40 ( .Y(n43), .A0(B_not_2_), .A1(n49) );
  inv01 U41 ( .Y(n31), .A(n43) );
  nor02 U42 ( .Y(n44), .A0(B_not_2_), .A1(A[2]) );
  inv01 U43 ( .Y(n33), .A(n44) );
  nor02 U44 ( .Y(n45), .A0(n25), .A1(n26) );
  inv01 U45 ( .Y(n35), .A(n45) );
  nor02 U46 ( .Y(n46), .A0(n28), .A1(n30) );
  inv01 U47 ( .Y(n36), .A(n46) );
  nor02 U48 ( .Y(n47), .A0(n32), .A1(n34) );
  inv01 U49 ( .Y(n37), .A(n47) );
  nor02 U50 ( .Y(n48), .A0(n38), .A1(n39) );
  inv01 U51 ( .Y(n41), .A(n48) );
  buf02 U52 ( .Y(n49), .A(carry_2_) );
  buf02 U53 ( .Y(n50), .A(carry_5_) );
  inv01 U54 ( .Y(B_not_0_), .A(B[0]) );
  inv02 U55 ( .Y(B_not_1_), .A(B[1]) );
  inv02 U56 ( .Y(B_not_2_), .A(B[2]) );
  inv02 U57 ( .Y(B_not_3_), .A(B[3]) );
  inv02 U58 ( .Y(B_not_4_), .A(B[4]) );
  or02 U59 ( .Y(carry_8_), .A0(A[7]), .A1(n21) );
  or02 U60 ( .Y(carry_7_), .A0(A[6]), .A1(n19) );
  fadd1 U2_1 ( .S(DIFF[1]), .CO(carry_2_), .A(A[1]), .B(B_not_1_), .CI(n16) );
  fadd1 U2_3 ( .S(DIFF[3]), .CO(carry_4_), .A(A[3]), .B(B_not_3_), .CI(
        carry_3_) );
  fadd1 U2_4 ( .S(DIFF[4]), .CO(carry_5_), .A(A[4]), .B(B_not_4_), .CI(n22) );
endmodule


module pre_norm_sqrt ( clk_i, opa_i, fracta_52_o, exp_o );
  input [31:0] opa_i;
  output [51:0] fracta_52_o;
  output [7:0] exp_o;
  input clk_i;
  wire   n3996, n3997, s_exp_tem_8_, s_exp_tem_7_, s_exp_tem_6_, s_exp_tem_5_,
         s_exp_tem_4_, s_exp_tem_3_, s_exp_tem_2_, s_exp_tem_1_,
         s_sqr_zeros_o_4_, s_sqr_zeros_o_3_, s_sqr_zeros_o_2_,
         s_sqr_zeros_o_1_, s_sqr_zeros_o_0_, n1468_4_, n____return1466_8_,
         n____return1466_6_, n____return1466_5_, n____return1466_3_,
         n____return1466_2_, n____return1466_1_, n____return1466_0_,
         s_exp_o1553_7_, s_exp_o1553_6_, s_exp_o1553_5_, s_exp_o1553_4_,
         s_exp_o1553_3_, s_exp_o1553_2_, s_exp_o1553_1_, s_exp_o1553_0_, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, SYNOPSYS_UNCONNECTED_1;
  assign fracta_52_o[0] = 1'b0;
  assign fracta_52_o[1] = 1'b0;
  assign fracta_52_o[2] = 1'b0;
  assign fracta_52_o[3] = 1'b0;
  assign fracta_52_o[4] = 1'b0;
  assign fracta_52_o[5] = 1'b0;
  assign fracta_52_o[6] = 1'b0;
  assign fracta_52_o[7] = 1'b0;
  assign fracta_52_o[8] = 1'b0;
  assign fracta_52_o[9] = 1'b0;
  assign fracta_52_o[10] = 1'b0;
  assign fracta_52_o[11] = 1'b0;
  assign fracta_52_o[12] = 1'b0;
  assign fracta_52_o[13] = 1'b0;
  assign fracta_52_o[14] = 1'b0;
  assign fracta_52_o[15] = 1'b0;
  assign fracta_52_o[16] = 1'b0;
  assign fracta_52_o[17] = 1'b0;
  assign fracta_52_o[18] = 1'b0;
  assign fracta_52_o[19] = 1'b0;
  assign fracta_52_o[20] = 1'b0;
  assign fracta_52_o[21] = 1'b0;
  assign fracta_52_o[22] = 1'b0;
  assign fracta_52_o[23] = 1'b0;
  assign fracta_52_o[24] = 1'b0;
  assign fracta_52_o[25] = 1'b0;
  assign fracta_52_o[26] = 1'b0;

  dff s_exp_o_reg_7_ ( .Q(exp_o[7]), .D(s_exp_o1553_7_), .CLK(clk_i) );
  dff s_exp_o_reg_6_ ( .Q(exp_o[6]), .D(s_exp_o1553_6_), .CLK(clk_i) );
  dff s_exp_o_reg_5_ ( .Q(exp_o[5]), .D(s_exp_o1553_5_), .CLK(clk_i) );
  dff s_exp_o_reg_4_ ( .Q(exp_o[4]), .D(s_exp_o1553_4_), .CLK(clk_i) );
  dff s_exp_o_reg_3_ ( .Q(exp_o[3]), .D(s_exp_o1553_3_), .CLK(clk_i) );
  dff s_exp_o_reg_2_ ( .Q(exp_o[2]), .D(s_exp_o1553_2_), .CLK(clk_i) );
  dff s_exp_o_reg_1_ ( .Q(exp_o[1]), .D(s_exp_o1553_1_), .CLK(clk_i) );
  dff s_exp_o_reg_0_ ( .Q(exp_o[0]), .D(s_exp_o1553_0_), .CLK(clk_i) );
  inv04 U686 ( .Y(n3798), .A(n3796) );
  nand02 U687 ( .Y(n3850), .A0(n2527), .A1(n2528) );
  inv02 U688 ( .Y(n2529), .A(opa_i[18]) );
  inv02 U689 ( .Y(n2530), .A(opa_i[17]) );
  inv02 U690 ( .Y(n2531), .A(n3799) );
  inv02 U691 ( .Y(n2532), .A(opa_i[19]) );
  inv02 U692 ( .Y(n2533), .A(n3824) );
  inv02 U693 ( .Y(n2534), .A(n3825) );
  nand02 U694 ( .Y(n2535), .A0(n2531), .A1(n2536) );
  nand02 U695 ( .Y(n2537), .A0(n2532), .A1(n2538) );
  nand02 U696 ( .Y(n2539), .A0(n2533), .A1(n2540) );
  nand02 U697 ( .Y(n2541), .A0(n2533), .A1(n2542) );
  nand02 U698 ( .Y(n2543), .A0(n2534), .A1(n2544) );
  nand02 U699 ( .Y(n2545), .A0(n2534), .A1(n2546) );
  nand02 U700 ( .Y(n2547), .A0(n2534), .A1(n2548) );
  nand02 U701 ( .Y(n2549), .A0(n2534), .A1(n2550) );
  nand02 U702 ( .Y(n2551), .A0(n2529), .A1(n2530) );
  inv01 U703 ( .Y(n2536), .A(n2551) );
  nand02 U704 ( .Y(n2552), .A0(n2529), .A1(n2530) );
  inv01 U705 ( .Y(n2538), .A(n2552) );
  nand02 U706 ( .Y(n2553), .A0(n2529), .A1(n2531) );
  inv01 U707 ( .Y(n2540), .A(n2553) );
  nand02 U708 ( .Y(n2554), .A0(n2529), .A1(n2532) );
  inv01 U709 ( .Y(n2542), .A(n2554) );
  nand02 U710 ( .Y(n2555), .A0(n2530), .A1(n2531) );
  inv01 U711 ( .Y(n2544), .A(n2555) );
  nand02 U712 ( .Y(n2556), .A0(n2530), .A1(n2532) );
  inv01 U713 ( .Y(n2546), .A(n2556) );
  nand02 U714 ( .Y(n2557), .A0(n2531), .A1(n2533) );
  inv01 U715 ( .Y(n2548), .A(n2557) );
  nand02 U716 ( .Y(n2558), .A0(n2532), .A1(n2533) );
  inv01 U717 ( .Y(n2550), .A(n2558) );
  nand02 U718 ( .Y(n2559), .A0(n2535), .A1(n2537) );
  inv01 U719 ( .Y(n2560), .A(n2559) );
  nand02 U720 ( .Y(n2561), .A0(n2539), .A1(n2541) );
  inv01 U721 ( .Y(n2562), .A(n2561) );
  nand02 U722 ( .Y(n2563), .A0(n2560), .A1(n2562) );
  inv01 U723 ( .Y(n2527), .A(n2563) );
  nand02 U724 ( .Y(n2564), .A0(n2543), .A1(n2545) );
  inv01 U725 ( .Y(n2565), .A(n2564) );
  nand02 U726 ( .Y(n2566), .A0(n2547), .A1(n2549) );
  inv01 U727 ( .Y(n2567), .A(n2566) );
  nand02 U728 ( .Y(n2568), .A0(n2565), .A1(n2567) );
  inv01 U729 ( .Y(n2528), .A(n2568) );
  inv04 U730 ( .Y(n3825), .A(n3798) );
  nand02 U731 ( .Y(n3872), .A0(n2569), .A1(n2570) );
  inv02 U732 ( .Y(n2571), .A(n3800) );
  inv02 U733 ( .Y(n2572), .A(n3825) );
  inv02 U734 ( .Y(n2573), .A(n3799) );
  inv02 U735 ( .Y(n2574), .A(opa_i[1]) );
  inv02 U736 ( .Y(n2575), .A(opa_i[0]) );
  inv02 U737 ( .Y(n2576), .A(opa_i[2]) );
  nand02 U738 ( .Y(n2577), .A0(n2573), .A1(n2578) );
  nand02 U739 ( .Y(n2579), .A0(n2574), .A1(n2580) );
  nand02 U740 ( .Y(n2581), .A0(n2575), .A1(n2582) );
  nand02 U741 ( .Y(n2583), .A0(n2575), .A1(n2584) );
  nand02 U742 ( .Y(n2585), .A0(n2576), .A1(n2586) );
  nand02 U743 ( .Y(n2587), .A0(n2576), .A1(n2588) );
  nand02 U744 ( .Y(n2589), .A0(n2576), .A1(n2590) );
  nand02 U745 ( .Y(n2591), .A0(n2576), .A1(n2592) );
  nand02 U746 ( .Y(n2593), .A0(n2571), .A1(n2572) );
  inv01 U747 ( .Y(n2578), .A(n2593) );
  nand02 U748 ( .Y(n2594), .A0(n2571), .A1(n2572) );
  inv01 U749 ( .Y(n2580), .A(n2594) );
  nand02 U750 ( .Y(n2595), .A0(n2571), .A1(n2573) );
  inv01 U751 ( .Y(n2582), .A(n2595) );
  nand02 U752 ( .Y(n2596), .A0(n2571), .A1(n2574) );
  inv01 U753 ( .Y(n2584), .A(n2596) );
  nand02 U754 ( .Y(n2597), .A0(n2572), .A1(n2573) );
  inv01 U755 ( .Y(n2586), .A(n2597) );
  nand02 U756 ( .Y(n2598), .A0(n2572), .A1(n2574) );
  inv01 U757 ( .Y(n2588), .A(n2598) );
  nand02 U758 ( .Y(n2599), .A0(n2573), .A1(n2575) );
  inv01 U759 ( .Y(n2590), .A(n2599) );
  nand02 U760 ( .Y(n2600), .A0(n2574), .A1(n2575) );
  inv01 U761 ( .Y(n2592), .A(n2600) );
  nand02 U762 ( .Y(n2601), .A0(n2577), .A1(n2579) );
  inv01 U763 ( .Y(n2602), .A(n2601) );
  nand02 U764 ( .Y(n2603), .A0(n2581), .A1(n2583) );
  inv01 U765 ( .Y(n2604), .A(n2603) );
  nand02 U766 ( .Y(n2605), .A0(n2602), .A1(n2604) );
  inv01 U767 ( .Y(n2569), .A(n2605) );
  nand02 U768 ( .Y(n2606), .A0(n2585), .A1(n2587) );
  inv01 U769 ( .Y(n2607), .A(n2606) );
  nand02 U770 ( .Y(n2608), .A0(n2589), .A1(n2591) );
  inv01 U771 ( .Y(n2609), .A(n2608) );
  nand02 U772 ( .Y(n2610), .A0(n2607), .A1(n2609) );
  inv01 U773 ( .Y(n2570), .A(n2610) );
  buf08 U774 ( .Y(n3800), .A(n3826) );
  nand02 U775 ( .Y(n3822), .A0(n2611), .A1(n2612) );
  inv02 U776 ( .Y(n2613), .A(opa_i[20]) );
  inv02 U777 ( .Y(n2614), .A(n3824) );
  inv02 U778 ( .Y(n2615), .A(n3799) );
  inv02 U779 ( .Y(n2616), .A(opa_i[21]) );
  inv02 U780 ( .Y(n2617), .A(opa_i[19]) );
  inv02 U781 ( .Y(n2618), .A(n3825) );
  nand02 U782 ( .Y(n2619), .A0(n2615), .A1(n2620) );
  nand02 U783 ( .Y(n2621), .A0(n2616), .A1(n2622) );
  nand02 U784 ( .Y(n2623), .A0(n2617), .A1(n2624) );
  nand02 U785 ( .Y(n2625), .A0(n2617), .A1(n2626) );
  nand02 U786 ( .Y(n2627), .A0(n2618), .A1(n2628) );
  nand02 U787 ( .Y(n2629), .A0(n2618), .A1(n2630) );
  nand02 U788 ( .Y(n2631), .A0(n2618), .A1(n2632) );
  nand02 U789 ( .Y(n2633), .A0(n2618), .A1(n2634) );
  nand02 U790 ( .Y(n2635), .A0(n2613), .A1(n2614) );
  inv01 U791 ( .Y(n2620), .A(n2635) );
  nand02 U792 ( .Y(n2636), .A0(n2613), .A1(n2614) );
  inv01 U793 ( .Y(n2622), .A(n2636) );
  nand02 U794 ( .Y(n2637), .A0(n2613), .A1(n2615) );
  inv01 U795 ( .Y(n2624), .A(n2637) );
  nand02 U796 ( .Y(n2638), .A0(n2613), .A1(n2616) );
  inv01 U797 ( .Y(n2626), .A(n2638) );
  nand02 U798 ( .Y(n2639), .A0(n2614), .A1(n2615) );
  inv01 U799 ( .Y(n2628), .A(n2639) );
  nand02 U800 ( .Y(n2640), .A0(n2614), .A1(n2616) );
  inv01 U801 ( .Y(n2630), .A(n2640) );
  nand02 U802 ( .Y(n2641), .A0(n2615), .A1(n2617) );
  inv01 U803 ( .Y(n2632), .A(n2641) );
  nand02 U804 ( .Y(n2642), .A0(n2616), .A1(n2617) );
  inv01 U805 ( .Y(n2634), .A(n2642) );
  nand02 U806 ( .Y(n2643), .A0(n2619), .A1(n2621) );
  inv01 U807 ( .Y(n2644), .A(n2643) );
  nand02 U808 ( .Y(n2645), .A0(n2623), .A1(n2625) );
  inv01 U809 ( .Y(n2646), .A(n2645) );
  nand02 U810 ( .Y(n2647), .A0(n2644), .A1(n2646) );
  inv01 U811 ( .Y(n2611), .A(n2647) );
  nand02 U812 ( .Y(n2648), .A0(n2627), .A1(n2629) );
  inv01 U813 ( .Y(n2649), .A(n2648) );
  nand02 U814 ( .Y(n2650), .A0(n2631), .A1(n2633) );
  inv01 U815 ( .Y(n2651), .A(n2650) );
  nand02 U816 ( .Y(n2652), .A0(n2649), .A1(n2651) );
  inv01 U817 ( .Y(n2612), .A(n2652) );
  nand02 U818 ( .Y(n3839), .A0(n2653), .A1(n2654) );
  inv02 U819 ( .Y(n2655), .A(n3825) );
  inv02 U820 ( .Y(n2656), .A(opa_i[18]) );
  inv02 U821 ( .Y(n2657), .A(opa_i[20]) );
  inv02 U822 ( .Y(n2658), .A(n3799) );
  inv02 U823 ( .Y(n2659), .A(n3824) );
  inv02 U824 ( .Y(n2660), .A(opa_i[19]) );
  nand02 U825 ( .Y(n2661), .A0(n2657), .A1(n2662) );
  nand02 U826 ( .Y(n2663), .A0(n2658), .A1(n2664) );
  nand02 U827 ( .Y(n2665), .A0(n2659), .A1(n2666) );
  nand02 U828 ( .Y(n2667), .A0(n2659), .A1(n2668) );
  nand02 U829 ( .Y(n2669), .A0(n2660), .A1(n2670) );
  nand02 U830 ( .Y(n2671), .A0(n2660), .A1(n2672) );
  nand02 U831 ( .Y(n2673), .A0(n2660), .A1(n2674) );
  nand02 U832 ( .Y(n2675), .A0(n2660), .A1(n2676) );
  nand02 U833 ( .Y(n2677), .A0(n2655), .A1(n2656) );
  inv01 U834 ( .Y(n2662), .A(n2677) );
  nand02 U835 ( .Y(n2678), .A0(n2655), .A1(n2656) );
  inv01 U836 ( .Y(n2664), .A(n2678) );
  nand02 U837 ( .Y(n2679), .A0(n2655), .A1(n2657) );
  inv01 U838 ( .Y(n2666), .A(n2679) );
  nand02 U839 ( .Y(n2680), .A0(n2655), .A1(n2658) );
  inv01 U840 ( .Y(n2668), .A(n2680) );
  nand02 U841 ( .Y(n2681), .A0(n2656), .A1(n2657) );
  inv01 U842 ( .Y(n2670), .A(n2681) );
  nand02 U843 ( .Y(n2682), .A0(n2656), .A1(n2658) );
  inv01 U844 ( .Y(n2672), .A(n2682) );
  nand02 U845 ( .Y(n2683), .A0(n2657), .A1(n2659) );
  inv01 U846 ( .Y(n2674), .A(n2683) );
  nand02 U847 ( .Y(n2684), .A0(n2658), .A1(n2659) );
  inv01 U848 ( .Y(n2676), .A(n2684) );
  nand02 U849 ( .Y(n2685), .A0(n2661), .A1(n2663) );
  inv01 U850 ( .Y(n2686), .A(n2685) );
  nand02 U851 ( .Y(n2687), .A0(n2665), .A1(n2667) );
  inv01 U852 ( .Y(n2688), .A(n2687) );
  nand02 U853 ( .Y(n2689), .A0(n2686), .A1(n2688) );
  inv01 U854 ( .Y(n2653), .A(n2689) );
  nand02 U855 ( .Y(n2690), .A0(n2669), .A1(n2671) );
  inv01 U856 ( .Y(n2691), .A(n2690) );
  nand02 U857 ( .Y(n2692), .A0(n2673), .A1(n2675) );
  inv01 U858 ( .Y(n2693), .A(n2692) );
  nand02 U859 ( .Y(n2694), .A0(n2691), .A1(n2693) );
  inv01 U860 ( .Y(n2654), .A(n2694) );
  buf08 U861 ( .Y(n3799), .A(n3823) );
  nand02 U862 ( .Y(n3997), .A0(n2695), .A1(n2696) );
  inv01 U863 ( .Y(n2697), .A(n3857) );
  inv01 U864 ( .Y(n2698), .A(n3801) );
  inv01 U865 ( .Y(n2699), .A(n3805) );
  inv01 U866 ( .Y(n2700), .A(n3869) );
  nand02 U867 ( .Y(n2695), .A0(n2697), .A1(n2698) );
  nand02 U868 ( .Y(n2696), .A0(n2699), .A1(n2700) );
  inv01 U869 ( .Y(n3996), .A(n2701) );
  nor02 U870 ( .Y(n2702), .A0(n3801), .A1(n3847) );
  nor02 U871 ( .Y(n2703), .A0(n3857), .A1(n3805) );
  nor02 U872 ( .Y(n2701), .A0(n2702), .A1(n2703) );
  inv02 U873 ( .Y(n3787), .A(n3888) );
  inv02 U874 ( .Y(n3791), .A(n3887) );
  inv02 U875 ( .Y(n2858), .A(opa_i[11]) );
  inv02 U876 ( .Y(n3638), .A(opa_i[16]) );
  inv02 U877 ( .Y(n3358), .A(n3357) );
  inv04 U878 ( .Y(n3984), .A(opa_i[14]) );
  or02 U879 ( .Y(n2704), .A0(n3801), .A1(n3613) );
  inv01 U880 ( .Y(fracta_52_o[27]), .A(n2704) );
  buf02 U881 ( .Y(n2706), .A(s_sqr_zeros_o_2_) );
  inv02 U882 ( .Y(n3601), .A(opa_i[18]) );
  inv02 U883 ( .Y(n2768), .A(opa_i[13]) );
  inv02 U884 ( .Y(n2847), .A(opa_i[13]) );
  buf02 U885 ( .Y(n2707), .A(opa_i[6]) );
  inv02 U886 ( .Y(n2708), .A(n2707) );
  inv01 U887 ( .Y(n3759), .A(n2709) );
  inv01 U888 ( .Y(n2710), .A(n3799) );
  inv01 U889 ( .Y(n2711), .A(opa_i[0]) );
  inv01 U890 ( .Y(n2712), .A(n3800) );
  inv01 U891 ( .Y(n2713), .A(opa_i[1]) );
  nor02 U892 ( .Y(n2714), .A0(n2710), .A1(n2711) );
  nor02 U893 ( .Y(n2715), .A0(n2712), .A1(n2713) );
  nor02 U894 ( .Y(n2709), .A0(n2714), .A1(n2715) );
  or02 U895 ( .Y(n2716), .A0(n3972), .A1(n3961) );
  inv01 U896 ( .Y(n2717), .A(n2716) );
  inv08 U897 ( .Y(n3769), .A(n3768) );
  inv02 U898 ( .Y(n3419), .A(opa_i[15]) );
  inv02 U899 ( .Y(n3658), .A(opa_i[15]) );
  ao22 U900 ( .Y(n2718), .A0(n3827), .A1(n3794), .B0(n3828), .B1(n3806) );
  inv01 U901 ( .Y(n2719), .A(n2718) );
  nand02 U902 ( .Y(n3848), .A0(n2720), .A1(n2721) );
  inv01 U903 ( .Y(n2722), .A(n3806) );
  inv01 U904 ( .Y(n2723), .A(n3794) );
  inv01 U905 ( .Y(n2724), .A(n3851) );
  inv01 U906 ( .Y(n2725), .A(n3852) );
  nand02 U907 ( .Y(n2726), .A0(n2722), .A1(n2723) );
  nand02 U908 ( .Y(n2727), .A0(n2722), .A1(n2724) );
  nand02 U909 ( .Y(n2728), .A0(n2723), .A1(n2725) );
  nand02 U910 ( .Y(n2729), .A0(n2724), .A1(n2725) );
  nand02 U911 ( .Y(n2730), .A0(n2726), .A1(n2727) );
  inv01 U912 ( .Y(n2720), .A(n2730) );
  nand02 U913 ( .Y(n2731), .A0(n2728), .A1(n2729) );
  inv01 U914 ( .Y(n2721), .A(n2731) );
  ao22 U915 ( .Y(n2732), .A0(n3840), .A1(n3794), .B0(n3841), .B1(n3806) );
  inv01 U916 ( .Y(n2733), .A(n2732) );
  nand02 U917 ( .Y(n3988), .A0(n2734), .A1(n2735) );
  inv01 U918 ( .Y(n2736), .A(opa_i[22]) );
  inv01 U919 ( .Y(n2737), .A(n3989) );
  inv01 U920 ( .Y(n2738), .A(opa_i[20]) );
  nand02 U921 ( .Y(n2734), .A0(n2736), .A1(n2737) );
  nand02 U922 ( .Y(n2735), .A0(n2736), .A1(n2738) );
  ao21 U923 ( .Y(n2739), .A0(n3960), .A1(n3961), .B0(n3938) );
  inv01 U924 ( .Y(n2740), .A(n2739) );
  nand02 U925 ( .Y(n2741), .A0(n3978), .A1(n2768) );
  inv02 U926 ( .Y(n2742), .A(n2741) );
  inv02 U927 ( .Y(n3302), .A(opa_i[19]) );
  nand02 U928 ( .Y(n3922), .A0(n2743), .A1(n2744) );
  inv01 U929 ( .Y(n2745), .A(opa_i[3]) );
  inv01 U930 ( .Y(n2746), .A(n3799) );
  inv01 U931 ( .Y(n2747), .A(n3800) );
  nand02 U932 ( .Y(n2748), .A0(n2745), .A1(n3309) );
  nand02 U933 ( .Y(n2749), .A0(n2745), .A1(n2746) );
  nand02 U934 ( .Y(n2750), .A0(n3309), .A1(n2747) );
  nand02 U935 ( .Y(n2751), .A0(n2746), .A1(n2747) );
  nand02 U936 ( .Y(n2752), .A0(n2748), .A1(n2749) );
  inv01 U937 ( .Y(n2743), .A(n2752) );
  nand02 U938 ( .Y(n2753), .A0(n2750), .A1(n2751) );
  inv01 U939 ( .Y(n2744), .A(n2753) );
  nand02 U940 ( .Y(n3912), .A0(n2754), .A1(n2755) );
  inv01 U941 ( .Y(n2756), .A(opa_i[8]) );
  inv01 U942 ( .Y(n2757), .A(opa_i[7]) );
  inv01 U943 ( .Y(n2758), .A(n3799) );
  inv01 U944 ( .Y(n2759), .A(n3800) );
  nand02 U945 ( .Y(n2760), .A0(n2756), .A1(n2757) );
  nand02 U946 ( .Y(n2761), .A0(n2756), .A1(n2758) );
  nand02 U947 ( .Y(n2762), .A0(n2757), .A1(n2759) );
  nand02 U948 ( .Y(n2763), .A0(n2758), .A1(n2759) );
  nand02 U949 ( .Y(n2764), .A0(n2760), .A1(n2761) );
  inv01 U950 ( .Y(n2754), .A(n2764) );
  nand02 U951 ( .Y(n2765), .A0(n2762), .A1(n2763) );
  inv01 U952 ( .Y(n2755), .A(n2765) );
  nand02 U953 ( .Y(n3898), .A0(n2766), .A1(n2767) );
  inv01 U954 ( .Y(n2769), .A(opa_i[12]) );
  inv01 U955 ( .Y(n2770), .A(n3799) );
  inv01 U956 ( .Y(n2771), .A(n3800) );
  nand02 U957 ( .Y(n2772), .A0(n2768), .A1(n2769) );
  nand02 U958 ( .Y(n2773), .A0(n2768), .A1(n2770) );
  nand02 U959 ( .Y(n2774), .A0(n2769), .A1(n2771) );
  nand02 U960 ( .Y(n2775), .A0(n2770), .A1(n2771) );
  nand02 U961 ( .Y(n2776), .A0(n2772), .A1(n2773) );
  inv01 U962 ( .Y(n2766), .A(n2776) );
  nand02 U963 ( .Y(n2777), .A0(n2774), .A1(n2775) );
  inv01 U964 ( .Y(n2767), .A(n2777) );
  nand02 U965 ( .Y(n3903), .A0(n2778), .A1(n2779) );
  inv01 U966 ( .Y(n2780), .A(opa_i[12]) );
  inv01 U967 ( .Y(n2781), .A(n3799) );
  inv01 U968 ( .Y(n2782), .A(n3800) );
  nand02 U969 ( .Y(n2783), .A0(n2780), .A1(n2858) );
  nand02 U970 ( .Y(n2784), .A0(n2780), .A1(n2781) );
  nand02 U971 ( .Y(n2785), .A0(n2858), .A1(n2782) );
  nand02 U972 ( .Y(n2786), .A0(n2781), .A1(n2782) );
  nand02 U973 ( .Y(n2787), .A0(n2783), .A1(n2784) );
  inv01 U974 ( .Y(n2778), .A(n2787) );
  nand02 U975 ( .Y(n2788), .A0(n2785), .A1(n2786) );
  inv01 U976 ( .Y(n2779), .A(n2788) );
  inv02 U977 ( .Y(n2789), .A(n____return1466_8_) );
  inv08 U978 ( .Y(n2790), .A(n2789) );
  nand02 U979 ( .Y(n3917), .A0(n2791), .A1(n2792) );
  inv01 U980 ( .Y(n2793), .A(opa_i[5]) );
  inv01 U981 ( .Y(n2794), .A(n3799) );
  inv01 U982 ( .Y(n2795), .A(n3800) );
  nand02 U983 ( .Y(n2796), .A0(n2793), .A1(n3767) );
  nand02 U984 ( .Y(n2797), .A0(n2793), .A1(n2794) );
  nand02 U985 ( .Y(n2798), .A0(n3767), .A1(n2795) );
  nand02 U986 ( .Y(n2799), .A0(n2794), .A1(n2795) );
  nand02 U987 ( .Y(n2800), .A0(n2796), .A1(n2797) );
  inv01 U988 ( .Y(n2791), .A(n2800) );
  nand02 U989 ( .Y(n2801), .A0(n2798), .A1(n2799) );
  inv01 U990 ( .Y(n2792), .A(n2801) );
  nand02 U991 ( .Y(n3908), .A0(n2802), .A1(n2803) );
  inv01 U992 ( .Y(n2804), .A(opa_i[10]) );
  inv01 U993 ( .Y(n2805), .A(n3799) );
  inv01 U994 ( .Y(n2806), .A(n3800) );
  nand02 U995 ( .Y(n2807), .A0(n2804), .A1(n3902) );
  nand02 U996 ( .Y(n2808), .A0(n2804), .A1(n2805) );
  nand02 U997 ( .Y(n2809), .A0(n3902), .A1(n2806) );
  nand02 U998 ( .Y(n2810), .A0(n2805), .A1(n2806) );
  nand02 U999 ( .Y(n2811), .A0(n2807), .A1(n2808) );
  inv01 U1000 ( .Y(n2802), .A(n2811) );
  nand02 U1001 ( .Y(n2812), .A0(n2809), .A1(n2810) );
  inv01 U1002 ( .Y(n2803), .A(n2812) );
  nand02 U1003 ( .Y(n3910), .A0(n2813), .A1(n2814) );
  inv01 U1004 ( .Y(n2815), .A(opa_i[9]) );
  inv01 U1005 ( .Y(n2816), .A(n3799) );
  inv01 U1006 ( .Y(n2817), .A(n3800) );
  nand02 U1007 ( .Y(n2818), .A0(n2815), .A1(n3905) );
  nand02 U1008 ( .Y(n2819), .A0(n2815), .A1(n2816) );
  nand02 U1009 ( .Y(n2820), .A0(n3905), .A1(n2817) );
  nand02 U1010 ( .Y(n2821), .A0(n2816), .A1(n2817) );
  nand02 U1011 ( .Y(n2822), .A0(n2818), .A1(n2819) );
  inv01 U1012 ( .Y(n2813), .A(n2822) );
  nand02 U1013 ( .Y(n2823), .A0(n2820), .A1(n2821) );
  inv01 U1014 ( .Y(n2814), .A(n2823) );
  nand02 U1015 ( .Y(n3920), .A0(n2824), .A1(n2825) );
  inv01 U1016 ( .Y(n2826), .A(opa_i[4]) );
  inv01 U1017 ( .Y(n2827), .A(n3799) );
  inv01 U1018 ( .Y(n2828), .A(n3800) );
  nand02 U1019 ( .Y(n2829), .A0(n2826), .A1(n3915) );
  nand02 U1020 ( .Y(n2830), .A0(n2826), .A1(n2827) );
  nand02 U1021 ( .Y(n2831), .A0(n3915), .A1(n2828) );
  nand02 U1022 ( .Y(n2832), .A0(n2827), .A1(n2828) );
  nand02 U1023 ( .Y(n2833), .A0(n2829), .A1(n2830) );
  inv01 U1024 ( .Y(n2824), .A(n2833) );
  nand02 U1025 ( .Y(n2834), .A0(n2831), .A1(n2832) );
  inv01 U1026 ( .Y(n2825), .A(n2834) );
  nand02 U1027 ( .Y(n3916), .A0(n2835), .A1(n2836) );
  inv01 U1028 ( .Y(n2837), .A(n3799) );
  inv01 U1029 ( .Y(n2838), .A(n3800) );
  nand02 U1030 ( .Y(n2839), .A0(n2708), .A1(n3312) );
  nand02 U1031 ( .Y(n2840), .A0(n2708), .A1(n2837) );
  nand02 U1032 ( .Y(n2841), .A0(n3312), .A1(n2838) );
  nand02 U1033 ( .Y(n2842), .A0(n2837), .A1(n2838) );
  nand02 U1034 ( .Y(n2843), .A0(n2839), .A1(n2840) );
  inv01 U1035 ( .Y(n2835), .A(n2843) );
  nand02 U1036 ( .Y(n2844), .A0(n2841), .A1(n2842) );
  inv01 U1037 ( .Y(n2836), .A(n2844) );
  nand02 U1038 ( .Y(n3895), .A0(n2845), .A1(n2846) );
  inv01 U1039 ( .Y(n2848), .A(n3799) );
  inv01 U1040 ( .Y(n2849), .A(n3800) );
  nand02 U1041 ( .Y(n2850), .A0(n3984), .A1(n2847) );
  nand02 U1042 ( .Y(n2851), .A0(n3984), .A1(n2848) );
  nand02 U1043 ( .Y(n2852), .A0(n2847), .A1(n2849) );
  nand02 U1044 ( .Y(n2853), .A0(n2848), .A1(n2849) );
  nand02 U1045 ( .Y(n2854), .A0(n2850), .A1(n2851) );
  inv01 U1046 ( .Y(n2845), .A(n2854) );
  nand02 U1047 ( .Y(n2855), .A0(n2852), .A1(n2853) );
  inv01 U1048 ( .Y(n2846), .A(n2855) );
  nand02 U1049 ( .Y(n3906), .A0(n2856), .A1(n2857) );
  inv01 U1050 ( .Y(n2859), .A(n3799) );
  inv01 U1051 ( .Y(n2860), .A(n3800) );
  nand02 U1052 ( .Y(n2861), .A0(n2858), .A1(n3754) );
  nand02 U1053 ( .Y(n2862), .A0(n2858), .A1(n2859) );
  nand02 U1054 ( .Y(n2863), .A0(n3754), .A1(n2860) );
  nand02 U1055 ( .Y(n2864), .A0(n2859), .A1(n2860) );
  nand02 U1056 ( .Y(n2865), .A0(n2861), .A1(n2862) );
  inv01 U1057 ( .Y(n2856), .A(n2865) );
  nand02 U1058 ( .Y(n2866), .A0(n2863), .A1(n2864) );
  inv01 U1059 ( .Y(n2857), .A(n2866) );
  buf02 U1060 ( .Y(fracta_52_o[45]), .A(n3997) );
  buf02 U1061 ( .Y(fracta_52_o[46]), .A(n3996) );
  inv01 U1062 ( .Y(fracta_52_o[47]), .A(n2869) );
  nor02 U1063 ( .Y(n2870), .A0(n3801), .A1(n3837) );
  nor02 U1064 ( .Y(n2871), .A0(n3847), .A1(n3805) );
  nor02 U1065 ( .Y(n2869), .A0(n2870), .A1(n2871) );
  or03 U1066 ( .Y(n2872), .A0(n3946), .A1(n3932), .A2(n3933) );
  inv01 U1067 ( .Y(n2873), .A(n2872) );
  nand02 U1068 ( .Y(n3891), .A0(n2874), .A1(n2875) );
  inv01 U1069 ( .Y(n2876), .A(n3799) );
  inv01 U1070 ( .Y(n2877), .A(n3800) );
  nand02 U1071 ( .Y(n2878), .A0(n3658), .A1(n3984) );
  nand02 U1072 ( .Y(n2879), .A0(n3419), .A1(n2876) );
  nand02 U1073 ( .Y(n2880), .A0(n3984), .A1(n2877) );
  nand02 U1074 ( .Y(n2881), .A0(n2876), .A1(n2877) );
  nand02 U1075 ( .Y(n2882), .A0(n2878), .A1(n2879) );
  inv01 U1076 ( .Y(n2874), .A(n2882) );
  nand02 U1077 ( .Y(n2883), .A0(n2880), .A1(n2881) );
  inv01 U1078 ( .Y(n2875), .A(n2883) );
  nand02 U1079 ( .Y(n3914), .A0(n2884), .A1(n2885) );
  inv01 U1080 ( .Y(n2886), .A(opa_i[7]) );
  inv01 U1081 ( .Y(n2887), .A(n3799) );
  inv01 U1082 ( .Y(n2888), .A(n3800) );
  nand02 U1083 ( .Y(n2889), .A0(n2886), .A1(n2708) );
  nand02 U1084 ( .Y(n2890), .A0(n2886), .A1(n2887) );
  nand02 U1085 ( .Y(n2891), .A0(n2708), .A1(n2888) );
  nand02 U1086 ( .Y(n2892), .A0(n2887), .A1(n2888) );
  nand02 U1087 ( .Y(n2893), .A0(n2889), .A1(n2890) );
  inv01 U1088 ( .Y(n2884), .A(n2893) );
  nand02 U1089 ( .Y(n2894), .A0(n2891), .A1(n2892) );
  inv01 U1090 ( .Y(n2885), .A(n2894) );
  inv01 U1091 ( .Y(fracta_52_o[44]), .A(n2895) );
  nor02 U1092 ( .Y(n2896), .A0(n3801), .A1(n3869) );
  nor02 U1093 ( .Y(n2897), .A0(n3875), .A1(n3805) );
  nor02 U1094 ( .Y(n2895), .A0(n2896), .A1(n2897) );
  inv01 U1095 ( .Y(fracta_52_o[49]), .A(n2898) );
  nor02 U1096 ( .Y(n2899), .A0(n3801), .A1(n3820) );
  nor02 U1097 ( .Y(n2900), .A0(n3819), .A1(n3805) );
  nor02 U1098 ( .Y(n2898), .A0(n2899), .A1(n2900) );
  nand02 U1099 ( .Y(n3867), .A0(n2901), .A1(n2902) );
  inv01 U1100 ( .Y(n2903), .A(n3800) );
  inv01 U1101 ( .Y(n2904), .A(n3799) );
  nand02 U1102 ( .Y(n2905), .A0(n2903), .A1(n3601) );
  nand02 U1103 ( .Y(n2906), .A0(n2903), .A1(n2904) );
  nand02 U1104 ( .Y(n2907), .A0(n3601), .A1(n3302) );
  nand02 U1105 ( .Y(n2908), .A0(n2904), .A1(n3302) );
  nand02 U1106 ( .Y(n2909), .A0(n2905), .A1(n2906) );
  inv01 U1107 ( .Y(n2901), .A(n2909) );
  nand02 U1108 ( .Y(n2910), .A0(n2907), .A1(n2908) );
  inv01 U1109 ( .Y(n2902), .A(n2910) );
  nand02 U1110 ( .Y(fracta_52_o[29]), .A0(n2911), .A1(n2912) );
  inv01 U1111 ( .Y(n2913), .A(n3612) );
  inv01 U1112 ( .Y(n2914), .A(n3762) );
  inv01 U1113 ( .Y(n2915), .A(n3780) );
  inv01 U1114 ( .Y(n2916), .A(n3801) );
  nand02 U1115 ( .Y(n2911), .A0(n2913), .A1(n2914) );
  nand02 U1116 ( .Y(n2912), .A0(n2915), .A1(n2916) );
  inv01 U1117 ( .Y(fracta_52_o[31]), .A(n2917) );
  nor02 U1118 ( .Y(n2918), .A0(n3860), .A1(n3612) );
  nor02 U1119 ( .Y(n2919), .A0(n3801), .A1(n3772) );
  nor02 U1120 ( .Y(n2917), .A0(n2918), .A1(n2919) );
  or02 U1121 ( .Y(n2920), .A0(n3784), .A1(n3785) );
  inv02 U1122 ( .Y(n2921), .A(n2920) );
  inv01 U1123 ( .Y(fracta_52_o[35]), .A(n2922) );
  nor02 U1124 ( .Y(n2923), .A0(n3699), .A1(n3775) );
  nor02 U1125 ( .Y(n2924), .A0(n3801), .A1(n3909) );
  nor02 U1126 ( .Y(n2922), .A0(n2923), .A1(n2924) );
  nand02 U1127 ( .Y(fracta_52_o[34]), .A0(n2925), .A1(n2926) );
  inv01 U1128 ( .Y(n2927), .A(n3775) );
  inv01 U1129 ( .Y(n2928), .A(n3596) );
  inv01 U1130 ( .Y(n2929), .A(n3699) );
  inv01 U1131 ( .Y(n2930), .A(n3801) );
  nand02 U1132 ( .Y(n2925), .A0(n2927), .A1(n2928) );
  nand02 U1133 ( .Y(n2926), .A0(n2929), .A1(n2930) );
  nand02 U1134 ( .Y(fracta_52_o[33]), .A0(n2931), .A1(n2932) );
  inv01 U1135 ( .Y(n2933), .A(n3775) );
  inv01 U1136 ( .Y(n2934), .A(n3611) );
  inv01 U1137 ( .Y(n2935), .A(n3596) );
  inv01 U1138 ( .Y(n2936), .A(n3801) );
  nand02 U1139 ( .Y(n2931), .A0(n2933), .A1(n2934) );
  nand02 U1140 ( .Y(n2932), .A0(n2935), .A1(n2936) );
  nand02 U1141 ( .Y(fracta_52_o[28]), .A0(n2937), .A1(n2938) );
  inv01 U1142 ( .Y(n2939), .A(n3612) );
  inv01 U1143 ( .Y(n2940), .A(n3613) );
  inv01 U1144 ( .Y(n2941), .A(n3762) );
  inv01 U1145 ( .Y(n2942), .A(n3801) );
  nand02 U1146 ( .Y(n2937), .A0(n2939), .A1(n2940) );
  nand02 U1147 ( .Y(n2938), .A0(n2941), .A1(n2942) );
  inv01 U1148 ( .Y(fracta_52_o[30]), .A(n2943) );
  nor02 U1149 ( .Y(n2944), .A0(n3780), .A1(n3612) );
  nor02 U1150 ( .Y(n2945), .A0(n3801), .A1(n3860) );
  nor02 U1151 ( .Y(n2943), .A0(n2944), .A1(n2945) );
  buf02 U1152 ( .Y(n3612), .A(n3918) );
  inv01 U1153 ( .Y(fracta_52_o[48]), .A(n2946) );
  nor02 U1154 ( .Y(n2947), .A0(n3801), .A1(n3819) );
  nor02 U1155 ( .Y(n2948), .A0(n3837), .A1(n3805) );
  nor02 U1156 ( .Y(n2946), .A0(n2947), .A1(n2948) );
  inv04 U1157 ( .Y(n3805), .A(n3769) );
  inv08 U1158 ( .Y(n3801), .A(n3805) );
  inv02 U1159 ( .Y(n3938), .A(n2949) );
  nand02 U1160 ( .Y(n2949), .A0(opa_i[9]), .A1(n2950) );
  nand02 U1161 ( .Y(n2951), .A0(n3975), .A1(n3754) );
  inv01 U1162 ( .Y(n2950), .A(n2951) );
  inv01 U1163 ( .Y(n3880), .A(n2952) );
  nor02 U1164 ( .Y(n2953), .A0(n3855), .A1(n3789) );
  nor02 U1165 ( .Y(n2954), .A0(n3613), .A1(n3700) );
  nor02 U1166 ( .Y(n2955), .A0(n3794), .A1(n3881) );
  nor02 U1167 ( .Y(n2952), .A0(n2955), .A1(n2956) );
  nor02 U1168 ( .Y(n2957), .A0(n2953), .A1(n2954) );
  inv01 U1169 ( .Y(n2956), .A(n2957) );
  buf02 U1170 ( .Y(n3613), .A(n3882) );
  buf02 U1171 ( .Y(n3789), .A(n3863) );
  inv01 U1172 ( .Y(n3858), .A(n2958) );
  nor02 U1173 ( .Y(n2959), .A0(n3862), .A1(n3789) );
  nor02 U1174 ( .Y(n2960), .A0(n3860), .A1(n3700) );
  nor02 U1175 ( .Y(n2961), .A0(n3794), .A1(n3859) );
  nor02 U1176 ( .Y(n2958), .A0(n2961), .A1(n2962) );
  nor02 U1177 ( .Y(n2963), .A0(n2959), .A1(n2960) );
  inv01 U1178 ( .Y(n2962), .A(n2963) );
  inv02 U1179 ( .Y(n3847), .A(n3858) );
  inv04 U1180 ( .Y(n3794), .A(n3793) );
  inv01 U1181 ( .Y(n3876), .A(n2964) );
  nor02 U1182 ( .Y(n2965), .A0(n3843), .A1(n3789) );
  nor02 U1183 ( .Y(n2966), .A0(n3761), .A1(n3861) );
  nor02 U1184 ( .Y(n2967), .A0(n3794), .A1(n3877) );
  nor02 U1185 ( .Y(n2964), .A0(n2967), .A1(n2968) );
  nor02 U1186 ( .Y(n2969), .A0(n2965), .A1(n2966) );
  inv01 U1187 ( .Y(n2968), .A(n2969) );
  inv02 U1188 ( .Y(n3869), .A(n3876) );
  inv01 U1189 ( .Y(n3870), .A(n2970) );
  nor02 U1190 ( .Y(n2971), .A0(n3831), .A1(n3789) );
  nor02 U1191 ( .Y(n2972), .A0(n3780), .A1(n3700) );
  nor02 U1192 ( .Y(n2973), .A0(n3794), .A1(n3871) );
  nor02 U1193 ( .Y(n2970), .A0(n2973), .A1(n2974) );
  nor02 U1194 ( .Y(n2975), .A0(n2971), .A1(n2972) );
  inv01 U1195 ( .Y(n2974), .A(n2975) );
  inv02 U1196 ( .Y(n3857), .A(n3870) );
  inv01 U1197 ( .Y(n3977), .A(n2976) );
  inv01 U1198 ( .Y(n2977), .A(opa_i[0]) );
  inv01 U1199 ( .Y(n2978), .A(n3919) );
  inv01 U1200 ( .Y(n2979), .A(n3980) );
  nor02 U1201 ( .Y(n2976), .A0(n2979), .A1(n2980) );
  nor02 U1202 ( .Y(n2981), .A0(n2977), .A1(n2978) );
  inv01 U1203 ( .Y(n2980), .A(n2981) );
  inv01 U1204 ( .Y(n3852), .A(n2982) );
  nor02 U1205 ( .Y(n2983), .A0(n3855), .A1(n3779) );
  nor02 U1206 ( .Y(n2984), .A0(n3854), .A1(n3750) );
  nor02 U1207 ( .Y(n2985), .A0(n3853), .A1(n3749) );
  nor02 U1208 ( .Y(n2982), .A0(n2985), .A1(n2986) );
  nor02 U1209 ( .Y(n2987), .A0(n2983), .A1(n2984) );
  inv01 U1210 ( .Y(n2986), .A(n2987) );
  buf02 U1211 ( .Y(n3779), .A(n3832) );
  buf02 U1212 ( .Y(n2988), .A(n3991) );
  inv01 U1213 ( .Y(n3841), .A(n2989) );
  nor02 U1214 ( .Y(n2990), .A0(n3844), .A1(n3749) );
  nor02 U1215 ( .Y(n2991), .A0(n3843), .A1(n3779) );
  nor02 U1216 ( .Y(n2992), .A0(n3842), .A1(n3830) );
  nor02 U1217 ( .Y(n2989), .A0(n2992), .A1(n2993) );
  nor02 U1218 ( .Y(n2994), .A0(n2990), .A1(n2991) );
  inv01 U1219 ( .Y(n2993), .A(n2994) );
  inv01 U1220 ( .Y(n3828), .A(n2995) );
  nor02 U1221 ( .Y(n2996), .A0(n3833), .A1(n3749) );
  nor02 U1222 ( .Y(n2997), .A0(n3831), .A1(n3779) );
  nor02 U1223 ( .Y(n2998), .A0(n3829), .A1(n3751) );
  nor02 U1224 ( .Y(n2995), .A0(n2998), .A1(n2999) );
  nor02 U1225 ( .Y(n3000), .A0(n2996), .A1(n2997) );
  inv01 U1226 ( .Y(n2999), .A(n3000) );
  buf02 U1227 ( .Y(n3749), .A(n3834) );
  nand02 U1228 ( .Y(n3001), .A0(n3979), .A1(n3312) );
  inv02 U1229 ( .Y(n3002), .A(n3001) );
  nand02 U1230 ( .Y(fracta_52_o[39]), .A0(n3003), .A1(n3004) );
  inv01 U1231 ( .Y(n3005), .A(n3801) );
  inv01 U1232 ( .Y(n3006), .A(n3899) );
  inv01 U1233 ( .Y(n3007), .A(n3056) );
  nand02 U1234 ( .Y(n3008), .A0(n3769), .A1(n3005) );
  nand02 U1235 ( .Y(n3009), .A0(n3801), .A1(n3006) );
  nand02 U1236 ( .Y(n3010), .A0(n3005), .A1(n3007) );
  nand02 U1237 ( .Y(n3011), .A0(n3006), .A1(n3007) );
  nand02 U1238 ( .Y(n3012), .A0(n3008), .A1(n3009) );
  inv01 U1239 ( .Y(n3003), .A(n3012) );
  nand02 U1240 ( .Y(n3013), .A0(n3010), .A1(n3011) );
  inv01 U1241 ( .Y(n3004), .A(n3013) );
  inv02 U1242 ( .Y(n3014), .A(n____return1466_6_) );
  inv08 U1243 ( .Y(n3015), .A(n3014) );
  inv02 U1244 ( .Y(n____return1466_5_), .A(n3016) );
  inv01 U1245 ( .Y(n3017), .A(n3993) );
  inv01 U1246 ( .Y(n3018), .A(opa_i[28]) );
  nor02 U1247 ( .Y(n3019), .A0(n3017), .A1(n3018) );
  nor02 U1248 ( .Y(n3016), .A0(n3019), .A1(n3111) );
  nand02 U1249 ( .Y(fracta_52_o[36]), .A0(n3020), .A1(n3021) );
  inv01 U1250 ( .Y(n3022), .A(n3801) );
  inv01 U1251 ( .Y(n3023), .A(n3909) );
  inv01 U1252 ( .Y(n3024), .A(n3907) );
  nand02 U1253 ( .Y(n3025), .A0(n3769), .A1(n3022) );
  nand02 U1254 ( .Y(n3026), .A0(n3769), .A1(n3023) );
  nand02 U1255 ( .Y(n3027), .A0(n3022), .A1(n3024) );
  nand02 U1256 ( .Y(n3028), .A0(n3023), .A1(n3024) );
  nand02 U1257 ( .Y(n3029), .A0(n3025), .A1(n3026) );
  inv01 U1258 ( .Y(n3020), .A(n3029) );
  nand02 U1259 ( .Y(n3030), .A0(n3027), .A1(n3028) );
  inv01 U1260 ( .Y(n3021), .A(n3030) );
  nand02 U1261 ( .Y(fracta_52_o[40]), .A0(n3031), .A1(n3032) );
  inv01 U1262 ( .Y(n3033), .A(n3801) );
  inv01 U1263 ( .Y(n3034), .A(n3056) );
  inv01 U1264 ( .Y(n3035), .A(n3892) );
  nand02 U1265 ( .Y(n3036), .A0(n3769), .A1(n3033) );
  nand02 U1266 ( .Y(n3037), .A0(n3769), .A1(n3034) );
  nand02 U1267 ( .Y(n3038), .A0(n3033), .A1(n3035) );
  nand02 U1268 ( .Y(n3039), .A0(n3034), .A1(n3035) );
  nand02 U1269 ( .Y(n3040), .A0(n3036), .A1(n3037) );
  inv01 U1270 ( .Y(n3031), .A(n3040) );
  nand02 U1271 ( .Y(n3041), .A0(n3038), .A1(n3039) );
  inv01 U1272 ( .Y(n3032), .A(n3041) );
  nand02 U1273 ( .Y(fracta_52_o[42]), .A0(n3042), .A1(n3043) );
  inv01 U1274 ( .Y(n3044), .A(n3801) );
  inv01 U1275 ( .Y(n3045), .A(n3886) );
  inv01 U1276 ( .Y(n3046), .A(n3360) );
  nand02 U1277 ( .Y(n3047), .A0(n3769), .A1(n3044) );
  nand02 U1278 ( .Y(n3048), .A0(n3769), .A1(n3045) );
  nand02 U1279 ( .Y(n3049), .A0(n3044), .A1(n3046) );
  nand02 U1280 ( .Y(n3050), .A0(n3045), .A1(n3046) );
  nand02 U1281 ( .Y(n3051), .A0(n3047), .A1(n3048) );
  inv01 U1282 ( .Y(n3042), .A(n3051) );
  nand02 U1283 ( .Y(n3052), .A0(n3049), .A1(n3050) );
  inv01 U1284 ( .Y(n3043), .A(n3052) );
  nand02 U1285 ( .Y(n3053), .A0(n3987), .A1(n3905) );
  inv02 U1286 ( .Y(n3054), .A(n3053) );
  ao21 U1287 ( .Y(n3055), .A0(n3792), .A1(n3856), .B0(n3900) );
  inv01 U1288 ( .Y(n3056), .A(n3055) );
  nand02 U1289 ( .Y(fracta_52_o[43]), .A0(n3057), .A1(n3058) );
  inv01 U1290 ( .Y(n3059), .A(n3801) );
  inv01 U1291 ( .Y(n3060), .A(n3360) );
  inv01 U1292 ( .Y(n3061), .A(n3875) );
  nand02 U1293 ( .Y(n3062), .A0(n3769), .A1(n3059) );
  nand02 U1294 ( .Y(n3063), .A0(n3769), .A1(n3060) );
  nand02 U1295 ( .Y(n3064), .A0(n3059), .A1(n3061) );
  nand02 U1296 ( .Y(n3065), .A0(n3060), .A1(n3061) );
  nand02 U1297 ( .Y(n3066), .A0(n3062), .A1(n3063) );
  inv01 U1298 ( .Y(n3057), .A(n3066) );
  nand02 U1299 ( .Y(n3067), .A0(n3064), .A1(n3065) );
  inv01 U1300 ( .Y(n3058), .A(n3067) );
  nand02 U1301 ( .Y(fracta_52_o[38]), .A0(n3068), .A1(n3069) );
  inv01 U1302 ( .Y(n3070), .A(n3801) );
  inv01 U1303 ( .Y(n3071), .A(n3904) );
  inv01 U1304 ( .Y(n3072), .A(n3899) );
  nand02 U1305 ( .Y(n3073), .A0(n3801), .A1(n3070) );
  nand02 U1306 ( .Y(n3074), .A0(n3801), .A1(n3071) );
  nand02 U1307 ( .Y(n3075), .A0(n3070), .A1(n3072) );
  nand02 U1308 ( .Y(n3076), .A0(n3071), .A1(n3072) );
  nand02 U1309 ( .Y(n3077), .A0(n3073), .A1(n3074) );
  inv01 U1310 ( .Y(n3068), .A(n3077) );
  nand02 U1311 ( .Y(n3078), .A0(n3075), .A1(n3076) );
  inv01 U1312 ( .Y(n3069), .A(n3078) );
  nand02 U1313 ( .Y(fracta_52_o[41]), .A0(n3079), .A1(n3080) );
  inv01 U1314 ( .Y(n3081), .A(n3801) );
  inv01 U1315 ( .Y(n3082), .A(n3892) );
  inv01 U1316 ( .Y(n3083), .A(n3886) );
  nand02 U1317 ( .Y(n3084), .A0(n3769), .A1(n3081) );
  nand02 U1318 ( .Y(n3085), .A0(n3769), .A1(n3082) );
  nand02 U1319 ( .Y(n3086), .A0(n3081), .A1(n3083) );
  nand02 U1320 ( .Y(n3087), .A0(n3082), .A1(n3083) );
  nand02 U1321 ( .Y(n3088), .A0(n3084), .A1(n3085) );
  inv01 U1322 ( .Y(n3079), .A(n3088) );
  nand02 U1323 ( .Y(n3089), .A0(n3086), .A1(n3087) );
  inv01 U1324 ( .Y(n3080), .A(n3089) );
  nand02 U1325 ( .Y(fracta_52_o[37]), .A0(n3090), .A1(n3091) );
  inv01 U1326 ( .Y(n3092), .A(n3801) );
  inv01 U1327 ( .Y(n3093), .A(n3907) );
  inv01 U1328 ( .Y(n3094), .A(n3904) );
  nand02 U1329 ( .Y(n3095), .A0(n3769), .A1(n3092) );
  nand02 U1330 ( .Y(n3096), .A0(n3769), .A1(n3093) );
  nand02 U1331 ( .Y(n3097), .A0(n3092), .A1(n3094) );
  nand02 U1332 ( .Y(n3098), .A0(n3093), .A1(n3094) );
  nand02 U1333 ( .Y(n3099), .A0(n3095), .A1(n3096) );
  inv01 U1334 ( .Y(n3090), .A(n3099) );
  nand02 U1335 ( .Y(n3100), .A0(n3097), .A1(n3098) );
  inv01 U1336 ( .Y(n3091), .A(n3100) );
  buf02 U1337 ( .Y(n3101), .A(n3973) );
  nor02 U1338 ( .Y(n3981), .A0(n3102), .A1(n3103) );
  nor02 U1339 ( .Y(n3104), .A0(n3986), .A1(n3925) );
  inv01 U1340 ( .Y(n3102), .A(n3104) );
  nor02 U1341 ( .Y(n3105), .A0(n3924), .A1(n3331) );
  inv01 U1342 ( .Y(n3103), .A(n3105) );
  or02 U1343 ( .Y(n3106), .A0(n3994), .A1(opa_i[26]) );
  inv01 U1344 ( .Y(n3107), .A(n3106) );
  or02 U1345 ( .Y(n3108), .A0(n3995), .A1(opa_i[25]) );
  inv01 U1346 ( .Y(n3109), .A(n3108) );
  or02 U1347 ( .Y(n3110), .A0(n3993), .A1(opa_i[28]) );
  inv01 U1348 ( .Y(n3111), .A(n3110) );
  nor02 U1349 ( .Y(n3982), .A0(n3112), .A1(n3113) );
  nor02 U1350 ( .Y(n3114), .A0(n3983), .A1(n3926) );
  inv01 U1351 ( .Y(n3112), .A(n3114) );
  nor02 U1352 ( .Y(n3115), .A0(n3928), .A1(n3927) );
  inv01 U1353 ( .Y(n3113), .A(n3115) );
  or02 U1354 ( .Y(n3116), .A0(n3794), .A1(n3749) );
  inv01 U1355 ( .Y(n3117), .A(n3116) );
  buf02 U1356 ( .Y(n3118), .A(opa_i[11]) );
  inv01 U1357 ( .Y(n3119), .A(n3118) );
  nand02 U1358 ( .Y(n3859), .A0(n3120), .A1(n3121) );
  inv02 U1359 ( .Y(n3122), .A(n3868) );
  inv02 U1360 ( .Y(n3123), .A(n3815) );
  inv02 U1361 ( .Y(n3124), .A(n3813) );
  inv02 U1362 ( .Y(n3125), .A(n3811) );
  inv02 U1363 ( .Y(n3126), .A(n3814) );
  inv02 U1364 ( .Y(n3127), .A(n3816) );
  nand02 U1365 ( .Y(n3128), .A0(n3124), .A1(n3129) );
  nand02 U1366 ( .Y(n3130), .A0(n3125), .A1(n3131) );
  nand02 U1367 ( .Y(n3132), .A0(n3126), .A1(n3133) );
  nand02 U1368 ( .Y(n3134), .A0(n3126), .A1(n3135) );
  nand02 U1369 ( .Y(n3136), .A0(n3127), .A1(n3137) );
  nand02 U1370 ( .Y(n3138), .A0(n3127), .A1(n3139) );
  nand02 U1371 ( .Y(n3140), .A0(n3127), .A1(n3141) );
  nand02 U1372 ( .Y(n3142), .A0(n3127), .A1(n3143) );
  nand02 U1373 ( .Y(n3144), .A0(n3122), .A1(n3123) );
  inv01 U1374 ( .Y(n3129), .A(n3144) );
  nand02 U1375 ( .Y(n3145), .A0(n3122), .A1(n3123) );
  inv01 U1376 ( .Y(n3131), .A(n3145) );
  nand02 U1377 ( .Y(n3146), .A0(n3122), .A1(n3124) );
  inv01 U1378 ( .Y(n3133), .A(n3146) );
  nand02 U1379 ( .Y(n3147), .A0(n3122), .A1(n3125) );
  inv01 U1380 ( .Y(n3135), .A(n3147) );
  nand02 U1381 ( .Y(n3148), .A0(n3123), .A1(n3124) );
  inv01 U1382 ( .Y(n3137), .A(n3148) );
  nand02 U1383 ( .Y(n3149), .A0(n3123), .A1(n3125) );
  inv01 U1384 ( .Y(n3139), .A(n3149) );
  nand02 U1385 ( .Y(n3150), .A0(n3124), .A1(n3126) );
  inv01 U1386 ( .Y(n3141), .A(n3150) );
  nand02 U1387 ( .Y(n3151), .A0(n3125), .A1(n3126) );
  inv01 U1388 ( .Y(n3143), .A(n3151) );
  nand02 U1389 ( .Y(n3152), .A0(n3128), .A1(n3130) );
  inv01 U1390 ( .Y(n3153), .A(n3152) );
  nand02 U1391 ( .Y(n3154), .A0(n3132), .A1(n3134) );
  inv01 U1392 ( .Y(n3155), .A(n3154) );
  nand02 U1393 ( .Y(n3156), .A0(n3153), .A1(n3155) );
  inv01 U1394 ( .Y(n3120), .A(n3156) );
  nand02 U1395 ( .Y(n3157), .A0(n3136), .A1(n3138) );
  inv01 U1396 ( .Y(n3158), .A(n3157) );
  nand02 U1397 ( .Y(n3159), .A0(n3140), .A1(n3142) );
  inv01 U1398 ( .Y(n3160), .A(n3159) );
  nand02 U1399 ( .Y(n3161), .A0(n3158), .A1(n3160) );
  inv01 U1400 ( .Y(n3121), .A(n3161) );
  nand02 U1401 ( .Y(n3871), .A0(n3162), .A1(n3163) );
  inv02 U1402 ( .Y(n3164), .A(n3874) );
  inv02 U1403 ( .Y(n3165), .A(n3835) );
  inv02 U1404 ( .Y(n3166), .A(n3836) );
  inv02 U1405 ( .Y(n3167), .A(n3811) );
  inv02 U1406 ( .Y(n3168), .A(n3814) );
  inv02 U1407 ( .Y(n3169), .A(n3816) );
  nand02 U1408 ( .Y(n3170), .A0(n3166), .A1(n3171) );
  nand02 U1409 ( .Y(n3172), .A0(n3167), .A1(n3173) );
  nand02 U1410 ( .Y(n3174), .A0(n3168), .A1(n3175) );
  nand02 U1411 ( .Y(n3176), .A0(n3168), .A1(n3177) );
  nand02 U1412 ( .Y(n3178), .A0(n3169), .A1(n3179) );
  nand02 U1413 ( .Y(n3180), .A0(n3169), .A1(n3181) );
  nand02 U1414 ( .Y(n3182), .A0(n3169), .A1(n3183) );
  nand02 U1415 ( .Y(n3184), .A0(n3169), .A1(n3185) );
  nand02 U1416 ( .Y(n3186), .A0(n3164), .A1(n3165) );
  inv01 U1417 ( .Y(n3171), .A(n3186) );
  nand02 U1418 ( .Y(n3187), .A0(n3164), .A1(n3165) );
  inv01 U1419 ( .Y(n3173), .A(n3187) );
  nand02 U1420 ( .Y(n3188), .A0(n3164), .A1(n3166) );
  inv01 U1421 ( .Y(n3175), .A(n3188) );
  nand02 U1422 ( .Y(n3189), .A0(n3164), .A1(n3167) );
  inv01 U1423 ( .Y(n3177), .A(n3189) );
  nand02 U1424 ( .Y(n3190), .A0(n3165), .A1(n3166) );
  inv01 U1425 ( .Y(n3179), .A(n3190) );
  nand02 U1426 ( .Y(n3191), .A0(n3165), .A1(n3167) );
  inv01 U1427 ( .Y(n3181), .A(n3191) );
  nand02 U1428 ( .Y(n3192), .A0(n3166), .A1(n3168) );
  inv01 U1429 ( .Y(n3183), .A(n3192) );
  nand02 U1430 ( .Y(n3193), .A0(n3167), .A1(n3168) );
  inv01 U1431 ( .Y(n3185), .A(n3193) );
  nand02 U1432 ( .Y(n3194), .A0(n3170), .A1(n3172) );
  inv01 U1433 ( .Y(n3195), .A(n3194) );
  nand02 U1434 ( .Y(n3196), .A0(n3174), .A1(n3176) );
  inv01 U1435 ( .Y(n3197), .A(n3196) );
  nand02 U1436 ( .Y(n3198), .A0(n3195), .A1(n3197) );
  inv01 U1437 ( .Y(n3162), .A(n3198) );
  nand02 U1438 ( .Y(n3199), .A0(n3178), .A1(n3180) );
  inv01 U1439 ( .Y(n3200), .A(n3199) );
  nand02 U1440 ( .Y(n3201), .A0(n3182), .A1(n3184) );
  inv01 U1441 ( .Y(n3202), .A(n3201) );
  nand02 U1442 ( .Y(n3203), .A0(n3200), .A1(n3202) );
  inv01 U1443 ( .Y(n3163), .A(n3203) );
  nand02 U1444 ( .Y(n3881), .A0(n3204), .A1(n3205) );
  inv02 U1445 ( .Y(n3206), .A(n3885) );
  inv02 U1446 ( .Y(n3207), .A(n3856) );
  inv02 U1447 ( .Y(n3208), .A(n3884) );
  inv02 U1448 ( .Y(n3209), .A(n3811) );
  inv02 U1449 ( .Y(n3210), .A(n3814) );
  inv02 U1450 ( .Y(n3211), .A(n3816) );
  nand02 U1451 ( .Y(n3212), .A0(n3208), .A1(n3213) );
  nand02 U1452 ( .Y(n3214), .A0(n3209), .A1(n3215) );
  nand02 U1453 ( .Y(n3216), .A0(n3210), .A1(n3217) );
  nand02 U1454 ( .Y(n3218), .A0(n3210), .A1(n3219) );
  nand02 U1455 ( .Y(n3220), .A0(n3211), .A1(n3221) );
  nand02 U1456 ( .Y(n3222), .A0(n3211), .A1(n3223) );
  nand02 U1457 ( .Y(n3224), .A0(n3211), .A1(n3225) );
  nand02 U1458 ( .Y(n3226), .A0(n3211), .A1(n3227) );
  nand02 U1459 ( .Y(n3228), .A0(n3206), .A1(n3207) );
  inv01 U1460 ( .Y(n3213), .A(n3228) );
  nand02 U1461 ( .Y(n3229), .A0(n3206), .A1(n3207) );
  inv01 U1462 ( .Y(n3215), .A(n3229) );
  nand02 U1463 ( .Y(n3230), .A0(n3206), .A1(n3208) );
  inv01 U1464 ( .Y(n3217), .A(n3230) );
  nand02 U1465 ( .Y(n3231), .A0(n3206), .A1(n3209) );
  inv01 U1466 ( .Y(n3219), .A(n3231) );
  nand02 U1467 ( .Y(n3232), .A0(n3207), .A1(n3208) );
  inv01 U1468 ( .Y(n3221), .A(n3232) );
  nand02 U1469 ( .Y(n3233), .A0(n3207), .A1(n3209) );
  inv01 U1470 ( .Y(n3223), .A(n3233) );
  nand02 U1471 ( .Y(n3234), .A0(n3208), .A1(n3210) );
  inv01 U1472 ( .Y(n3225), .A(n3234) );
  nand02 U1473 ( .Y(n3235), .A0(n3209), .A1(n3210) );
  inv01 U1474 ( .Y(n3227), .A(n3235) );
  nand02 U1475 ( .Y(n3236), .A0(n3212), .A1(n3214) );
  inv01 U1476 ( .Y(n3237), .A(n3236) );
  nand02 U1477 ( .Y(n3238), .A0(n3216), .A1(n3218) );
  inv01 U1478 ( .Y(n3239), .A(n3238) );
  nand02 U1479 ( .Y(n3240), .A0(n3237), .A1(n3239) );
  inv01 U1480 ( .Y(n3204), .A(n3240) );
  nand02 U1481 ( .Y(n3241), .A0(n3220), .A1(n3222) );
  inv01 U1482 ( .Y(n3242), .A(n3241) );
  nand02 U1483 ( .Y(n3243), .A0(n3224), .A1(n3226) );
  inv01 U1484 ( .Y(n3244), .A(n3243) );
  nand02 U1485 ( .Y(n3245), .A0(n3242), .A1(n3244) );
  inv01 U1486 ( .Y(n3205), .A(n3245) );
  nand02 U1487 ( .Y(n3877), .A0(n3246), .A1(n3247) );
  inv02 U1488 ( .Y(n3248), .A(n3879) );
  inv02 U1489 ( .Y(n3249), .A(n3845) );
  inv02 U1490 ( .Y(n3250), .A(n3846) );
  inv02 U1491 ( .Y(n3251), .A(n3811) );
  inv02 U1492 ( .Y(n3252), .A(n3814) );
  inv02 U1493 ( .Y(n3253), .A(n3816) );
  nand02 U1494 ( .Y(n3254), .A0(n3250), .A1(n3255) );
  nand02 U1495 ( .Y(n3256), .A0(n3251), .A1(n3257) );
  nand02 U1496 ( .Y(n3258), .A0(n3252), .A1(n3259) );
  nand02 U1497 ( .Y(n3260), .A0(n3252), .A1(n3261) );
  nand02 U1498 ( .Y(n3262), .A0(n3253), .A1(n3263) );
  nand02 U1499 ( .Y(n3264), .A0(n3253), .A1(n3265) );
  nand02 U1500 ( .Y(n3266), .A0(n3253), .A1(n3267) );
  nand02 U1501 ( .Y(n3268), .A0(n3253), .A1(n3269) );
  nand02 U1502 ( .Y(n3270), .A0(n3248), .A1(n3249) );
  inv01 U1503 ( .Y(n3255), .A(n3270) );
  nand02 U1504 ( .Y(n3271), .A0(n3248), .A1(n3249) );
  inv01 U1505 ( .Y(n3257), .A(n3271) );
  nand02 U1506 ( .Y(n3272), .A0(n3248), .A1(n3250) );
  inv01 U1507 ( .Y(n3259), .A(n3272) );
  nand02 U1508 ( .Y(n3273), .A0(n3248), .A1(n3251) );
  inv01 U1509 ( .Y(n3261), .A(n3273) );
  nand02 U1510 ( .Y(n3274), .A0(n3249), .A1(n3250) );
  inv01 U1511 ( .Y(n3263), .A(n3274) );
  nand02 U1512 ( .Y(n3275), .A0(n3249), .A1(n3251) );
  inv01 U1513 ( .Y(n3265), .A(n3275) );
  nand02 U1514 ( .Y(n3276), .A0(n3250), .A1(n3252) );
  inv01 U1515 ( .Y(n3267), .A(n3276) );
  nand02 U1516 ( .Y(n3277), .A0(n3251), .A1(n3252) );
  inv01 U1517 ( .Y(n3269), .A(n3277) );
  nand02 U1518 ( .Y(n3278), .A0(n3254), .A1(n3256) );
  inv01 U1519 ( .Y(n3279), .A(n3278) );
  nand02 U1520 ( .Y(n3280), .A0(n3258), .A1(n3260) );
  inv01 U1521 ( .Y(n3281), .A(n3280) );
  nand02 U1522 ( .Y(n3282), .A0(n3279), .A1(n3281) );
  inv01 U1523 ( .Y(n3246), .A(n3282) );
  nand02 U1524 ( .Y(n3283), .A0(n3262), .A1(n3264) );
  inv01 U1525 ( .Y(n3284), .A(n3283) );
  nand02 U1526 ( .Y(n3285), .A0(n3266), .A1(n3268) );
  inv01 U1527 ( .Y(n3286), .A(n3285) );
  nand02 U1528 ( .Y(n3287), .A0(n3284), .A1(n3286) );
  inv01 U1529 ( .Y(n3247), .A(n3287) );
  or02 U1530 ( .Y(n3288), .A0(n3804), .A1(opa_i[27]) );
  inv01 U1531 ( .Y(n3289), .A(n3288) );
  inv01 U1532 ( .Y(n3900), .A(n3290) );
  nor02 U1533 ( .Y(n3291), .A0(n3771), .A1(n3292) );
  nor02 U1534 ( .Y(n3293), .A0(n3854), .A1(n3789) );
  nor02 U1535 ( .Y(n3290), .A0(n3291), .A1(n3293) );
  nor02 U1536 ( .Y(n3294), .A0(n3794), .A1(n3901) );
  inv01 U1537 ( .Y(n3292), .A(n3294) );
  buf02 U1538 ( .Y(n3295), .A(n3839) );
  inv02 U1539 ( .Y(n3975), .A(n3296) );
  nand02 U1540 ( .Y(n3296), .A0(n2742), .A1(n3297) );
  nand02 U1541 ( .Y(n3298), .A0(n3119), .A1(n3758) );
  inv01 U1542 ( .Y(n3297), .A(n3298) );
  nand02 U1543 ( .Y(n3986), .A0(n3299), .A1(n3300) );
  inv01 U1544 ( .Y(n3301), .A(n3972) );
  inv01 U1545 ( .Y(n3303), .A(n3601) );
  inv01 U1546 ( .Y(n3304), .A(n3817) );
  inv01 U1547 ( .Y(n3305), .A(n3988) );
  nand02 U1548 ( .Y(n3299), .A0(n3303), .A1(n3306) );
  nand02 U1549 ( .Y(n3300), .A0(n3304), .A1(n3305) );
  nand02 U1550 ( .Y(n3307), .A0(n3301), .A1(n3302) );
  inv01 U1551 ( .Y(n3306), .A(n3307) );
  buf02 U1552 ( .Y(n3308), .A(opa_i[2]) );
  inv02 U1553 ( .Y(n3309), .A(n3308) );
  buf02 U1554 ( .Y(n3780), .A(n3872) );
  buf02 U1555 ( .Y(n3310), .A(n3822) );
  inv02 U1556 ( .Y(n3905), .A(opa_i[8]) );
  buf02 U1557 ( .Y(n3311), .A(opa_i[5]) );
  inv02 U1558 ( .Y(n3312), .A(n3311) );
  buf02 U1559 ( .Y(n3313), .A(n3850) );
  inv02 U1560 ( .Y(n____return1466_2_), .A(n3314) );
  inv01 U1561 ( .Y(n3315), .A(n3995) );
  inv01 U1562 ( .Y(n3316), .A(opa_i[25]) );
  nor02 U1563 ( .Y(n3317), .A0(n3315), .A1(n3316) );
  nor02 U1564 ( .Y(n3314), .A0(n3317), .A1(n3109) );
  inv02 U1565 ( .Y(n____return1466_1_), .A(n3318) );
  inv01 U1566 ( .Y(n3319), .A(opa_i[23]) );
  inv01 U1567 ( .Y(n3320), .A(opa_i[24]) );
  nor02 U1568 ( .Y(n3321), .A0(n3319), .A1(n3320) );
  nor02 U1569 ( .Y(n3318), .A0(n3321), .A1(n3347) );
  inv02 U1570 ( .Y(n1468_4_), .A(n3322) );
  inv01 U1571 ( .Y(n3323), .A(n3804) );
  inv01 U1572 ( .Y(n3324), .A(opa_i[27]) );
  nor02 U1573 ( .Y(n3325), .A0(n3323), .A1(n3324) );
  nor02 U1574 ( .Y(n3322), .A0(n3325), .A1(n3289) );
  inv02 U1575 ( .Y(n____return1466_3_), .A(n3326) );
  inv01 U1576 ( .Y(n3327), .A(n3994) );
  inv01 U1577 ( .Y(n3328), .A(opa_i[26]) );
  nor02 U1578 ( .Y(n3329), .A0(n3327), .A1(n3328) );
  nor02 U1579 ( .Y(n3326), .A0(n3329), .A1(n3107) );
  nand02 U1580 ( .Y(n3330), .A0(opa_i[8]), .A1(n3987) );
  inv02 U1581 ( .Y(n3331), .A(n3330) );
  nand02 U1582 ( .Y(fracta_52_o[32]), .A0(n3332), .A1(n3333) );
  inv01 U1583 ( .Y(n3334), .A(n3771) );
  inv01 U1584 ( .Y(n3335), .A(n3781) );
  inv01 U1585 ( .Y(n3336), .A(n3775) );
  inv01 U1586 ( .Y(n3337), .A(n3611) );
  inv01 U1587 ( .Y(n3338), .A(n____return1466_0_) );
  nand02 U1588 ( .Y(n3332), .A0(n3336), .A1(n3339) );
  nand02 U1589 ( .Y(n3333), .A0(n3337), .A1(n3338) );
  nand02 U1590 ( .Y(n3340), .A0(n3334), .A1(n3335) );
  inv01 U1591 ( .Y(n3339), .A(n3340) );
  buf04 U1592 ( .Y(n3781), .A(s_sqr_zeros_o_3_) );
  inv01 U1593 ( .Y(fracta_52_o[51]), .A(n3341) );
  nor02 U1594 ( .Y(n3342), .A0(n3699), .A1(n3343) );
  nor02 U1595 ( .Y(n3344), .A0(n3807), .A1(n3775) );
  nor02 U1596 ( .Y(n3341), .A0(n3342), .A1(n3344) );
  nor02 U1597 ( .Y(n3345), .A0(n3805), .A1(n3806) );
  inv01 U1598 ( .Y(n3343), .A(n3345) );
  buf02 U1599 ( .Y(n3775), .A(n3808) );
  or02 U1600 ( .Y(n3346), .A0(opa_i[24]), .A1(opa_i[23]) );
  inv01 U1601 ( .Y(n3347), .A(n3346) );
  inv01 U1602 ( .Y(n3807), .A(n3348) );
  inv01 U1603 ( .Y(n3349), .A(opa_i[21]) );
  inv01 U1604 ( .Y(n3350), .A(opa_i[22]) );
  inv01 U1605 ( .Y(n3351), .A(n3810) );
  inv01 U1606 ( .Y(n3352), .A(n3809) );
  nand02 U1607 ( .Y(n3348), .A0(n3353), .A1(n3354) );
  nand02 U1608 ( .Y(n3355), .A0(n3349), .A1(n3350) );
  inv01 U1609 ( .Y(n3353), .A(n3355) );
  nand02 U1610 ( .Y(n3356), .A0(n3351), .A1(n3352) );
  inv01 U1611 ( .Y(n3354), .A(n3356) );
  xor2 U1612 ( .Y(n3357), .A0(n3774), .A1(opa_i[30]) );
  ao221 U1613 ( .Y(n3359), .A0(n3815), .A1(n3792), .B0(n3868), .B1(n3788), 
        .C0(n3889) );
  inv01 U1614 ( .Y(n3360), .A(n3359) );
  nand02 U1615 ( .Y(n3892), .A0(n3361), .A1(n3362) );
  inv02 U1616 ( .Y(n3363), .A(n3896) );
  inv01 U1617 ( .Y(n3364), .A(n3788) );
  inv01 U1618 ( .Y(n3365), .A(n3792) );
  inv01 U1619 ( .Y(n3366), .A(n3845) );
  inv01 U1620 ( .Y(n3367), .A(n3879) );
  nand02 U1621 ( .Y(n3368), .A0(n3365), .A1(n3369) );
  nand02 U1622 ( .Y(n3370), .A0(n3366), .A1(n3371) );
  nand02 U1623 ( .Y(n3372), .A0(n3367), .A1(n3373) );
  nand02 U1624 ( .Y(n3374), .A0(n3367), .A1(n3375) );
  nand02 U1625 ( .Y(n3376), .A0(n3363), .A1(n3364) );
  inv01 U1626 ( .Y(n3369), .A(n3376) );
  nand02 U1627 ( .Y(n3377), .A0(n3363), .A1(n3364) );
  inv01 U1628 ( .Y(n3371), .A(n3377) );
  nand02 U1629 ( .Y(n3378), .A0(n3363), .A1(n3365) );
  inv01 U1630 ( .Y(n3373), .A(n3378) );
  nand02 U1631 ( .Y(n3379), .A0(n3363), .A1(n3366) );
  inv01 U1632 ( .Y(n3375), .A(n3379) );
  nand02 U1633 ( .Y(n3380), .A0(n3368), .A1(n3370) );
  inv01 U1634 ( .Y(n3361), .A(n3380) );
  nand02 U1635 ( .Y(n3381), .A0(n3372), .A1(n3374) );
  inv01 U1636 ( .Y(n3362), .A(n3381) );
  nand02 U1637 ( .Y(n3886), .A0(n3382), .A1(n3383) );
  inv02 U1638 ( .Y(n3384), .A(n3893) );
  inv01 U1639 ( .Y(n3385), .A(n3788) );
  inv01 U1640 ( .Y(n3386), .A(n3792) );
  inv01 U1641 ( .Y(n3387), .A(n3835) );
  inv01 U1642 ( .Y(n3388), .A(n3874) );
  nand02 U1643 ( .Y(n3389), .A0(n3386), .A1(n3390) );
  nand02 U1644 ( .Y(n3391), .A0(n3387), .A1(n3392) );
  nand02 U1645 ( .Y(n3393), .A0(n3388), .A1(n3394) );
  nand02 U1646 ( .Y(n3395), .A0(n3388), .A1(n3396) );
  nand02 U1647 ( .Y(n3397), .A0(n3384), .A1(n3385) );
  inv01 U1648 ( .Y(n3390), .A(n3397) );
  nand02 U1649 ( .Y(n3398), .A0(n3384), .A1(n3385) );
  inv01 U1650 ( .Y(n3392), .A(n3398) );
  nand02 U1651 ( .Y(n3399), .A0(n3384), .A1(n3386) );
  inv01 U1652 ( .Y(n3394), .A(n3399) );
  nand02 U1653 ( .Y(n3400), .A0(n3384), .A1(n3387) );
  inv01 U1654 ( .Y(n3396), .A(n3400) );
  nand02 U1655 ( .Y(n3401), .A0(n3389), .A1(n3391) );
  inv01 U1656 ( .Y(n3382), .A(n3401) );
  nand02 U1657 ( .Y(n3402), .A0(n3393), .A1(n3395) );
  inv01 U1658 ( .Y(n3383), .A(n3402) );
  nand02 U1659 ( .Y(n3812), .A0(n3867), .A1(n3403) );
  inv01 U1660 ( .Y(n3404), .A(n3798) );
  inv01 U1661 ( .Y(n3405), .A(n3865) );
  inv01 U1662 ( .Y(n3406), .A(n3795) );
  inv01 U1663 ( .Y(n3407), .A(n3638) );
  nand02 U1664 ( .Y(n3408), .A0(n3404), .A1(n3405) );
  nand02 U1665 ( .Y(n3409), .A0(n3406), .A1(n3407) );
  nand02 U1666 ( .Y(n3410), .A0(n3408), .A1(n3409) );
  inv01 U1667 ( .Y(n3403), .A(n3410) );
  inv02 U1668 ( .Y(n3884), .A(n3411) );
  nor02 U1669 ( .Y(n3412), .A0(n3754), .A1(n3797) );
  nor02 U1670 ( .Y(n3413), .A0(n3902), .A1(n3795) );
  inv01 U1671 ( .Y(n3414), .A(n3903) );
  nor02 U1672 ( .Y(n3411), .A0(n3414), .A1(n3415) );
  nor02 U1673 ( .Y(n3416), .A0(n3412), .A1(n3413) );
  inv01 U1674 ( .Y(n3415), .A(n3416) );
  inv02 U1675 ( .Y(n3854), .A(n3884) );
  buf04 U1676 ( .Y(n3795), .A(n3864) );
  inv01 U1677 ( .Y(n3978), .A(n3417) );
  inv01 U1678 ( .Y(n3418), .A(n3974) );
  nand02 U1679 ( .Y(n3417), .A0(n3984), .A1(n3420) );
  nand02 U1680 ( .Y(n3421), .A0(n3418), .A1(n3419) );
  inv01 U1681 ( .Y(n3420), .A(n3421) );
  inv01 U1682 ( .Y(n3927), .A(n3422) );
  inv01 U1683 ( .Y(n3423), .A(n3984) );
  inv01 U1684 ( .Y(n3424), .A(n3974) );
  nand02 U1685 ( .Y(n3422), .A0(n3424), .A1(n3425) );
  nand02 U1686 ( .Y(n3426), .A0(n3423), .A1(n3419) );
  inv01 U1687 ( .Y(n3425), .A(n3426) );
  nand02 U1688 ( .Y(n3907), .A0(n3427), .A1(n3428) );
  inv02 U1689 ( .Y(n3429), .A(n3792) );
  inv02 U1690 ( .Y(n3430), .A(n3790) );
  inv02 U1691 ( .Y(n3431), .A(n3788) );
  inv02 U1692 ( .Y(n3432), .A(n3897) );
  inv02 U1693 ( .Y(n3433), .A(n3845) );
  inv02 U1694 ( .Y(n3434), .A(n3879) );
  nand02 U1695 ( .Y(n3435), .A0(n3431), .A1(n3436) );
  nand02 U1696 ( .Y(n3437), .A0(n3432), .A1(n3438) );
  nand02 U1697 ( .Y(n3439), .A0(n3433), .A1(n3440) );
  nand02 U1698 ( .Y(n3441), .A0(n3433), .A1(n3442) );
  nand02 U1699 ( .Y(n3443), .A0(n3434), .A1(n3444) );
  nand02 U1700 ( .Y(n3445), .A0(n3434), .A1(n3446) );
  nand02 U1701 ( .Y(n3447), .A0(n3434), .A1(n3448) );
  nand02 U1702 ( .Y(n3449), .A0(n3434), .A1(n3450) );
  nand02 U1703 ( .Y(n3451), .A0(n3429), .A1(n3430) );
  inv01 U1704 ( .Y(n3436), .A(n3451) );
  nand02 U1705 ( .Y(n3452), .A0(n3429), .A1(n3430) );
  inv01 U1706 ( .Y(n3438), .A(n3452) );
  nand02 U1707 ( .Y(n3453), .A0(n3429), .A1(n3431) );
  inv01 U1708 ( .Y(n3440), .A(n3453) );
  nand02 U1709 ( .Y(n3454), .A0(n3429), .A1(n3432) );
  inv01 U1710 ( .Y(n3442), .A(n3454) );
  nand02 U1711 ( .Y(n3455), .A0(n3430), .A1(n3431) );
  inv01 U1712 ( .Y(n3444), .A(n3455) );
  nand02 U1713 ( .Y(n3456), .A0(n3430), .A1(n3432) );
  inv01 U1714 ( .Y(n3446), .A(n3456) );
  nand02 U1715 ( .Y(n3457), .A0(n3431), .A1(n3433) );
  inv01 U1716 ( .Y(n3448), .A(n3457) );
  nand02 U1717 ( .Y(n3458), .A0(n3432), .A1(n3433) );
  inv01 U1718 ( .Y(n3450), .A(n3458) );
  nand02 U1719 ( .Y(n3459), .A0(n3435), .A1(n3437) );
  inv01 U1720 ( .Y(n3460), .A(n3459) );
  nand02 U1721 ( .Y(n3461), .A0(n3439), .A1(n3441) );
  inv01 U1722 ( .Y(n3462), .A(n3461) );
  nand02 U1723 ( .Y(n3463), .A0(n3460), .A1(n3462) );
  inv01 U1724 ( .Y(n3427), .A(n3463) );
  nand02 U1725 ( .Y(n3464), .A0(n3443), .A1(n3445) );
  inv01 U1726 ( .Y(n3465), .A(n3464) );
  nand02 U1727 ( .Y(n3466), .A0(n3447), .A1(n3449) );
  inv01 U1728 ( .Y(n3467), .A(n3466) );
  nand02 U1729 ( .Y(n3468), .A0(n3465), .A1(n3467) );
  inv01 U1730 ( .Y(n3428), .A(n3468) );
  inv01 U1731 ( .Y(n3904), .A(n3469) );
  nor02 U1732 ( .Y(n3470), .A0(n3792), .A1(n3471) );
  nor02 U1733 ( .Y(n3472), .A0(n3792), .A1(n3473) );
  nor02 U1734 ( .Y(n3474), .A0(n3792), .A1(n3475) );
  nor02 U1735 ( .Y(n3476), .A0(n3792), .A1(n3477) );
  nor02 U1736 ( .Y(n3478), .A0(n3874), .A1(n3479) );
  nor02 U1737 ( .Y(n3480), .A0(n3874), .A1(n3481) );
  nor02 U1738 ( .Y(n3482), .A0(n3874), .A1(n3483) );
  nor02 U1739 ( .Y(n3484), .A0(n3874), .A1(n3485) );
  nor02 U1740 ( .Y(n3469), .A0(n3486), .A1(n3487) );
  nor02 U1741 ( .Y(n3488), .A0(n3788), .A1(n3790) );
  inv01 U1742 ( .Y(n3471), .A(n3488) );
  nor02 U1743 ( .Y(n3489), .A0(n3894), .A1(n3790) );
  inv01 U1744 ( .Y(n3473), .A(n3489) );
  nor02 U1745 ( .Y(n3490), .A0(n3788), .A1(n3835) );
  inv01 U1746 ( .Y(n3475), .A(n3490) );
  nor02 U1747 ( .Y(n3491), .A0(n3894), .A1(n3835) );
  inv01 U1748 ( .Y(n3477), .A(n3491) );
  nor02 U1749 ( .Y(n3492), .A0(n3788), .A1(n3790) );
  inv01 U1750 ( .Y(n3479), .A(n3492) );
  nor02 U1751 ( .Y(n3493), .A0(n3894), .A1(n3790) );
  inv01 U1752 ( .Y(n3481), .A(n3493) );
  nor02 U1753 ( .Y(n3494), .A0(n3788), .A1(n3835) );
  inv01 U1754 ( .Y(n3483), .A(n3494) );
  nor02 U1755 ( .Y(n3495), .A0(n3894), .A1(n3835) );
  inv01 U1756 ( .Y(n3485), .A(n3495) );
  nor02 U1757 ( .Y(n3496), .A0(n3470), .A1(n3472) );
  inv01 U1758 ( .Y(n3497), .A(n3496) );
  nor02 U1759 ( .Y(n3498), .A0(n3474), .A1(n3476) );
  inv01 U1760 ( .Y(n3499), .A(n3498) );
  nor02 U1761 ( .Y(n3500), .A0(n3497), .A1(n3499) );
  inv01 U1762 ( .Y(n3486), .A(n3500) );
  nor02 U1763 ( .Y(n3501), .A0(n3478), .A1(n3480) );
  inv01 U1764 ( .Y(n3502), .A(n3501) );
  nor02 U1765 ( .Y(n3503), .A0(n3482), .A1(n3484) );
  inv01 U1766 ( .Y(n3504), .A(n3503) );
  nor02 U1767 ( .Y(n3505), .A0(n3502), .A1(n3504) );
  inv01 U1768 ( .Y(n3487), .A(n3505) );
  nand02 U1769 ( .Y(n3899), .A0(n3506), .A1(n3507) );
  inv02 U1770 ( .Y(n3508), .A(n3792) );
  inv02 U1771 ( .Y(n3509), .A(n3790) );
  inv02 U1772 ( .Y(n3510), .A(n3788) );
  inv02 U1773 ( .Y(n3511), .A(n3890) );
  inv02 U1774 ( .Y(n3512), .A(n3815) );
  inv02 U1775 ( .Y(n3513), .A(n3868) );
  nand02 U1776 ( .Y(n3514), .A0(n3510), .A1(n3515) );
  nand02 U1777 ( .Y(n3516), .A0(n3511), .A1(n3517) );
  nand02 U1778 ( .Y(n3518), .A0(n3512), .A1(n3519) );
  nand02 U1779 ( .Y(n3520), .A0(n3512), .A1(n3521) );
  nand02 U1780 ( .Y(n3522), .A0(n3513), .A1(n3523) );
  nand02 U1781 ( .Y(n3524), .A0(n3513), .A1(n3525) );
  nand02 U1782 ( .Y(n3526), .A0(n3513), .A1(n3527) );
  nand02 U1783 ( .Y(n3528), .A0(n3513), .A1(n3529) );
  nand02 U1784 ( .Y(n3530), .A0(n3508), .A1(n3509) );
  inv01 U1785 ( .Y(n3515), .A(n3530) );
  nand02 U1786 ( .Y(n3531), .A0(n3508), .A1(n3509) );
  inv01 U1787 ( .Y(n3517), .A(n3531) );
  nand02 U1788 ( .Y(n3532), .A0(n3508), .A1(n3510) );
  inv01 U1789 ( .Y(n3519), .A(n3532) );
  nand02 U1790 ( .Y(n3533), .A0(n3508), .A1(n3511) );
  inv01 U1791 ( .Y(n3521), .A(n3533) );
  nand02 U1792 ( .Y(n3534), .A0(n3509), .A1(n3510) );
  inv01 U1793 ( .Y(n3523), .A(n3534) );
  nand02 U1794 ( .Y(n3535), .A0(n3509), .A1(n3511) );
  inv01 U1795 ( .Y(n3525), .A(n3535) );
  nand02 U1796 ( .Y(n3536), .A0(n3510), .A1(n3512) );
  inv01 U1797 ( .Y(n3527), .A(n3536) );
  nand02 U1798 ( .Y(n3537), .A0(n3511), .A1(n3512) );
  inv01 U1799 ( .Y(n3529), .A(n3537) );
  nand02 U1800 ( .Y(n3538), .A0(n3514), .A1(n3516) );
  inv01 U1801 ( .Y(n3539), .A(n3538) );
  nand02 U1802 ( .Y(n3540), .A0(n3518), .A1(n3520) );
  inv01 U1803 ( .Y(n3541), .A(n3540) );
  nand02 U1804 ( .Y(n3542), .A0(n3539), .A1(n3541) );
  inv01 U1805 ( .Y(n3506), .A(n3542) );
  nand02 U1806 ( .Y(n3543), .A0(n3522), .A1(n3524) );
  inv01 U1807 ( .Y(n3544), .A(n3543) );
  nand02 U1808 ( .Y(n3545), .A0(n3526), .A1(n3528) );
  inv01 U1809 ( .Y(n3546), .A(n3545) );
  nand02 U1810 ( .Y(n3547), .A0(n3544), .A1(n3546) );
  inv01 U1811 ( .Y(n3507), .A(n3547) );
  inv01 U1812 ( .Y(n3960), .A(n3548) );
  inv01 U1813 ( .Y(n3549), .A(opa_i[22]) );
  inv01 U1814 ( .Y(n3550), .A(n3990) );
  nand02 U1815 ( .Y(n3548), .A0(n3550), .A1(n3551) );
  nand02 U1816 ( .Y(n3552), .A0(n3304), .A1(n3549) );
  inv01 U1817 ( .Y(n3551), .A(n3552) );
  nand02 U1818 ( .Y(n3909), .A0(n3553), .A1(n3554) );
  inv02 U1819 ( .Y(n3555), .A(n3792) );
  inv02 U1820 ( .Y(n3556), .A(n3790) );
  inv02 U1821 ( .Y(n3557), .A(n3788) );
  inv02 U1822 ( .Y(n3558), .A(n3911) );
  inv02 U1823 ( .Y(n3559), .A(n3856) );
  inv02 U1824 ( .Y(n3560), .A(n3885) );
  nand02 U1825 ( .Y(n3561), .A0(n3557), .A1(n3562) );
  nand02 U1826 ( .Y(n3563), .A0(n3558), .A1(n3564) );
  nand02 U1827 ( .Y(n3565), .A0(n3559), .A1(n3566) );
  nand02 U1828 ( .Y(n3567), .A0(n3559), .A1(n3568) );
  nand02 U1829 ( .Y(n3569), .A0(n3560), .A1(n3570) );
  nand02 U1830 ( .Y(n3571), .A0(n3560), .A1(n3572) );
  nand02 U1831 ( .Y(n3573), .A0(n3560), .A1(n3574) );
  nand02 U1832 ( .Y(n3575), .A0(n3560), .A1(n3576) );
  nand02 U1833 ( .Y(n3577), .A0(n3555), .A1(n3556) );
  inv02 U1834 ( .Y(n3562), .A(n3577) );
  nand02 U1835 ( .Y(n3578), .A0(n3555), .A1(n3556) );
  inv01 U1836 ( .Y(n3564), .A(n3578) );
  nand02 U1837 ( .Y(n3579), .A0(n3555), .A1(n3557) );
  inv01 U1838 ( .Y(n3566), .A(n3579) );
  nand02 U1839 ( .Y(n3580), .A0(n3555), .A1(n3558) );
  inv01 U1840 ( .Y(n3568), .A(n3580) );
  nand02 U1841 ( .Y(n3581), .A0(n3556), .A1(n3557) );
  inv01 U1842 ( .Y(n3570), .A(n3581) );
  nand02 U1843 ( .Y(n3582), .A0(n3556), .A1(n3558) );
  inv01 U1844 ( .Y(n3572), .A(n3582) );
  nand02 U1845 ( .Y(n3583), .A0(n3557), .A1(n3559) );
  inv01 U1846 ( .Y(n3574), .A(n3583) );
  nand02 U1847 ( .Y(n3584), .A0(n3558), .A1(n3559) );
  inv01 U1848 ( .Y(n3576), .A(n3584) );
  nand02 U1849 ( .Y(n3585), .A0(n3561), .A1(n3563) );
  inv02 U1850 ( .Y(n3586), .A(n3585) );
  nand02 U1851 ( .Y(n3587), .A0(n3565), .A1(n3567) );
  inv02 U1852 ( .Y(n3588), .A(n3587) );
  nand02 U1853 ( .Y(n3589), .A0(n3586), .A1(n3588) );
  inv02 U1854 ( .Y(n3553), .A(n3589) );
  nand02 U1855 ( .Y(n3590), .A0(n3569), .A1(n3571) );
  inv01 U1856 ( .Y(n3591), .A(n3590) );
  nand02 U1857 ( .Y(n3592), .A0(n3573), .A1(n3575) );
  inv02 U1858 ( .Y(n3593), .A(n3592) );
  nand02 U1859 ( .Y(n3594), .A0(n3591), .A1(n3593) );
  inv02 U1860 ( .Y(n3554), .A(n3594) );
  ao22 U1861 ( .Y(n3595), .A0(n3894), .A1(n3811), .B0(n3874), .B1(n3764) );
  inv02 U1862 ( .Y(n3596), .A(n3595) );
  nand02 U1863 ( .Y(n3971), .A0(n3597), .A1(n3598) );
  inv01 U1864 ( .Y(n3599), .A(n3865) );
  inv01 U1865 ( .Y(n3600), .A(n3972) );
  inv01 U1866 ( .Y(n3602), .A(n3101) );
  inv01 U1867 ( .Y(n3603), .A(opa_i[22]) );
  nand02 U1868 ( .Y(n3597), .A0(n3604), .A1(n3605) );
  nand02 U1869 ( .Y(n3598), .A0(n3304), .A1(n3606) );
  nand02 U1870 ( .Y(n3607), .A0(n3599), .A1(n3600) );
  inv01 U1871 ( .Y(n3604), .A(n3607) );
  nand02 U1872 ( .Y(n3608), .A0(n3601), .A1(n3302) );
  inv01 U1873 ( .Y(n3605), .A(n3608) );
  nand02 U1874 ( .Y(n3609), .A0(n3602), .A1(n3603) );
  inv01 U1875 ( .Y(n3606), .A(n3609) );
  ao22 U1876 ( .Y(n3610), .A0(n3879), .A1(n3765), .B0(n3897), .B1(n3811) );
  inv02 U1877 ( .Y(n3611), .A(n3610) );
  inv02 U1878 ( .Y(n3972), .A(n3960) );
  buf02 U1879 ( .Y(n3614), .A(s_sqr_zeros_o_0_) );
  inv02 U1880 ( .Y(n3846), .A(n3615) );
  nor02 U1881 ( .Y(n3616), .A0(n3119), .A1(n3797) );
  nor02 U1882 ( .Y(n3617), .A0(n3754), .A1(n3795) );
  inv01 U1883 ( .Y(n3618), .A(n3898) );
  nor02 U1884 ( .Y(n3615), .A0(n3618), .A1(n3619) );
  nor02 U1885 ( .Y(n3620), .A0(n3616), .A1(n3617) );
  inv01 U1886 ( .Y(n3619), .A(n3620) );
  inv02 U1887 ( .Y(n3797), .A(n3796) );
  inv02 U1888 ( .Y(n3836), .A(n3621) );
  nor02 U1889 ( .Y(n3622), .A0(n3758), .A1(n3798) );
  nor02 U1890 ( .Y(n3623), .A0(n3119), .A1(n3795) );
  inv01 U1891 ( .Y(n3624), .A(n3895) );
  nor02 U1892 ( .Y(n3621), .A0(n3624), .A1(n3625) );
  nor02 U1893 ( .Y(n3626), .A0(n3622), .A1(n3623) );
  inv01 U1894 ( .Y(n3625), .A(n3626) );
  inv02 U1895 ( .Y(n3885), .A(n3627) );
  nor02 U1896 ( .Y(n3628), .A0(n3309), .A1(n3798) );
  nor02 U1897 ( .Y(n3629), .A0(n3919), .A1(n3795) );
  inv01 U1898 ( .Y(n3630), .A(n3920) );
  nor02 U1899 ( .Y(n3627), .A0(n3630), .A1(n3631) );
  nor02 U1900 ( .Y(n3632), .A0(n3628), .A1(n3629) );
  inv01 U1901 ( .Y(n3631), .A(n3632) );
  nand02 U1902 ( .Y(n3831), .A0(n3633), .A1(n3634) );
  inv02 U1903 ( .Y(n3635), .A(n3873) );
  inv01 U1904 ( .Y(n3636), .A(n3825) );
  inv01 U1905 ( .Y(n3637), .A(n3824) );
  nand02 U1906 ( .Y(n3639), .A0(n3637), .A1(n3640) );
  nand02 U1907 ( .Y(n3641), .A0(n3419), .A1(n3642) );
  nand02 U1908 ( .Y(n3643), .A0(n3638), .A1(n3644) );
  nand02 U1909 ( .Y(n3645), .A0(n3638), .A1(n3646) );
  nand02 U1910 ( .Y(n3647), .A0(n3635), .A1(n3636) );
  inv01 U1911 ( .Y(n3640), .A(n3647) );
  nand02 U1912 ( .Y(n3648), .A0(n3635), .A1(n3636) );
  inv01 U1913 ( .Y(n3642), .A(n3648) );
  nand02 U1914 ( .Y(n3649), .A0(n3635), .A1(n3637) );
  inv01 U1915 ( .Y(n3644), .A(n3649) );
  nand02 U1916 ( .Y(n3650), .A0(n3635), .A1(n3658) );
  inv01 U1917 ( .Y(n3646), .A(n3650) );
  nand02 U1918 ( .Y(n3651), .A0(n3639), .A1(n3641) );
  inv02 U1919 ( .Y(n3633), .A(n3651) );
  nand02 U1920 ( .Y(n3652), .A0(n3643), .A1(n3645) );
  inv02 U1921 ( .Y(n3634), .A(n3652) );
  nand02 U1922 ( .Y(n3843), .A0(n3653), .A1(n3654) );
  inv02 U1923 ( .Y(n3655), .A(n3878) );
  inv01 U1924 ( .Y(n3656), .A(n3825) );
  inv01 U1925 ( .Y(n3657), .A(n3824) );
  nand02 U1926 ( .Y(n3659), .A0(n3657), .A1(n3660) );
  nand02 U1927 ( .Y(n3661), .A0(n3984), .A1(n3662) );
  nand02 U1928 ( .Y(n3663), .A0(n3658), .A1(n3664) );
  nand02 U1929 ( .Y(n3665), .A0(n3658), .A1(n3666) );
  nand02 U1930 ( .Y(n3667), .A0(n3655), .A1(n3656) );
  inv01 U1931 ( .Y(n3660), .A(n3667) );
  nand02 U1932 ( .Y(n3668), .A0(n3655), .A1(n3656) );
  inv01 U1933 ( .Y(n3662), .A(n3668) );
  nand02 U1934 ( .Y(n3669), .A0(n3655), .A1(n3657) );
  inv01 U1935 ( .Y(n3664), .A(n3669) );
  nand02 U1936 ( .Y(n3670), .A0(n3655), .A1(n3984) );
  inv01 U1937 ( .Y(n3666), .A(n3670) );
  nand02 U1938 ( .Y(n3671), .A0(n3659), .A1(n3661) );
  inv02 U1939 ( .Y(n3653), .A(n3671) );
  nand02 U1940 ( .Y(n3672), .A0(n3663), .A1(n3665) );
  inv02 U1941 ( .Y(n3654), .A(n3672) );
  nand02 U1942 ( .Y(n3855), .A0(n3673), .A1(n3674) );
  inv02 U1943 ( .Y(n3675), .A(n3883) );
  inv01 U1944 ( .Y(n3676), .A(n3825) );
  inv01 U1945 ( .Y(n3677), .A(n3824) );
  nand02 U1946 ( .Y(n3678), .A0(n3677), .A1(n3679) );
  nand02 U1947 ( .Y(n3680), .A0(n2847), .A1(n3681) );
  nand02 U1948 ( .Y(n3682), .A0(n3984), .A1(n3683) );
  nand02 U1949 ( .Y(n3684), .A0(n3984), .A1(n3685) );
  nand02 U1950 ( .Y(n3686), .A0(n3675), .A1(n3676) );
  inv01 U1951 ( .Y(n3679), .A(n3686) );
  nand02 U1952 ( .Y(n3687), .A0(n3675), .A1(n3676) );
  inv01 U1953 ( .Y(n3681), .A(n3687) );
  nand02 U1954 ( .Y(n3688), .A0(n3675), .A1(n3677) );
  inv01 U1955 ( .Y(n3683), .A(n3688) );
  nand02 U1956 ( .Y(n3689), .A0(n3675), .A1(n2847) );
  inv01 U1957 ( .Y(n3685), .A(n3689) );
  nand02 U1958 ( .Y(n3690), .A0(n3678), .A1(n3680) );
  inv02 U1959 ( .Y(n3673), .A(n3690) );
  nand02 U1960 ( .Y(n3691), .A0(n3682), .A1(n3684) );
  inv02 U1961 ( .Y(n3674), .A(n3691) );
  inv02 U1962 ( .Y(n3813), .A(n3692) );
  nor02 U1963 ( .Y(n3693), .A0(n2768), .A1(n3798) );
  nor02 U1964 ( .Y(n3694), .A0(n3758), .A1(n3795) );
  inv01 U1965 ( .Y(n3695), .A(n3891) );
  nor02 U1966 ( .Y(n3692), .A0(n3695), .A1(n3696) );
  nor02 U1967 ( .Y(n3697), .A0(n3693), .A1(n3694) );
  inv01 U1968 ( .Y(n3696), .A(n3697) );
  ao22 U1969 ( .Y(n3698), .A0(n3890), .A1(n3811), .B0(n3868), .B1(n3764) );
  inv02 U1970 ( .Y(n3699), .A(n3698) );
  buf02 U1971 ( .Y(n3700), .A(n3861) );
  inv02 U1972 ( .Y(n3890), .A(n3701) );
  nor02 U1973 ( .Y(n3702), .A0(n3919), .A1(n3797) );
  nor02 U1974 ( .Y(n3703), .A0(n3921), .A1(n3795) );
  inv01 U1975 ( .Y(n3704), .A(n3922) );
  nor02 U1976 ( .Y(n3701), .A0(n3704), .A1(n3705) );
  nor02 U1977 ( .Y(n3706), .A0(n3702), .A1(n3703) );
  inv01 U1978 ( .Y(n3705), .A(n3706) );
  inv02 U1979 ( .Y(n3860), .A(n3890) );
  inv02 U1980 ( .Y(n3835), .A(n3707) );
  nor02 U1981 ( .Y(n3708), .A0(n3905), .A1(n3798) );
  nor02 U1982 ( .Y(n3709), .A0(n3756), .A1(n3795) );
  inv01 U1983 ( .Y(n3710), .A(n3908) );
  nor02 U1984 ( .Y(n3707), .A0(n3710), .A1(n3711) );
  nor02 U1985 ( .Y(n3712), .A0(n3708), .A1(n3709) );
  inv01 U1986 ( .Y(n3711), .A(n3712) );
  inv02 U1987 ( .Y(n3856), .A(n3713) );
  nor02 U1988 ( .Y(n3714), .A0(n2708), .A1(n3797) );
  nor02 U1989 ( .Y(n3715), .A0(n3312), .A1(n3795) );
  inv01 U1990 ( .Y(n3716), .A(n3912) );
  nor02 U1991 ( .Y(n3713), .A0(n3716), .A1(n3717) );
  nor02 U1992 ( .Y(n3718), .A0(n3714), .A1(n3715) );
  inv01 U1993 ( .Y(n3717), .A(n3718) );
  inv02 U1994 ( .Y(n3845), .A(n3719) );
  nor02 U1995 ( .Y(n3720), .A0(n3756), .A1(n3798) );
  nor02 U1996 ( .Y(n3721), .A0(n2708), .A1(n3795) );
  inv01 U1997 ( .Y(n3722), .A(n3910) );
  nor02 U1998 ( .Y(n3719), .A0(n3722), .A1(n3723) );
  nor02 U1999 ( .Y(n3724), .A0(n3720), .A1(n3721) );
  inv01 U2000 ( .Y(n3723), .A(n3724) );
  inv02 U2001 ( .Y(n3874), .A(n3725) );
  nor02 U2002 ( .Y(n3726), .A0(n3767), .A1(n3797) );
  nor02 U2003 ( .Y(n3727), .A0(n3915), .A1(n3795) );
  inv01 U2004 ( .Y(n3728), .A(n3916) );
  nor02 U2005 ( .Y(n3725), .A0(n3728), .A1(n3729) );
  nor02 U2006 ( .Y(n3730), .A0(n3726), .A1(n3727) );
  inv01 U2007 ( .Y(n3729), .A(n3730) );
  inv02 U2008 ( .Y(n3879), .A(n3731) );
  nor02 U2009 ( .Y(n3732), .A0(n3915), .A1(n3797) );
  nor02 U2010 ( .Y(n3733), .A0(n3309), .A1(n3795) );
  inv01 U2011 ( .Y(n3734), .A(n3917) );
  nor02 U2012 ( .Y(n3731), .A0(n3734), .A1(n3735) );
  nor02 U2013 ( .Y(n3736), .A0(n3732), .A1(n3733) );
  inv01 U2014 ( .Y(n3735), .A(n3736) );
  inv02 U2015 ( .Y(n3915), .A(opa_i[3]) );
  inv02 U2016 ( .Y(n3868), .A(n3737) );
  nor02 U2017 ( .Y(n3738), .A0(n3312), .A1(n3797) );
  nor02 U2018 ( .Y(n3739), .A0(n3767), .A1(n3795) );
  inv01 U2019 ( .Y(n3740), .A(n3914) );
  nor02 U2020 ( .Y(n3737), .A0(n3740), .A1(n3741) );
  nor02 U2021 ( .Y(n3742), .A0(n3738), .A1(n3739) );
  inv01 U2022 ( .Y(n3741), .A(n3742) );
  inv02 U2023 ( .Y(n3815), .A(n3743) );
  nor02 U2024 ( .Y(n3744), .A0(n3902), .A1(n3798) );
  nor02 U2025 ( .Y(n3745), .A0(n3905), .A1(n3795) );
  inv01 U2026 ( .Y(n3746), .A(n3906) );
  nor02 U2027 ( .Y(n3743), .A0(n3746), .A1(n3747) );
  nor02 U2028 ( .Y(n3748), .A0(n3744), .A1(n3745) );
  inv01 U2029 ( .Y(n3747), .A(n3748) );
  inv02 U2030 ( .Y(n3902), .A(opa_i[9]) );
  nand02 U2031 ( .Y(n3751), .A0(n3781), .A1(n3913) );
  nand02 U2032 ( .Y(n3750), .A0(n3781), .A1(n3913) );
  inv04 U2033 ( .Y(n3913), .A(n3778) );
  inv02 U2034 ( .Y(n3816), .A(n3749) );
  inv02 U2035 ( .Y(n3814), .A(n3751) );
  buf02 U2036 ( .Y(n3752), .A(s_sqr_zeros_o_1_) );
  buf02 U2037 ( .Y(n3753), .A(opa_i[10]) );
  inv02 U2038 ( .Y(n3754), .A(n3753) );
  buf02 U2039 ( .Y(n3755), .A(opa_i[7]) );
  inv02 U2040 ( .Y(n3756), .A(n3755) );
  buf02 U2041 ( .Y(n3757), .A(opa_i[12]) );
  inv02 U2042 ( .Y(n3758), .A(n3757) );
  inv01 U2043 ( .Y(n3760), .A(n3759) );
  inv01 U2044 ( .Y(n3762), .A(n3759) );
  inv01 U2045 ( .Y(n3761), .A(n3759) );
  inv02 U2046 ( .Y(n3897), .A(n3760) );
  or02 U2047 ( .Y(n3763), .A0(n3777), .A1(n3781) );
  inv01 U2048 ( .Y(n3764), .A(n3763) );
  inv02 U2049 ( .Y(n3765), .A(n3763) );
  buf02 U2050 ( .Y(n3766), .A(opa_i[4]) );
  inv02 U2051 ( .Y(n3767), .A(n3766) );
  buf02 U2052 ( .Y(n3768), .A(opa_i[23]) );
  ao22 U2053 ( .Y(n3770), .A0(n3911), .A1(n3777), .B0(n3885), .B1(n3913) );
  inv02 U2054 ( .Y(n3771), .A(n3770) );
  inv01 U2055 ( .Y(n3772), .A(n3770) );
  or02 U2056 ( .Y(n3773), .A0(n3992), .A1(opa_i[29]) );
  inv02 U2057 ( .Y(n3774), .A(n3773) );
  inv02 U2058 ( .Y(n3776), .A(n2706) );
  inv02 U2059 ( .Y(n3777), .A(n3776) );
  inv02 U2060 ( .Y(n3778), .A(n3776) );
  inv04 U2061 ( .Y(n3790), .A(n3789) );
  inv02 U2062 ( .Y(n3894), .A(n3780) );
  inv04 U2063 ( .Y(n3803), .A(n2921) );
  inv01 U2064 ( .Y(n3782), .A(n3980) );
  inv01 U2065 ( .Y(n3783), .A(n3919) );
  inv01 U2066 ( .Y(n3784), .A(n3921) );
  nor02 U2067 ( .Y(n3786), .A0(n3782), .A1(n3783) );
  inv02 U2068 ( .Y(n3785), .A(n3786) );
  inv02 U2069 ( .Y(n3919), .A(opa_i[1]) );
  inv04 U2070 ( .Y(n3811), .A(n3779) );
  inv04 U2071 ( .Y(n3788), .A(n3787) );
  inv04 U2072 ( .Y(n3792), .A(n3791) );
  inv02 U2073 ( .Y(n3793), .A(s_sqr_zeros_o_4_) );
  inv02 U2074 ( .Y(n3806), .A(n3794) );
  inv02 U2075 ( .Y(n3824), .A(n3795) );
  inv04 U2076 ( .Y(n3796), .A(n3866) );
  inv01 U2077 ( .Y(n3969), .A(n3331) );
  inv01 U2078 ( .Y(n3968), .A(n3924) );
  nor02 U2079 ( .Y(n3967), .A0(n3929), .A1(n3928) );
  nor02 U2080 ( .Y(n3966), .A0(n3938), .A1(n3971) );
  inv01 U2081 ( .Y(n3964), .A(n3939) );
  nor02 U2082 ( .Y(n3963), .A0(n3932), .A1(n3930) );
  inv01 U2083 ( .Y(n3962), .A(n3935) );
  and03 U2084 ( .Y(n3957), .A0(n3959), .A1(n2740), .A2(n3958) );
  inv01 U2085 ( .Y(n3959), .A(n3926) );
  nor02 U2086 ( .Y(n3958), .A0(n3924), .A1(n3331) );
  nor02 U2087 ( .Y(n3956), .A0(n3939), .A1(n3940) );
  nor02 U2088 ( .Y(n3955), .A0(n3935), .A1(n3934) );
  inv01 U2089 ( .Y(n3954), .A(n3931) );
  nand03 U2090 ( .Y(s_sqr_zeros_o_3_), .A0(n3948), .A1(n3949), .A2(n3947) );
  inv01 U2091 ( .Y(n3953), .A(n3331) );
  nor02 U2092 ( .Y(n3952), .A0(n3926), .A1(n3927) );
  inv01 U2093 ( .Y(n3951), .A(n3928) );
  nor02 U2094 ( .Y(n3950), .A0(n3930), .A1(n3931) );
  inv01 U2095 ( .Y(n3948), .A(n3933) );
  nor02 U2096 ( .Y(n3947), .A0(n3936), .A1(n3938) );
  nand03 U2097 ( .Y(s_sqr_zeros_o_4_), .A0(n2873), .A1(n3942), .A2(n3941) );
  and03 U2098 ( .Y(n3942), .A0(n3944), .A1(n3945), .A2(n3943) );
  inv01 U2099 ( .Y(n3945), .A(n3925) );
  inv01 U2100 ( .Y(n3944), .A(n3929) );
  nor02 U2101 ( .Y(n3943), .A0(n3939), .A1(n3940) );
  or02 U2102 ( .Y(n3946), .A0(n3935), .A1(n3934) );
  inv01 U2103 ( .Y(n3941), .A(n3937) );
  and02 U2105 ( .Y(s_exp_o1553_7_), .A0(s_exp_tem_8_), .A1(n3803) );
  and02 U2106 ( .Y(s_exp_o1553_6_), .A0(s_exp_tem_7_), .A1(n3803) );
  and02 U2107 ( .Y(s_exp_o1553_5_), .A0(s_exp_tem_6_), .A1(n3803) );
  and02 U2108 ( .Y(s_exp_o1553_4_), .A0(s_exp_tem_5_), .A1(n3803) );
  and02 U2109 ( .Y(s_exp_o1553_3_), .A0(s_exp_tem_4_), .A1(n3803) );
  and02 U2110 ( .Y(s_exp_o1553_2_), .A0(s_exp_tem_3_), .A1(n3803) );
  and02 U2111 ( .Y(s_exp_o1553_1_), .A0(s_exp_tem_2_), .A1(n3803) );
  and02 U2112 ( .Y(s_exp_o1553_0_), .A0(s_exp_tem_1_), .A1(n3803) );
  ao21 U2113 ( .Y(n3810), .A0(n3811), .A1(n3812), .B0(opa_i[20]) );
  ao221 U2114 ( .Y(n3809), .A0(n3813), .A1(n3814), .B0(n3815), .B1(n3816), 
        .C0(n3817) );
  ao21 U2115 ( .Y(fracta_52_o[50]), .A0(n3769), .A1(n3818), .B0(opa_i[23]) );
  inv01 U2116 ( .Y(n3820), .A(n3818) );
  nand03 U2117 ( .Y(n3818), .A0(n2719), .A1(n3821), .A2(n3310) );
  nand02 U2118 ( .Y(n3821), .A0(opa_i[22]), .A1(n3800) );
  inv01 U2119 ( .Y(n3833), .A(n3835) );
  inv01 U2120 ( .Y(n3829), .A(n3836) );
  inv01 U2121 ( .Y(n3827), .A(n3596) );
  and03 U2122 ( .Y(n3819), .A0(n2733), .A1(n3838), .A2(n3295) );
  nand02 U2123 ( .Y(n3838), .A0(opa_i[21]), .A1(n3800) );
  inv01 U2124 ( .Y(n3844), .A(n3845) );
  inv01 U2125 ( .Y(n3842), .A(n3846) );
  inv01 U2126 ( .Y(n3840), .A(n3611) );
  and03 U2127 ( .Y(n3837), .A0(n3848), .A1(n3849), .A2(n3313) );
  nand02 U2128 ( .Y(n3849), .A0(n3800), .A1(opa_i[20]) );
  inv01 U2129 ( .Y(n3853), .A(n3856) );
  nor02 U2130 ( .Y(n3851), .A0(n3781), .A1(n3772) );
  inv01 U2131 ( .Y(n3862), .A(n3812) );
  ao22 U2132 ( .Y(n3873), .A0(n3799), .A1(opa_i[17]), .B0(n3800), .B1(
        opa_i[18]) );
  ao22 U2133 ( .Y(n3878), .A0(n3799), .A1(opa_i[16]), .B0(n3800), .B1(
        opa_i[17]) );
  inv01 U2134 ( .Y(n3875), .A(n3880) );
  ao22 U2135 ( .Y(n3883), .A0(n3799), .A1(opa_i[15]), .B0(n3800), .B1(
        opa_i[16]) );
  nand02 U2136 ( .Y(n3861), .A0(n3765), .A1(n3794) );
  ao22 U2137 ( .Y(n3889), .A0(n3790), .A1(n3813), .B0(n3117), .B1(n3890) );
  ao22 U2138 ( .Y(n3893), .A0(n3790), .A1(n3836), .B0(n3117), .B1(n3894) );
  ao22 U2139 ( .Y(n3896), .A0(n3117), .A1(n3897), .B0(n3790), .B1(n3846) );
  nand02 U2140 ( .Y(n3834), .A0(n3781), .A1(n3777) );
  nor02 U2141 ( .Y(n3887), .A0(n3794), .A1(n3779) );
  nor02 U2142 ( .Y(n3888), .A0(n3794), .A1(n3830) );
  nand02 U2143 ( .Y(n3830), .A0(n3781), .A1(n3913) );
  nand02 U2144 ( .Y(n3832), .A0(n3778), .A1(n3901) );
  inv01 U2145 ( .Y(n3901), .A(n3781) );
  nand02 U2146 ( .Y(n3808), .A0(n3769), .A1(n3806) );
  inv01 U2147 ( .Y(n3911), .A(n3613) );
  nand02 U2148 ( .Y(n3864), .A0(n3752), .A1(n3614) );
  nand02 U2149 ( .Y(n3866), .A0(n3752), .A1(n3923) );
  nand02 U2150 ( .Y(n3918), .A0(n3790), .A1(n3801) );
  nand02 U2151 ( .Y(n3863), .A0(n3765), .A1(n3806) );
  and04 U2152 ( .Y(n3949), .A0(n3950), .A1(n3951), .A2(n3952), .A3(n3953) );
  nand04 U2153 ( .Y(s_sqr_zeros_o_2_), .A0(n3954), .A1(n3955), .A2(n3956), 
        .A3(n3957) );
  nor02 U2154 ( .Y(n3823), .A0(n3923), .A1(n3752) );
  inv01 U2155 ( .Y(n3923), .A(n3614) );
  nand02 U2156 ( .Y(n3882), .A0(n3800), .A1(opa_i[0]) );
  nor02 U2157 ( .Y(n3826), .A0(n3614), .A1(n3752) );
  nand04 U2158 ( .Y(s_sqr_zeros_o_1_), .A0(n3962), .A1(n3963), .A2(n3964), 
        .A3(n3965) );
  and04 U2159 ( .Y(n3965), .A0(n3966), .A1(n3967), .A2(n3968), .A3(n3969) );
  and03 U2160 ( .Y(n3934), .A0(n3002), .A1(n3767), .A2(opa_i[3]) );
  inv01 U2161 ( .Y(n3929), .A(n3970) );
  inv01 U2162 ( .Y(n3865), .A(opa_i[17]) );
  and02 U2163 ( .Y(n3937), .A0(opa_i[7]), .A1(n3054) );
  nor02 U2164 ( .Y(n3936), .A0(n3658), .A1(n3974) );
  inv01 U2165 ( .Y(n3940), .A(n3976) );
  inv01 U2166 ( .Y(n3939), .A(n3977) );
  and03 U2167 ( .Y(n3931), .A0(n2742), .A1(n3758), .A2(opa_i[11]) );
  and02 U2168 ( .Y(n3930), .A0(opa_i[13]), .A1(n3978) );
  and02 U2169 ( .Y(n3932), .A0(opa_i[5]), .A1(n3979) );
  and02 U2170 ( .Y(n3935), .A0(opa_i[1]), .A1(n3980) );
  inv01 U2171 ( .Y(n3933), .A(n3803) );
  inv01 U2172 ( .Y(n3921), .A(opa_i[0]) );
  nand02 U2173 ( .Y(s_sqr_zeros_o_0_), .A0(n3981), .A1(n3982) );
  and02 U2174 ( .Y(n3928), .A0(opa_i[12]), .A1(n2742) );
  and02 U2175 ( .Y(n3926), .A0(opa_i[10]), .A1(n3975) );
  nand03 U2176 ( .Y(n3983), .A0(n3976), .A1(n3977), .A2(n3944) );
  nand02 U2177 ( .Y(n3970), .A0(opa_i[4]), .A1(n3002) );
  nand02 U2178 ( .Y(n3976), .A0(opa_i[2]), .A1(n3985) );
  and02 U2179 ( .Y(n3980), .A0(n3985), .A1(n3309) );
  and03 U2180 ( .Y(n3985), .A0(n3915), .A1(n3767), .A2(n3002) );
  and03 U2181 ( .Y(n3979), .A0(n2708), .A1(n3756), .A2(n3054) );
  and02 U2182 ( .Y(n3924), .A0(opa_i[16]), .A1(n2717) );
  and03 U2183 ( .Y(n3925), .A0(n3054), .A1(n3756), .A2(opa_i[6]) );
  and03 U2184 ( .Y(n3987), .A0(n3754), .A1(n3902), .A2(n3975) );
  nand02 U2185 ( .Y(n3974), .A0(n2717), .A1(n3638) );
  or03 U2186 ( .Y(n3961), .A0(opa_i[18]), .A1(opa_i[19]), .A2(opa_i[17]) );
  inv01 U2187 ( .Y(n3989), .A(opa_i[21]) );
  nand02 U2188 ( .Y(n3817), .A0(n3774), .A1(n2988) );
  inv01 U2189 ( .Y(n3990), .A(n3101) );
  nor02 U2190 ( .Y(n3973), .A0(opa_i[21]), .A1(opa_i[20]) );
  nor02 U2191 ( .Y(n____return1466_8_), .A0(n3774), .A1(n2988) );
  inv01 U2192 ( .Y(n3991), .A(opa_i[30]) );
  ao21 U2193 ( .Y(n____return1466_6_), .A0(opa_i[29]), .A1(n3992), .B0(n3774)
         );
  inv01 U2194 ( .Y(n3992), .A(n3111) );
  inv01 U2195 ( .Y(n3993), .A(n3289) );
  inv01 U2196 ( .Y(n3804), .A(n3107) );
  inv01 U2197 ( .Y(n3994), .A(n3109) );
  inv01 U2198 ( .Y(n3995), .A(n3347) );
  inv01 U2199 ( .Y(n____return1466_0_), .A(opa_i[23]) );
  pre_norm_sqrt_DW01_sub_9_0 sub_0_root_sub_92_minus_minus ( .A({n2790, n3358, 
        n3015, n____return1466_5_, n1468_4_, n____return1466_3_, 
        n____return1466_2_, n____return1466_1_, n3801}), .B({1'b0, 1'b0, 1'b0, 
        1'b0, n3794, n3781, n3778, n3752, n3614}), .CI(1'b0), .DIFF({
        s_exp_tem_8_, s_exp_tem_7_, s_exp_tem_6_, s_exp_tem_5_, s_exp_tem_4_, 
        s_exp_tem_3_, s_exp_tem_2_, s_exp_tem_1_, SYNOPSYS_UNCONNECTED_1}) );
endmodule


module post_norm_sqrt_DW01_inc_23_0 ( A, SUM );
  input [22:0] A;
  output [22:0] SUM;
  wire   carry_22_, carry_21_, carry_20_, carry_19_, carry_18_, carry_17_,
         carry_16_, carry_15_, carry_14_, carry_13_, carry_12_, carry_11_,
         carry_10_, carry_9_, carry_8_, carry_7_, carry_6_, carry_5_, carry_4_,
         carry_3_, carry_2_;

  inv04 U5 ( .Y(SUM[0]), .A(A[0]) );
  xor2 U6 ( .Y(SUM[22]), .A0(carry_22_), .A1(A[22]) );
  hadd1 U1_1_1 ( .S(SUM[1]), .CO(carry_2_), .A(A[1]), .B(A[0]) );
  hadd1 U1_1_2 ( .S(SUM[2]), .CO(carry_3_), .A(A[2]), .B(carry_2_) );
  hadd1 U1_1_3 ( .S(SUM[3]), .CO(carry_4_), .A(A[3]), .B(carry_3_) );
  hadd1 U1_1_4 ( .S(SUM[4]), .CO(carry_5_), .A(A[4]), .B(carry_4_) );
  hadd1 U1_1_5 ( .S(SUM[5]), .CO(carry_6_), .A(A[5]), .B(carry_5_) );
  hadd1 U1_1_6 ( .S(SUM[6]), .CO(carry_7_), .A(A[6]), .B(carry_6_) );
  hadd1 U1_1_7 ( .S(SUM[7]), .CO(carry_8_), .A(A[7]), .B(carry_7_) );
  hadd1 U1_1_8 ( .S(SUM[8]), .CO(carry_9_), .A(A[8]), .B(carry_8_) );
  hadd1 U1_1_9 ( .S(SUM[9]), .CO(carry_10_), .A(A[9]), .B(carry_9_) );
  hadd1 U1_1_10 ( .S(SUM[10]), .CO(carry_11_), .A(A[10]), .B(carry_10_) );
  hadd1 U1_1_11 ( .S(SUM[11]), .CO(carry_12_), .A(A[11]), .B(carry_11_) );
  hadd1 U1_1_12 ( .S(SUM[12]), .CO(carry_13_), .A(A[12]), .B(carry_12_) );
  hadd1 U1_1_13 ( .S(SUM[13]), .CO(carry_14_), .A(A[13]), .B(carry_13_) );
  hadd1 U1_1_14 ( .S(SUM[14]), .CO(carry_15_), .A(A[14]), .B(carry_14_) );
  hadd1 U1_1_15 ( .S(SUM[15]), .CO(carry_16_), .A(A[15]), .B(carry_15_) );
  hadd1 U1_1_16 ( .S(SUM[16]), .CO(carry_17_), .A(A[16]), .B(carry_16_) );
  hadd1 U1_1_17 ( .S(SUM[17]), .CO(carry_18_), .A(A[17]), .B(carry_17_) );
  hadd1 U1_1_18 ( .S(SUM[18]), .CO(carry_19_), .A(A[18]), .B(carry_18_) );
  hadd1 U1_1_19 ( .S(SUM[19]), .CO(carry_20_), .A(A[19]), .B(carry_19_) );
  hadd1 U1_1_20 ( .S(SUM[20]), .CO(carry_21_), .A(A[20]), .B(carry_20_) );
  hadd1 U1_1_21 ( .S(SUM[21]), .CO(carry_22_), .A(A[21]), .B(carry_21_) );
endmodule


module post_norm_sqrt ( clk_i, opa_i, fract_26_i, exp_i, ine_i, rmode_i, 
        output_o, ine_o );
  input [31:0] opa_i;
  input [25:0] fract_26_i;
  input [7:0] exp_i;
  input [1:0] rmode_i;
  output [31:0] output_o;
  input clk_i, ine_i;
  output ine_o;
  wire   s_output_o_30_, s_output_o_29_, s_output_o_28_, s_output_o_27_,
         s_output_o_26_, s_output_o_25_, s_output_o_24_, s_output_o_23_,
         s_output_o_22_, s_ine_o, s_fraco1_24_, s_fraco1_23_, s_fraco1_22_,
         s_fraco1_21_, s_fraco1_20_, s_fraco1_19_, s_fraco1_18_, s_fraco1_17_,
         s_fraco1_16_, s_fraco1_15_, s_fraco1_14_, s_fraco1_13_, s_fraco1_12_,
         s_fraco1_11_, s_fraco1_10_, s_fraco1_9_, s_fraco1_8_, s_fraco1_7_,
         s_fraco1_6_, s_fraco1_5_, s_fraco1_4_, s_fraco1_3_, s_fraco1_2_,
         s_guard, s_round, s_sticky, s_sign_i, s_frac_rnd_22_, s_opa_i_28_,
         s_opa_i_27_, s_opa_i_26_, s_opa_i_25_, s_opa_i_24_, s_opa_i_23_,
         s_opa_i_21_, s_opa_i_20_, s_opa_i_16_, s_opa_i_15_, s_opa_i_14_,
         s_opa_i_11_, s_opa_i_10_, s_opa_i_6_, s_opa_i_5_, s_opa_i_4_,
         s_opa_i_1_, s_opa_i_0_, s_rmode_i_1_, s_rmode_i_0_, s_frac_rnd254_22_,
         s_frac_rnd254_21_, s_frac_rnd254_20_, s_frac_rnd254_19_,
         s_frac_rnd254_18_, s_frac_rnd254_17_, s_frac_rnd254_16_,
         s_frac_rnd254_15_, s_frac_rnd254_14_, s_frac_rnd254_13_,
         s_frac_rnd254_12_, s_frac_rnd254_11_, s_frac_rnd254_10_,
         s_frac_rnd254_9_, s_frac_rnd254_8_, s_frac_rnd254_7_,
         s_frac_rnd254_6_, s_frac_rnd254_5_, s_frac_rnd254_4_,
         s_frac_rnd254_3_, s_frac_rnd254_2_, s_frac_rnd254_1_,
         s_frac_rnd254_0_, n283_22_, n____return281_21_, n____return281_20_,
         n____return281_19_, n____return281_18_, n____return281_17_,
         n____return281_16_, n____return281_15_, n____return281_14_,
         n____return281_13_, n____return281_12_, n____return281_11_,
         n____return281_10_, n____return281_9_, n____return281_8_,
         n____return281_7_, n____return281_6_, n____return281_5_,
         n____return281_4_, n____return281_3_, n____return281_2_,
         n____return281_1_, n____return281_0_, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908;

  dff s_expa_reg_7_ ( .QB(n869), .D(opa_i[30]), .CLK(clk_i) );
  dff s_expa_reg_6_ ( .QB(n868), .D(opa_i[29]), .CLK(clk_i) );
  dff s_expa_reg_5_ ( .QB(n867), .D(opa_i[28]), .CLK(clk_i) );
  dff s_expa_reg_4_ ( .QB(n866), .D(opa_i[27]), .CLK(clk_i) );
  dff s_expa_reg_3_ ( .QB(n873), .D(opa_i[26]), .CLK(clk_i) );
  dff s_expa_reg_2_ ( .QB(n872), .D(opa_i[25]), .CLK(clk_i) );
  dff s_expa_reg_1_ ( .QB(n871), .D(opa_i[24]), .CLK(clk_i) );
  dff s_expa_reg_0_ ( .QB(n870), .D(opa_i[23]), .CLK(clk_i) );
  dff s_fract_26_i_reg_24_ ( .Q(s_fraco1_24_), .QB(n895), .D(fract_26_i[24]), 
        .CLK(clk_i) );
  dff s_fract_26_i_reg_23_ ( .Q(s_fraco1_23_), .QB(n896), .D(fract_26_i[23]), 
        .CLK(clk_i) );
  dff s_fract_26_i_reg_22_ ( .Q(s_fraco1_22_), .QB(n897), .D(fract_26_i[22]), 
        .CLK(clk_i) );
  dff s_fract_26_i_reg_21_ ( .Q(s_fraco1_21_), .QB(n898), .D(fract_26_i[21]), 
        .CLK(clk_i) );
  dff s_fract_26_i_reg_20_ ( .Q(s_fraco1_20_), .QB(n899), .D(fract_26_i[20]), 
        .CLK(clk_i) );
  dff s_fract_26_i_reg_19_ ( .Q(s_fraco1_19_), .QB(n900), .D(fract_26_i[19]), 
        .CLK(clk_i) );
  dff s_fract_26_i_reg_18_ ( .Q(s_fraco1_18_), .QB(n901), .D(fract_26_i[18]), 
        .CLK(clk_i) );
  dff s_fract_26_i_reg_17_ ( .Q(s_fraco1_17_), .QB(n902), .D(fract_26_i[17]), 
        .CLK(clk_i) );
  dff s_fract_26_i_reg_16_ ( .Q(s_fraco1_16_), .QB(n903), .D(fract_26_i[16]), 
        .CLK(clk_i) );
  dff s_fract_26_i_reg_15_ ( .Q(s_fraco1_15_), .QB(n904), .D(fract_26_i[15]), 
        .CLK(clk_i) );
  dff s_fract_26_i_reg_14_ ( .Q(s_fraco1_14_), .QB(n905), .D(fract_26_i[14]), 
        .CLK(clk_i) );
  dff s_fract_26_i_reg_13_ ( .Q(s_fraco1_13_), .QB(n906), .D(fract_26_i[13]), 
        .CLK(clk_i) );
  dff s_fract_26_i_reg_12_ ( .Q(s_fraco1_12_), .QB(n907), .D(fract_26_i[12]), 
        .CLK(clk_i) );
  dff s_fract_26_i_reg_11_ ( .Q(s_fraco1_11_), .QB(n887), .D(fract_26_i[11]), 
        .CLK(clk_i) );
  dff s_fract_26_i_reg_10_ ( .Q(s_fraco1_10_), .QB(n888), .D(fract_26_i[10]), 
        .CLK(clk_i) );
  dff s_fract_26_i_reg_9_ ( .Q(s_fraco1_9_), .QB(n889), .D(fract_26_i[9]), 
        .CLK(clk_i) );
  dff s_fract_26_i_reg_8_ ( .Q(s_fraco1_8_), .QB(n890), .D(fract_26_i[8]), 
        .CLK(clk_i) );
  dff s_fract_26_i_reg_7_ ( .Q(s_fraco1_7_), .QB(n891), .D(fract_26_i[7]), 
        .CLK(clk_i) );
  dff s_fract_26_i_reg_6_ ( .Q(s_fraco1_6_), .QB(n892), .D(fract_26_i[6]), 
        .CLK(clk_i) );
  dff s_fract_26_i_reg_5_ ( .Q(s_fraco1_5_), .QB(n893), .D(fract_26_i[5]), 
        .CLK(clk_i) );
  dff s_fract_26_i_reg_4_ ( .Q(s_fraco1_4_), .QB(n894), .D(fract_26_i[4]), 
        .CLK(clk_i) );
  dff s_fract_26_i_reg_3_ ( .Q(s_fraco1_3_), .D(fract_26_i[3]), .CLK(clk_i) );
  dff s_fract_26_i_reg_2_ ( .Q(s_fraco1_2_), .QB(n908), .D(fract_26_i[2]), 
        .CLK(clk_i) );
  dff s_fract_26_i_reg_1_ ( .Q(s_guard), .D(fract_26_i[1]), .CLK(clk_i) );
  dff s_fract_26_i_reg_0_ ( .Q(s_round), .D(fract_26_i[0]), .CLK(clk_i) );
  dff s_exp_i_reg_7_ ( .QB(n843), .D(exp_i[7]), .CLK(clk_i) );
  dff s_exp_i_reg_6_ ( .QB(n845), .D(exp_i[6]), .CLK(clk_i) );
  dff s_exp_i_reg_5_ ( .QB(n846), .D(exp_i[5]), .CLK(clk_i) );
  dff s_exp_i_reg_4_ ( .QB(n847), .D(exp_i[4]), .CLK(clk_i) );
  dff s_exp_i_reg_3_ ( .QB(n848), .D(exp_i[3]), .CLK(clk_i) );
  dff s_exp_i_reg_2_ ( .QB(n849), .D(exp_i[2]), .CLK(clk_i) );
  dff s_exp_i_reg_1_ ( .QB(n850), .D(exp_i[1]), .CLK(clk_i) );
  dff s_exp_i_reg_0_ ( .QB(n851), .D(exp_i[0]), .CLK(clk_i) );
  dff s_rmode_i_reg_1_ ( .Q(s_rmode_i_1_), .D(rmode_i[1]), .CLK(clk_i) );
  dff s_rmode_i_reg_0_ ( .Q(s_rmode_i_0_), .D(rmode_i[0]), .CLK(clk_i) );
  dff output_o_reg_31_ ( .Q(output_o[31]), .D(s_sign_i), .CLK(clk_i) );
  dff output_o_reg_30_ ( .Q(output_o[30]), .D(s_output_o_30_), .CLK(clk_i) );
  dff output_o_reg_29_ ( .Q(output_o[29]), .D(s_output_o_29_), .CLK(clk_i) );
  dff output_o_reg_28_ ( .Q(output_o[28]), .D(s_output_o_28_), .CLK(clk_i) );
  dff output_o_reg_27_ ( .Q(output_o[27]), .D(s_output_o_27_), .CLK(clk_i) );
  dff output_o_reg_26_ ( .Q(output_o[26]), .D(s_output_o_26_), .CLK(clk_i) );
  dff output_o_reg_25_ ( .Q(output_o[25]), .D(s_output_o_25_), .CLK(clk_i) );
  dff output_o_reg_24_ ( .Q(output_o[24]), .D(s_output_o_24_), .CLK(clk_i) );
  dff output_o_reg_23_ ( .Q(output_o[23]), .D(s_output_o_23_), .CLK(clk_i) );
  dff output_o_reg_22_ ( .Q(output_o[22]), .D(s_output_o_22_), .CLK(clk_i) );
  dff output_o_reg_21_ ( .Q(output_o[21]), .D(n689), .CLK(clk_i) );
  dff output_o_reg_20_ ( .Q(output_o[20]), .D(n697), .CLK(clk_i) );
  dff output_o_reg_19_ ( .Q(output_o[19]), .D(n677), .CLK(clk_i) );
  dff output_o_reg_18_ ( .Q(output_o[18]), .D(n679), .CLK(clk_i) );
  dff output_o_reg_17_ ( .Q(output_o[17]), .D(n663), .CLK(clk_i) );
  dff output_o_reg_16_ ( .Q(output_o[16]), .D(n693), .CLK(clk_i) );
  dff output_o_reg_15_ ( .Q(output_o[15]), .D(n683), .CLK(clk_i) );
  dff output_o_reg_14_ ( .Q(output_o[14]), .D(n673), .CLK(clk_i) );
  dff output_o_reg_13_ ( .Q(output_o[13]), .D(n699), .CLK(clk_i) );
  dff output_o_reg_12_ ( .Q(output_o[12]), .D(n691), .CLK(clk_i) );
  dff output_o_reg_11_ ( .Q(output_o[11]), .D(n681), .CLK(clk_i) );
  dff output_o_reg_10_ ( .Q(output_o[10]), .D(n667), .CLK(clk_i) );
  dff output_o_reg_9_ ( .Q(output_o[9]), .D(n705), .CLK(clk_i) );
  dff output_o_reg_8_ ( .Q(output_o[8]), .D(n669), .CLK(clk_i) );
  dff output_o_reg_7_ ( .Q(output_o[7]), .D(n675), .CLK(clk_i) );
  dff output_o_reg_6_ ( .Q(output_o[6]), .D(n687), .CLK(clk_i) );
  dff output_o_reg_5_ ( .Q(output_o[5]), .D(n703), .CLK(clk_i) );
  dff output_o_reg_4_ ( .Q(output_o[4]), .D(n665), .CLK(clk_i) );
  dff output_o_reg_3_ ( .Q(output_o[3]), .D(n685), .CLK(clk_i) );
  dff output_o_reg_2_ ( .Q(output_o[2]), .D(n701), .CLK(clk_i) );
  dff output_o_reg_1_ ( .Q(output_o[1]), .D(n695), .CLK(clk_i) );
  dff output_o_reg_0_ ( .Q(output_o[0]), .D(n671), .CLK(clk_i) );
  dff s_opa_i_reg_30_ ( .QB(n886), .D(opa_i[30]), .CLK(clk_i) );
  dff s_opa_i_reg_29_ ( .QB(n885), .D(opa_i[29]), .CLK(clk_i) );
  dff s_opa_i_reg_28_ ( .Q(s_opa_i_28_), .D(opa_i[28]), .CLK(clk_i) );
  dff s_opa_i_reg_27_ ( .Q(s_opa_i_27_), .D(opa_i[27]), .CLK(clk_i) );
  dff s_opa_i_reg_26_ ( .Q(s_opa_i_26_), .D(opa_i[26]), .CLK(clk_i) );
  dff s_opa_i_reg_25_ ( .Q(s_opa_i_25_), .D(opa_i[25]), .CLK(clk_i) );
  dff s_opa_i_reg_24_ ( .Q(s_opa_i_24_), .D(opa_i[24]), .CLK(clk_i) );
  dff s_opa_i_reg_23_ ( .Q(s_opa_i_23_), .D(opa_i[23]), .CLK(clk_i) );
  dff s_opa_i_reg_22_ ( .QB(n877), .D(opa_i[22]), .CLK(clk_i) );
  dff s_opa_i_reg_21_ ( .Q(s_opa_i_21_), .D(opa_i[21]), .CLK(clk_i) );
  dff s_opa_i_reg_20_ ( .Q(s_opa_i_20_), .D(opa_i[20]), .CLK(clk_i) );
  dff s_opa_i_reg_19_ ( .QB(n882), .D(opa_i[19]), .CLK(clk_i) );
  dff s_opa_i_reg_18_ ( .QB(n881), .D(opa_i[18]), .CLK(clk_i) );
  dff s_opa_i_reg_17_ ( .QB(n880), .D(opa_i[17]), .CLK(clk_i) );
  dff s_opa_i_reg_16_ ( .Q(s_opa_i_16_), .D(opa_i[16]), .CLK(clk_i) );
  dff s_opa_i_reg_15_ ( .Q(s_opa_i_15_), .D(opa_i[15]), .CLK(clk_i) );
  dff s_opa_i_reg_14_ ( .Q(s_opa_i_14_), .D(opa_i[14]), .CLK(clk_i) );
  dff s_opa_i_reg_13_ ( .QB(n884), .D(opa_i[13]), .CLK(clk_i) );
  dff s_opa_i_reg_12_ ( .QB(n883), .D(opa_i[12]), .CLK(clk_i) );
  dff s_opa_i_reg_11_ ( .Q(s_opa_i_11_), .D(opa_i[11]), .CLK(clk_i) );
  dff s_opa_i_reg_10_ ( .Q(s_opa_i_10_), .D(opa_i[10]), .CLK(clk_i) );
  dff s_opa_i_reg_9_ ( .QB(n876), .D(opa_i[9]), .CLK(clk_i) );
  dff s_opa_i_reg_8_ ( .QB(n875), .D(opa_i[8]), .CLK(clk_i) );
  dff s_opa_i_reg_7_ ( .QB(n874), .D(opa_i[7]), .CLK(clk_i) );
  dff s_opa_i_reg_6_ ( .Q(s_opa_i_6_), .D(opa_i[6]), .CLK(clk_i) );
  dff s_opa_i_reg_5_ ( .Q(s_opa_i_5_), .D(opa_i[5]), .CLK(clk_i) );
  dff s_opa_i_reg_4_ ( .Q(s_opa_i_4_), .D(opa_i[4]), .CLK(clk_i) );
  dff s_opa_i_reg_3_ ( .QB(n879), .D(opa_i[3]), .CLK(clk_i) );
  dff s_opa_i_reg_2_ ( .QB(n878), .D(opa_i[2]), .CLK(clk_i) );
  dff s_opa_i_reg_1_ ( .Q(s_opa_i_1_), .D(opa_i[1]), .CLK(clk_i) );
  dff s_opa_i_reg_0_ ( .Q(s_opa_i_0_), .D(opa_i[0]), .CLK(clk_i) );
  dff s_sign_i_reg ( .Q(s_sign_i), .D(opa_i[31]), .CLK(clk_i) );
  dff s_ine_i_reg ( .Q(s_sticky), .D(ine_i), .CLK(clk_i) );
  dff ine_o_reg ( .Q(ine_o), .D(s_ine_o), .CLK(clk_i) );
  dff s_frac_rnd_reg_22_ ( .Q(s_frac_rnd_22_), .D(n722), .CLK(clk_i) );
  dff s_frac_rnd_reg_21_ ( .QB(n852), .D(n720), .CLK(clk_i) );
  dff s_frac_rnd_reg_20_ ( .QB(n853), .D(n728), .CLK(clk_i) );
  dff s_frac_rnd_reg_19_ ( .QB(n855), .D(n721), .CLK(clk_i) );
  dff s_frac_rnd_reg_18_ ( .QB(n856), .D(s_frac_rnd254_18_), .CLK(clk_i) );
  dff s_frac_rnd_reg_17_ ( .QB(n857), .D(n709), .CLK(clk_i) );
  dff s_frac_rnd_reg_16_ ( .QB(n858), .D(n725), .CLK(clk_i) );
  dff s_frac_rnd_reg_15_ ( .QB(n859), .D(n726), .CLK(clk_i) );
  dff s_frac_rnd_reg_14_ ( .QB(n860), .D(n723), .CLK(clk_i) );
  dff s_frac_rnd_reg_13_ ( .QB(n861), .D(n729), .CLK(clk_i) );
  dff s_frac_rnd_reg_12_ ( .QB(n862), .D(n715), .CLK(clk_i) );
  dff s_frac_rnd_reg_11_ ( .QB(n863), .D(n713), .CLK(clk_i) );
  dff s_frac_rnd_reg_10_ ( .QB(n864), .D(n710), .CLK(clk_i) );
  dff s_frac_rnd_reg_9_ ( .QB(n836), .D(n712), .CLK(clk_i) );
  dff s_frac_rnd_reg_8_ ( .QB(n837), .D(n717), .CLK(clk_i) );
  dff s_frac_rnd_reg_7_ ( .QB(n838), .D(n718), .CLK(clk_i) );
  dff s_frac_rnd_reg_6_ ( .QB(n839), .D(n719), .CLK(clk_i) );
  dff s_frac_rnd_reg_5_ ( .QB(n840), .D(n724), .CLK(clk_i) );
  dff s_frac_rnd_reg_4_ ( .QB(n841), .D(n711), .CLK(clk_i) );
  dff s_frac_rnd_reg_3_ ( .QB(n842), .D(n727), .CLK(clk_i) );
  dff s_frac_rnd_reg_2_ ( .QB(n844), .D(n714), .CLK(clk_i) );
  dff s_frac_rnd_reg_1_ ( .QB(n854), .D(s_frac_rnd254_1_), .CLK(clk_i) );
  dff s_frac_rnd_reg_0_ ( .QB(n865), .D(n716), .CLK(clk_i) );
  xor2 U295 ( .Y(n660), .A0(s_sign_i), .A1(s_rmode_i_0_) );
  inv01 U296 ( .Y(n661), .A(n660) );
  or02 U297 ( .Y(n662), .A0(n793), .A1(n857) );
  inv01 U298 ( .Y(n663), .A(n662) );
  or02 U299 ( .Y(n664), .A0(n793), .A1(n841) );
  inv01 U300 ( .Y(n665), .A(n664) );
  or02 U301 ( .Y(n666), .A0(n793), .A1(n864) );
  inv01 U302 ( .Y(n667), .A(n666) );
  or02 U303 ( .Y(n668), .A0(n793), .A1(n837) );
  inv01 U304 ( .Y(n669), .A(n668) );
  or02 U305 ( .Y(n670), .A0(n793), .A1(n865) );
  inv01 U306 ( .Y(n671), .A(n670) );
  or02 U307 ( .Y(n672), .A0(n793), .A1(n860) );
  inv01 U308 ( .Y(n673), .A(n672) );
  or02 U309 ( .Y(n674), .A0(n793), .A1(n838) );
  inv01 U310 ( .Y(n675), .A(n674) );
  or02 U311 ( .Y(n676), .A0(n793), .A1(n855) );
  inv01 U312 ( .Y(n677), .A(n676) );
  or02 U313 ( .Y(n678), .A0(n793), .A1(n856) );
  inv01 U314 ( .Y(n679), .A(n678) );
  or02 U315 ( .Y(n680), .A0(n793), .A1(n863) );
  inv01 U316 ( .Y(n681), .A(n680) );
  or02 U317 ( .Y(n682), .A0(n793), .A1(n859) );
  inv01 U318 ( .Y(n683), .A(n682) );
  or02 U319 ( .Y(n684), .A0(n793), .A1(n842) );
  inv01 U320 ( .Y(n685), .A(n684) );
  or02 U321 ( .Y(n686), .A0(n793), .A1(n839) );
  inv01 U322 ( .Y(n687), .A(n686) );
  or02 U323 ( .Y(n688), .A0(n793), .A1(n852) );
  inv01 U324 ( .Y(n689), .A(n688) );
  or02 U325 ( .Y(n690), .A0(n793), .A1(n862) );
  inv01 U326 ( .Y(n691), .A(n690) );
  or02 U327 ( .Y(n692), .A0(n793), .A1(n858) );
  inv01 U328 ( .Y(n693), .A(n692) );
  or02 U329 ( .Y(n694), .A0(n793), .A1(n854) );
  inv01 U330 ( .Y(n695), .A(n694) );
  or02 U331 ( .Y(n696), .A0(n793), .A1(n853) );
  inv01 U332 ( .Y(n697), .A(n696) );
  or02 U333 ( .Y(n698), .A0(n793), .A1(n861) );
  inv01 U334 ( .Y(n699), .A(n698) );
  or02 U335 ( .Y(n700), .A0(n793), .A1(n844) );
  inv01 U336 ( .Y(n701), .A(n700) );
  or02 U337 ( .Y(n702), .A0(n793), .A1(n840) );
  inv01 U338 ( .Y(n703), .A(n702) );
  or02 U339 ( .Y(n704), .A0(n793), .A1(n836) );
  inv01 U340 ( .Y(n705), .A(n704) );
  inv01 U341 ( .Y(n833), .A(n706) );
  nor02 U342 ( .Y(n707), .A0(s_round), .A1(s_sticky) );
  inv01 U343 ( .Y(n708), .A(n834) );
  nor02 U344 ( .Y(n706), .A0(n707), .A1(n708) );
  buf02 U345 ( .Y(n709), .A(s_frac_rnd254_17_) );
  buf02 U346 ( .Y(n710), .A(s_frac_rnd254_10_) );
  buf02 U347 ( .Y(n711), .A(s_frac_rnd254_4_) );
  buf02 U348 ( .Y(n712), .A(s_frac_rnd254_9_) );
  buf02 U349 ( .Y(n713), .A(s_frac_rnd254_11_) );
  buf02 U350 ( .Y(n714), .A(s_frac_rnd254_2_) );
  buf02 U351 ( .Y(n715), .A(s_frac_rnd254_12_) );
  buf02 U352 ( .Y(n716), .A(s_frac_rnd254_0_) );
  buf02 U353 ( .Y(n717), .A(s_frac_rnd254_8_) );
  buf02 U354 ( .Y(n718), .A(s_frac_rnd254_7_) );
  buf02 U355 ( .Y(n719), .A(s_frac_rnd254_6_) );
  buf02 U356 ( .Y(n720), .A(s_frac_rnd254_21_) );
  buf02 U357 ( .Y(n721), .A(s_frac_rnd254_19_) );
  buf02 U358 ( .Y(n722), .A(s_frac_rnd254_22_) );
  buf02 U359 ( .Y(n723), .A(s_frac_rnd254_14_) );
  buf02 U360 ( .Y(n724), .A(s_frac_rnd254_5_) );
  buf02 U361 ( .Y(n725), .A(s_frac_rnd254_16_) );
  buf02 U362 ( .Y(n726), .A(s_frac_rnd254_15_) );
  buf02 U363 ( .Y(n727), .A(s_frac_rnd254_3_) );
  buf02 U364 ( .Y(n728), .A(s_frac_rnd254_20_) );
  buf02 U365 ( .Y(n729), .A(s_frac_rnd254_13_) );
  nand02 U366 ( .Y(s_frac_rnd254_18_), .A0(n730), .A1(n731) );
  inv01 U367 ( .Y(n732), .A(n899) );
  inv01 U368 ( .Y(n733), .A(n822) );
  inv01 U369 ( .Y(n734), .A(n794) );
  nand02 U370 ( .Y(n730), .A0(n794), .A1(n732) );
  nand02 U371 ( .Y(n731), .A0(n733), .A1(n734) );
  inv01 U372 ( .Y(n735), .A(n739) );
  or04 U373 ( .Y(n736), .A0(n866), .A1(n867), .A2(n868), .A3(n869) );
  inv01 U374 ( .Y(n737), .A(n736) );
  inv01 U375 ( .Y(n801), .A(n738) );
  inv01 U376 ( .Y(n739), .A(n799) );
  inv01 U377 ( .Y(n740), .A(s_opa_i_23_) );
  inv01 U378 ( .Y(n741), .A(s_opa_i_24_) );
  inv01 U379 ( .Y(n742), .A(s_opa_i_25_) );
  nand02 U380 ( .Y(n738), .A0(n743), .A1(n744) );
  nand02 U381 ( .Y(n745), .A0(n739), .A1(n740) );
  inv01 U382 ( .Y(n743), .A(n745) );
  nand02 U383 ( .Y(n746), .A0(n741), .A1(n742) );
  inv01 U384 ( .Y(n744), .A(n746) );
  or04 U385 ( .Y(n747), .A0(n870), .A1(n871), .A2(n872), .A3(n873) );
  inv01 U386 ( .Y(n748), .A(n747) );
  or04 U387 ( .Y(n749), .A0(s_opa_i_28_), .A1(n803), .A2(s_opa_i_27_), .A3(
        s_opa_i_26_) );
  inv01 U388 ( .Y(n750), .A(n749) );
  or03 U389 ( .Y(n751), .A0(s_rmode_i_0_), .A1(s_rmode_i_1_), .A2(n835) );
  inv01 U390 ( .Y(n752), .A(n751) );
  or04 U391 ( .Y(n753), .A0(s_opa_i_11_), .A1(n807), .A2(s_opa_i_10_), .A3(
        s_opa_i_0_) );
  inv01 U392 ( .Y(n754), .A(n753) );
  or04 U393 ( .Y(n755), .A0(n806), .A1(s_opa_i_14_), .A2(s_opa_i_16_), .A3(
        s_opa_i_15_) );
  inv01 U394 ( .Y(n756), .A(n755) );
  or04 U395 ( .Y(n757), .A0(n805), .A1(s_opa_i_1_), .A2(s_opa_i_21_), .A3(
        s_opa_i_20_) );
  inv01 U396 ( .Y(n758), .A(n757) );
  or04 U397 ( .Y(n759), .A0(n804), .A1(s_opa_i_4_), .A2(s_opa_i_6_), .A3(
        s_opa_i_5_) );
  inv01 U398 ( .Y(n760), .A(n759) );
  nand02 U399 ( .Y(n809), .A0(n761), .A1(n762) );
  inv02 U400 ( .Y(n763), .A(n832) );
  inv02 U401 ( .Y(n764), .A(s_fraco1_3_) );
  inv01 U402 ( .Y(n765), .A(n661) );
  inv01 U403 ( .Y(n766), .A(s_guard) );
  inv01 U404 ( .Y(n767), .A(s_rmode_i_1_) );
  inv01 U405 ( .Y(n768), .A(n752) );
  nand02 U406 ( .Y(n769), .A0(n765), .A1(n770) );
  nand02 U407 ( .Y(n771), .A0(n766), .A1(n772) );
  nand02 U408 ( .Y(n773), .A0(n767), .A1(n774) );
  nand02 U409 ( .Y(n775), .A0(n768), .A1(n776) );
  nand02 U410 ( .Y(n777), .A0(n768), .A1(n778) );
  nand02 U411 ( .Y(n779), .A0(n768), .A1(n780) );
  nand02 U412 ( .Y(n781), .A0(n763), .A1(n764) );
  inv01 U413 ( .Y(n770), .A(n781) );
  nand02 U414 ( .Y(n782), .A0(n763), .A1(n764) );
  inv01 U415 ( .Y(n772), .A(n782) );
  nand02 U416 ( .Y(n783), .A0(n763), .A1(n764) );
  inv01 U417 ( .Y(n774), .A(n783) );
  nand02 U418 ( .Y(n784), .A0(n763), .A1(n765) );
  inv01 U419 ( .Y(n776), .A(n784) );
  nand02 U420 ( .Y(n785), .A0(n763), .A1(n766) );
  inv01 U421 ( .Y(n778), .A(n785) );
  nand02 U422 ( .Y(n786), .A0(n763), .A1(n767) );
  inv01 U423 ( .Y(n780), .A(n786) );
  nand02 U424 ( .Y(n787), .A0(n769), .A1(n771) );
  inv01 U425 ( .Y(n788), .A(n787) );
  nand02 U426 ( .Y(n789), .A0(n773), .A1(n788) );
  inv01 U427 ( .Y(n761), .A(n789) );
  nand02 U428 ( .Y(n790), .A0(n775), .A1(n777) );
  inv01 U429 ( .Y(n791), .A(n790) );
  nand02 U430 ( .Y(n792), .A0(n779), .A1(n791) );
  inv01 U431 ( .Y(n762), .A(n792) );
  buf12 U432 ( .Y(n794), .A(n809) );
  buf16 U433 ( .Y(n793), .A(n795) );
  inv02 U434 ( .Y(n796), .A(n793) );
  nand02 U435 ( .Y(s_output_o_30_), .A0(n796), .A1(n843) );
  nand02 U436 ( .Y(s_output_o_29_), .A0(n796), .A1(n845) );
  nand02 U437 ( .Y(s_output_o_28_), .A0(n796), .A1(n846) );
  nand02 U438 ( .Y(s_output_o_27_), .A0(n796), .A1(n847) );
  nand02 U439 ( .Y(s_output_o_26_), .A0(n796), .A1(n848) );
  nand02 U440 ( .Y(s_output_o_25_), .A0(n796), .A1(n849) );
  nand02 U441 ( .Y(s_output_o_24_), .A0(n796), .A1(n850) );
  nand02 U442 ( .Y(s_output_o_23_), .A0(n796), .A1(n851) );
  nand02 U443 ( .Y(s_output_o_22_), .A0(n797), .A1(n798) );
  mux21 U444 ( .Y(n797), .A0(n735), .A1(s_frac_rnd_22_), .S0(n800) );
  and02 U445 ( .Y(s_ine_o), .A0(n796), .A1(s_sticky) );
  nand02 U446 ( .Y(n795), .A0(n798), .A1(n800) );
  nand02 U447 ( .Y(n800), .A0(n737), .A1(n748) );
  ao21 U448 ( .Y(n798), .A0(n801), .A1(n750), .B0(n802) );
  inv01 U449 ( .Y(n802), .A(s_sign_i) );
  nand02 U450 ( .Y(n803), .A0(n885), .A1(n886) );
  nand04 U451 ( .Y(n799), .A0(n754), .A1(n756), .A2(n758), .A3(n760) );
  nand03 U452 ( .Y(n804), .A0(n875), .A1(n876), .A2(n874) );
  nand03 U453 ( .Y(n805), .A0(n878), .A1(n879), .A2(n877) );
  nand03 U454 ( .Y(n806), .A0(n881), .A1(n882), .A2(n880) );
  nand02 U455 ( .Y(n807), .A0(n883), .A1(n884) );
  mux21 U456 ( .Y(s_frac_rnd254_9_), .A0(n808), .A1(n887), .S0(n794) );
  inv01 U457 ( .Y(n808), .A(n____return281_9_) );
  mux21 U458 ( .Y(s_frac_rnd254_8_), .A0(n810), .A1(n888), .S0(n794) );
  inv01 U459 ( .Y(n810), .A(n____return281_8_) );
  mux21 U460 ( .Y(s_frac_rnd254_7_), .A0(n811), .A1(n889), .S0(n794) );
  inv01 U461 ( .Y(n811), .A(n____return281_7_) );
  mux21 U462 ( .Y(s_frac_rnd254_6_), .A0(n812), .A1(n890), .S0(n794) );
  inv01 U463 ( .Y(n812), .A(n____return281_6_) );
  mux21 U464 ( .Y(s_frac_rnd254_5_), .A0(n813), .A1(n891), .S0(n794) );
  inv01 U465 ( .Y(n813), .A(n____return281_5_) );
  mux21 U466 ( .Y(s_frac_rnd254_4_), .A0(n814), .A1(n892), .S0(n794) );
  inv01 U467 ( .Y(n814), .A(n____return281_4_) );
  mux21 U468 ( .Y(s_frac_rnd254_3_), .A0(n815), .A1(n893), .S0(n794) );
  inv01 U469 ( .Y(n815), .A(n____return281_3_) );
  mux21 U470 ( .Y(s_frac_rnd254_2_), .A0(n816), .A1(n894), .S0(n794) );
  inv01 U471 ( .Y(n816), .A(n____return281_2_) );
  mux21 U472 ( .Y(s_frac_rnd254_22_), .A0(n817), .A1(n895), .S0(n794) );
  inv01 U473 ( .Y(n817), .A(n283_22_) );
  mux21 U474 ( .Y(s_frac_rnd254_21_), .A0(n818), .A1(n896), .S0(n794) );
  inv01 U475 ( .Y(n818), .A(n____return281_21_) );
  mux21 U476 ( .Y(s_frac_rnd254_20_), .A0(n819), .A1(n897), .S0(n794) );
  inv01 U477 ( .Y(n819), .A(n____return281_20_) );
  inv01 U478 ( .Y(s_frac_rnd254_1_), .A(n820) );
  mux21 U479 ( .Y(n820), .A0(n____return281_1_), .A1(s_fraco1_3_), .S0(n794)
         );
  mux21 U480 ( .Y(s_frac_rnd254_19_), .A0(n821), .A1(n898), .S0(n794) );
  inv01 U481 ( .Y(n821), .A(n____return281_19_) );
  inv01 U482 ( .Y(n822), .A(n____return281_18_) );
  mux21 U483 ( .Y(s_frac_rnd254_17_), .A0(n823), .A1(n900), .S0(n794) );
  inv01 U484 ( .Y(n823), .A(n____return281_17_) );
  mux21 U485 ( .Y(s_frac_rnd254_16_), .A0(n824), .A1(n901), .S0(n794) );
  inv01 U486 ( .Y(n824), .A(n____return281_16_) );
  mux21 U487 ( .Y(s_frac_rnd254_15_), .A0(n825), .A1(n902), .S0(n794) );
  inv01 U488 ( .Y(n825), .A(n____return281_15_) );
  mux21 U489 ( .Y(s_frac_rnd254_14_), .A0(n826), .A1(n903), .S0(n794) );
  inv01 U490 ( .Y(n826), .A(n____return281_14_) );
  mux21 U491 ( .Y(s_frac_rnd254_13_), .A0(n827), .A1(n904), .S0(n794) );
  inv01 U492 ( .Y(n827), .A(n____return281_13_) );
  mux21 U493 ( .Y(s_frac_rnd254_12_), .A0(n828), .A1(n905), .S0(n794) );
  inv01 U494 ( .Y(n828), .A(n____return281_12_) );
  mux21 U495 ( .Y(s_frac_rnd254_11_), .A0(n829), .A1(n906), .S0(n794) );
  inv01 U496 ( .Y(n829), .A(n____return281_11_) );
  mux21 U497 ( .Y(s_frac_rnd254_10_), .A0(n830), .A1(n907), .S0(n794) );
  inv01 U498 ( .Y(n830), .A(n____return281_10_) );
  mux21 U499 ( .Y(s_frac_rnd254_0_), .A0(n831), .A1(n908), .S0(n794) );
  inv01 U500 ( .Y(n832), .A(n833) );
  ao21 U501 ( .Y(n834), .A0(s_rmode_i_1_), .A1(n661), .B0(n752) );
  inv01 U502 ( .Y(n835), .A(s_guard) );
  inv01 U503 ( .Y(n831), .A(n____return281_0_) );
  post_norm_sqrt_DW01_inc_23_0 add_136_plus_plus ( .A({s_fraco1_24_, 
        s_fraco1_23_, s_fraco1_22_, s_fraco1_21_, s_fraco1_20_, s_fraco1_19_, 
        s_fraco1_18_, s_fraco1_17_, s_fraco1_16_, s_fraco1_15_, s_fraco1_14_, 
        s_fraco1_13_, s_fraco1_12_, s_fraco1_11_, s_fraco1_10_, s_fraco1_9_, 
        s_fraco1_8_, s_fraco1_7_, s_fraco1_6_, s_fraco1_5_, s_fraco1_4_, 
        s_fraco1_3_, s_fraco1_2_}), .SUM({n283_22_, n____return281_21_, 
        n____return281_20_, n____return281_19_, n____return281_18_, 
        n____return281_17_, n____return281_16_, n____return281_15_, 
        n____return281_14_, n____return281_13_, n____return281_12_, 
        n____return281_11_, n____return281_10_, n____return281_9_, 
        n____return281_8_, n____return281_7_, n____return281_6_, 
        n____return281_5_, n____return281_4_, n____return281_3_, 
        n____return281_2_, n____return281_1_, n____return281_0_}) );
endmodule


module mul_24_DW01_add_48_2 ( A, B, CI, SUM, CO );
  input [47:0] A;
  input [47:0] B;
  output [47:0] SUM;
  input CI;
  output CO;
  wire   carry_47_, carry_37_, carry_36_, carry_35_, carry_34_, carry_33_,
         carry_32_, carry_31_, carry_30_, carry_29_, carry_28_, carry_27_,
         carry_26_, carry_25_, carry_24_, carry_23_, carry_22_, carry_21_,
         carry_20_, carry_19_, carry_18_, carry_17_, carry_16_, carry_15_,
         carry_14_, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_,
         B_1_, B_0_, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380;
  assign SUM[11] = B_11_;
  assign B_11_ = B[11];
  assign SUM[10] = B_10_;
  assign B_10_ = B[10];
  assign SUM[9] = B_9_;
  assign B_9_ = B[9];
  assign SUM[8] = B_8_;
  assign B_8_ = B[8];
  assign SUM[7] = B_7_;
  assign B_7_ = B[7];
  assign SUM[6] = B_6_;
  assign B_6_ = B[6];
  assign SUM[5] = B_5_;
  assign B_5_ = B[5];
  assign SUM[4] = B_4_;
  assign B_4_ = B[4];
  assign SUM[3] = B_3_;
  assign B_3_ = B[3];
  assign SUM[2] = B_2_;
  assign B_2_ = B[2];
  assign SUM[1] = B_1_;
  assign B_1_ = B[1];
  assign SUM[0] = B_0_;
  assign B_0_ = B[0];

  buf02 U4 ( .Y(SUM[19]), .A(n385) );
  buf02 U5 ( .Y(SUM[16]), .A(n388) );
  buf02 U6 ( .Y(SUM[18]), .A(n386) );
  buf02 U7 ( .Y(SUM[14]), .A(n390) );
  buf02 U8 ( .Y(SUM[23]), .A(n381) );
  buf02 U9 ( .Y(SUM[21]), .A(n383) );
  buf02 U10 ( .Y(SUM[17]), .A(n387) );
  buf02 U11 ( .Y(SUM[22]), .A(n382) );
  buf02 U12 ( .Y(SUM[13]), .A(n391) );
  buf02 U13 ( .Y(SUM[15]), .A(n389) );
  buf02 U14 ( .Y(SUM[20]), .A(n384) );
  nand02 U15 ( .Y(n12), .A0(A[12]), .A1(B[12]) );
  inv02 U16 ( .Y(n13), .A(n12) );
  nand02 U17 ( .Y(n14), .A0(n23), .A1(A[40]) );
  inv02 U18 ( .Y(n15), .A(n14) );
  nand02 U19 ( .Y(n16), .A0(n25), .A1(A[43]) );
  inv02 U20 ( .Y(n17), .A(n16) );
  nand02 U21 ( .Y(n18), .A0(n29), .A1(A[45]) );
  inv02 U22 ( .Y(n19), .A(n18) );
  nand02 U23 ( .Y(n20), .A0(carry_37_), .A1(A[37]) );
  inv02 U24 ( .Y(n21), .A(n20) );
  nand02 U25 ( .Y(n22), .A0(n27), .A1(A[39]) );
  inv02 U26 ( .Y(n23), .A(n22) );
  nand02 U27 ( .Y(n24), .A0(n31), .A1(A[42]) );
  inv02 U28 ( .Y(n25), .A(n24) );
  nand02 U29 ( .Y(n26), .A0(n21), .A1(A[38]) );
  inv02 U30 ( .Y(n27), .A(n26) );
  nand02 U31 ( .Y(n28), .A0(n17), .A1(A[44]) );
  inv02 U32 ( .Y(n29), .A(n28) );
  nand02 U33 ( .Y(n30), .A0(n15), .A1(A[41]) );
  inv02 U34 ( .Y(n31), .A(n30) );
  buf02 U35 ( .Y(n32), .A(carry_23_) );
  buf02 U36 ( .Y(n33), .A(carry_22_) );
  buf02 U37 ( .Y(n34), .A(carry_21_) );
  buf02 U38 ( .Y(n35), .A(carry_20_) );
  buf02 U39 ( .Y(n36), .A(carry_19_) );
  buf02 U40 ( .Y(n37), .A(carry_18_) );
  buf02 U41 ( .Y(n38), .A(carry_17_) );
  buf02 U42 ( .Y(n39), .A(carry_16_) );
  buf02 U43 ( .Y(n40), .A(carry_15_) );
  buf02 U44 ( .Y(n41), .A(carry_14_) );
  buf02 U45 ( .Y(n42), .A(carry_24_) );
  inv01 U46 ( .Y(SUM[24]), .A(n43) );
  inv02 U47 ( .Y(carry_25_), .A(n44) );
  inv02 U48 ( .Y(n45), .A(B[24]) );
  inv02 U49 ( .Y(n46), .A(A[24]) );
  inv02 U50 ( .Y(n47), .A(n42) );
  nor02 U51 ( .Y(n48), .A0(n45), .A1(n49) );
  nor02 U52 ( .Y(n50), .A0(n46), .A1(n51) );
  nor02 U53 ( .Y(n52), .A0(n47), .A1(n53) );
  nor02 U54 ( .Y(n54), .A0(n47), .A1(n55) );
  nor02 U55 ( .Y(n43), .A0(n56), .A1(n57) );
  nor02 U56 ( .Y(n58), .A0(n46), .A1(n47) );
  nor02 U57 ( .Y(n59), .A0(n45), .A1(n47) );
  nor02 U58 ( .Y(n60), .A0(n45), .A1(n46) );
  nor02 U59 ( .Y(n44), .A0(n60), .A1(n61) );
  nor02 U60 ( .Y(n62), .A0(A[24]), .A1(n42) );
  inv01 U61 ( .Y(n49), .A(n62) );
  nor02 U62 ( .Y(n63), .A0(B[24]), .A1(n42) );
  inv01 U63 ( .Y(n51), .A(n63) );
  nor02 U64 ( .Y(n64), .A0(B[24]), .A1(A[24]) );
  inv01 U65 ( .Y(n53), .A(n64) );
  nor02 U66 ( .Y(n65), .A0(n45), .A1(n46) );
  inv01 U67 ( .Y(n55), .A(n65) );
  nor02 U68 ( .Y(n66), .A0(n48), .A1(n50) );
  inv01 U69 ( .Y(n56), .A(n66) );
  nor02 U70 ( .Y(n67), .A0(n52), .A1(n54) );
  inv01 U71 ( .Y(n57), .A(n67) );
  nor02 U72 ( .Y(n68), .A0(n58), .A1(n59) );
  inv01 U73 ( .Y(n61), .A(n68) );
  inv01 U74 ( .Y(SUM[25]), .A(n69) );
  inv02 U75 ( .Y(carry_26_), .A(n70) );
  inv02 U76 ( .Y(n71), .A(B[25]) );
  inv02 U77 ( .Y(n72), .A(A[25]) );
  inv02 U78 ( .Y(n73), .A(carry_25_) );
  nor02 U79 ( .Y(n74), .A0(n71), .A1(n75) );
  nor02 U80 ( .Y(n76), .A0(n72), .A1(n77) );
  nor02 U81 ( .Y(n78), .A0(n73), .A1(n79) );
  nor02 U82 ( .Y(n80), .A0(n73), .A1(n81) );
  nor02 U83 ( .Y(n69), .A0(n82), .A1(n83) );
  nor02 U84 ( .Y(n84), .A0(n72), .A1(n73) );
  nor02 U85 ( .Y(n85), .A0(n71), .A1(n73) );
  nor02 U86 ( .Y(n86), .A0(n71), .A1(n72) );
  nor02 U87 ( .Y(n70), .A0(n86), .A1(n87) );
  nor02 U88 ( .Y(n88), .A0(A[25]), .A1(carry_25_) );
  inv01 U89 ( .Y(n75), .A(n88) );
  nor02 U90 ( .Y(n89), .A0(B[25]), .A1(carry_25_) );
  inv01 U91 ( .Y(n77), .A(n89) );
  nor02 U92 ( .Y(n90), .A0(B[25]), .A1(A[25]) );
  inv01 U93 ( .Y(n79), .A(n90) );
  nor02 U94 ( .Y(n91), .A0(n71), .A1(n72) );
  inv01 U95 ( .Y(n81), .A(n91) );
  nor02 U96 ( .Y(n92), .A0(n74), .A1(n76) );
  inv01 U97 ( .Y(n82), .A(n92) );
  nor02 U98 ( .Y(n93), .A0(n78), .A1(n80) );
  inv01 U99 ( .Y(n83), .A(n93) );
  nor02 U100 ( .Y(n94), .A0(n84), .A1(n85) );
  inv01 U101 ( .Y(n87), .A(n94) );
  inv01 U102 ( .Y(SUM[26]), .A(n95) );
  inv02 U103 ( .Y(carry_27_), .A(n96) );
  inv02 U104 ( .Y(n97), .A(B[26]) );
  inv02 U105 ( .Y(n98), .A(A[26]) );
  inv02 U106 ( .Y(n99), .A(carry_26_) );
  nor02 U107 ( .Y(n100), .A0(n97), .A1(n101) );
  nor02 U108 ( .Y(n102), .A0(n98), .A1(n103) );
  nor02 U109 ( .Y(n104), .A0(n99), .A1(n105) );
  nor02 U110 ( .Y(n106), .A0(n99), .A1(n107) );
  nor02 U111 ( .Y(n95), .A0(n108), .A1(n109) );
  nor02 U112 ( .Y(n110), .A0(n98), .A1(n99) );
  nor02 U113 ( .Y(n111), .A0(n97), .A1(n99) );
  nor02 U114 ( .Y(n112), .A0(n97), .A1(n98) );
  nor02 U115 ( .Y(n96), .A0(n112), .A1(n113) );
  nor02 U116 ( .Y(n114), .A0(A[26]), .A1(carry_26_) );
  inv01 U117 ( .Y(n101), .A(n114) );
  nor02 U118 ( .Y(n115), .A0(B[26]), .A1(carry_26_) );
  inv01 U119 ( .Y(n103), .A(n115) );
  nor02 U120 ( .Y(n116), .A0(B[26]), .A1(A[26]) );
  inv01 U121 ( .Y(n105), .A(n116) );
  nor02 U122 ( .Y(n117), .A0(n97), .A1(n98) );
  inv01 U123 ( .Y(n107), .A(n117) );
  nor02 U124 ( .Y(n118), .A0(n100), .A1(n102) );
  inv01 U125 ( .Y(n108), .A(n118) );
  nor02 U126 ( .Y(n119), .A0(n104), .A1(n106) );
  inv01 U127 ( .Y(n109), .A(n119) );
  nor02 U128 ( .Y(n120), .A0(n110), .A1(n111) );
  inv01 U129 ( .Y(n113), .A(n120) );
  inv01 U130 ( .Y(SUM[27]), .A(n121) );
  inv02 U131 ( .Y(carry_28_), .A(n122) );
  inv02 U132 ( .Y(n123), .A(B[27]) );
  inv02 U133 ( .Y(n124), .A(A[27]) );
  inv02 U134 ( .Y(n125), .A(carry_27_) );
  nor02 U135 ( .Y(n126), .A0(n123), .A1(n127) );
  nor02 U136 ( .Y(n128), .A0(n124), .A1(n129) );
  nor02 U137 ( .Y(n130), .A0(n125), .A1(n131) );
  nor02 U138 ( .Y(n132), .A0(n125), .A1(n133) );
  nor02 U139 ( .Y(n121), .A0(n134), .A1(n135) );
  nor02 U140 ( .Y(n136), .A0(n124), .A1(n125) );
  nor02 U141 ( .Y(n137), .A0(n123), .A1(n125) );
  nor02 U142 ( .Y(n138), .A0(n123), .A1(n124) );
  nor02 U143 ( .Y(n122), .A0(n138), .A1(n139) );
  nor02 U144 ( .Y(n140), .A0(A[27]), .A1(carry_27_) );
  inv01 U145 ( .Y(n127), .A(n140) );
  nor02 U146 ( .Y(n141), .A0(B[27]), .A1(carry_27_) );
  inv01 U147 ( .Y(n129), .A(n141) );
  nor02 U148 ( .Y(n142), .A0(B[27]), .A1(A[27]) );
  inv01 U149 ( .Y(n131), .A(n142) );
  nor02 U150 ( .Y(n143), .A0(n123), .A1(n124) );
  inv01 U151 ( .Y(n133), .A(n143) );
  nor02 U152 ( .Y(n144), .A0(n126), .A1(n128) );
  inv01 U153 ( .Y(n134), .A(n144) );
  nor02 U154 ( .Y(n145), .A0(n130), .A1(n132) );
  inv01 U155 ( .Y(n135), .A(n145) );
  nor02 U156 ( .Y(n146), .A0(n136), .A1(n137) );
  inv01 U157 ( .Y(n139), .A(n146) );
  inv01 U158 ( .Y(SUM[28]), .A(n147) );
  inv02 U159 ( .Y(carry_29_), .A(n148) );
  inv02 U160 ( .Y(n149), .A(B[28]) );
  inv02 U161 ( .Y(n150), .A(A[28]) );
  inv02 U162 ( .Y(n151), .A(carry_28_) );
  nor02 U163 ( .Y(n152), .A0(n149), .A1(n153) );
  nor02 U164 ( .Y(n154), .A0(n150), .A1(n155) );
  nor02 U165 ( .Y(n156), .A0(n151), .A1(n157) );
  nor02 U166 ( .Y(n158), .A0(n151), .A1(n159) );
  nor02 U167 ( .Y(n147), .A0(n160), .A1(n161) );
  nor02 U168 ( .Y(n162), .A0(n150), .A1(n151) );
  nor02 U169 ( .Y(n163), .A0(n149), .A1(n151) );
  nor02 U170 ( .Y(n164), .A0(n149), .A1(n150) );
  nor02 U171 ( .Y(n148), .A0(n164), .A1(n165) );
  nor02 U172 ( .Y(n166), .A0(A[28]), .A1(carry_28_) );
  inv01 U173 ( .Y(n153), .A(n166) );
  nor02 U174 ( .Y(n167), .A0(B[28]), .A1(carry_28_) );
  inv01 U175 ( .Y(n155), .A(n167) );
  nor02 U176 ( .Y(n168), .A0(B[28]), .A1(A[28]) );
  inv01 U177 ( .Y(n157), .A(n168) );
  nor02 U178 ( .Y(n169), .A0(n149), .A1(n150) );
  inv01 U179 ( .Y(n159), .A(n169) );
  nor02 U180 ( .Y(n170), .A0(n152), .A1(n154) );
  inv01 U181 ( .Y(n160), .A(n170) );
  nor02 U182 ( .Y(n171), .A0(n156), .A1(n158) );
  inv01 U183 ( .Y(n161), .A(n171) );
  nor02 U184 ( .Y(n172), .A0(n162), .A1(n163) );
  inv01 U185 ( .Y(n165), .A(n172) );
  inv01 U186 ( .Y(SUM[29]), .A(n173) );
  inv02 U187 ( .Y(carry_30_), .A(n174) );
  inv02 U188 ( .Y(n175), .A(B[29]) );
  inv02 U189 ( .Y(n176), .A(A[29]) );
  inv02 U190 ( .Y(n177), .A(carry_29_) );
  nor02 U191 ( .Y(n178), .A0(n175), .A1(n179) );
  nor02 U192 ( .Y(n180), .A0(n176), .A1(n181) );
  nor02 U193 ( .Y(n182), .A0(n177), .A1(n183) );
  nor02 U194 ( .Y(n184), .A0(n177), .A1(n185) );
  nor02 U195 ( .Y(n173), .A0(n186), .A1(n187) );
  nor02 U196 ( .Y(n188), .A0(n176), .A1(n177) );
  nor02 U197 ( .Y(n189), .A0(n175), .A1(n177) );
  nor02 U198 ( .Y(n190), .A0(n175), .A1(n176) );
  nor02 U199 ( .Y(n174), .A0(n190), .A1(n191) );
  nor02 U200 ( .Y(n192), .A0(A[29]), .A1(carry_29_) );
  inv01 U201 ( .Y(n179), .A(n192) );
  nor02 U202 ( .Y(n193), .A0(B[29]), .A1(carry_29_) );
  inv01 U203 ( .Y(n181), .A(n193) );
  nor02 U204 ( .Y(n194), .A0(B[29]), .A1(A[29]) );
  inv01 U205 ( .Y(n183), .A(n194) );
  nor02 U206 ( .Y(n195), .A0(n175), .A1(n176) );
  inv01 U207 ( .Y(n185), .A(n195) );
  nor02 U208 ( .Y(n196), .A0(n178), .A1(n180) );
  inv01 U209 ( .Y(n186), .A(n196) );
  nor02 U210 ( .Y(n197), .A0(n182), .A1(n184) );
  inv01 U211 ( .Y(n187), .A(n197) );
  nor02 U212 ( .Y(n198), .A0(n188), .A1(n189) );
  inv01 U213 ( .Y(n191), .A(n198) );
  inv01 U214 ( .Y(SUM[30]), .A(n199) );
  inv02 U215 ( .Y(carry_31_), .A(n200) );
  inv02 U216 ( .Y(n201), .A(B[30]) );
  inv02 U217 ( .Y(n202), .A(A[30]) );
  inv02 U218 ( .Y(n203), .A(carry_30_) );
  nor02 U219 ( .Y(n204), .A0(n201), .A1(n205) );
  nor02 U220 ( .Y(n206), .A0(n202), .A1(n207) );
  nor02 U221 ( .Y(n208), .A0(n203), .A1(n209) );
  nor02 U222 ( .Y(n210), .A0(n203), .A1(n211) );
  nor02 U223 ( .Y(n199), .A0(n212), .A1(n213) );
  nor02 U224 ( .Y(n214), .A0(n202), .A1(n203) );
  nor02 U225 ( .Y(n215), .A0(n201), .A1(n203) );
  nor02 U226 ( .Y(n216), .A0(n201), .A1(n202) );
  nor02 U227 ( .Y(n200), .A0(n216), .A1(n217) );
  nor02 U228 ( .Y(n218), .A0(A[30]), .A1(carry_30_) );
  inv01 U229 ( .Y(n205), .A(n218) );
  nor02 U230 ( .Y(n219), .A0(B[30]), .A1(carry_30_) );
  inv01 U231 ( .Y(n207), .A(n219) );
  nor02 U232 ( .Y(n220), .A0(B[30]), .A1(A[30]) );
  inv01 U233 ( .Y(n209), .A(n220) );
  nor02 U234 ( .Y(n221), .A0(n201), .A1(n202) );
  inv01 U235 ( .Y(n211), .A(n221) );
  nor02 U236 ( .Y(n222), .A0(n204), .A1(n206) );
  inv01 U237 ( .Y(n212), .A(n222) );
  nor02 U238 ( .Y(n223), .A0(n208), .A1(n210) );
  inv01 U239 ( .Y(n213), .A(n223) );
  nor02 U240 ( .Y(n224), .A0(n214), .A1(n215) );
  inv01 U241 ( .Y(n217), .A(n224) );
  inv01 U242 ( .Y(SUM[31]), .A(n225) );
  inv02 U243 ( .Y(carry_32_), .A(n226) );
  inv02 U244 ( .Y(n227), .A(B[31]) );
  inv02 U245 ( .Y(n228), .A(A[31]) );
  inv02 U246 ( .Y(n229), .A(carry_31_) );
  nor02 U247 ( .Y(n230), .A0(n227), .A1(n231) );
  nor02 U248 ( .Y(n232), .A0(n228), .A1(n233) );
  nor02 U249 ( .Y(n234), .A0(n229), .A1(n235) );
  nor02 U250 ( .Y(n236), .A0(n229), .A1(n237) );
  nor02 U251 ( .Y(n225), .A0(n238), .A1(n239) );
  nor02 U252 ( .Y(n240), .A0(n228), .A1(n229) );
  nor02 U253 ( .Y(n241), .A0(n227), .A1(n229) );
  nor02 U254 ( .Y(n242), .A0(n227), .A1(n228) );
  nor02 U255 ( .Y(n226), .A0(n242), .A1(n243) );
  nor02 U256 ( .Y(n244), .A0(A[31]), .A1(carry_31_) );
  inv01 U257 ( .Y(n231), .A(n244) );
  nor02 U258 ( .Y(n245), .A0(B[31]), .A1(carry_31_) );
  inv01 U259 ( .Y(n233), .A(n245) );
  nor02 U260 ( .Y(n246), .A0(B[31]), .A1(A[31]) );
  inv01 U261 ( .Y(n235), .A(n246) );
  nor02 U262 ( .Y(n247), .A0(n227), .A1(n228) );
  inv01 U263 ( .Y(n237), .A(n247) );
  nor02 U264 ( .Y(n248), .A0(n230), .A1(n232) );
  inv01 U265 ( .Y(n238), .A(n248) );
  nor02 U266 ( .Y(n249), .A0(n234), .A1(n236) );
  inv01 U267 ( .Y(n239), .A(n249) );
  nor02 U268 ( .Y(n250), .A0(n240), .A1(n241) );
  inv01 U269 ( .Y(n243), .A(n250) );
  inv01 U270 ( .Y(SUM[32]), .A(n251) );
  inv02 U271 ( .Y(carry_33_), .A(n252) );
  inv02 U272 ( .Y(n253), .A(B[32]) );
  inv02 U273 ( .Y(n254), .A(A[32]) );
  inv02 U274 ( .Y(n255), .A(carry_32_) );
  nor02 U275 ( .Y(n256), .A0(n253), .A1(n257) );
  nor02 U276 ( .Y(n258), .A0(n254), .A1(n259) );
  nor02 U277 ( .Y(n260), .A0(n255), .A1(n261) );
  nor02 U278 ( .Y(n262), .A0(n255), .A1(n263) );
  nor02 U279 ( .Y(n251), .A0(n264), .A1(n265) );
  nor02 U280 ( .Y(n266), .A0(n254), .A1(n255) );
  nor02 U281 ( .Y(n267), .A0(n253), .A1(n255) );
  nor02 U282 ( .Y(n268), .A0(n253), .A1(n254) );
  nor02 U283 ( .Y(n252), .A0(n268), .A1(n269) );
  nor02 U284 ( .Y(n270), .A0(A[32]), .A1(carry_32_) );
  inv01 U285 ( .Y(n257), .A(n270) );
  nor02 U286 ( .Y(n271), .A0(B[32]), .A1(carry_32_) );
  inv01 U287 ( .Y(n259), .A(n271) );
  nor02 U288 ( .Y(n272), .A0(B[32]), .A1(A[32]) );
  inv01 U289 ( .Y(n261), .A(n272) );
  nor02 U290 ( .Y(n273), .A0(n253), .A1(n254) );
  inv01 U291 ( .Y(n263), .A(n273) );
  nor02 U292 ( .Y(n274), .A0(n256), .A1(n258) );
  inv01 U293 ( .Y(n264), .A(n274) );
  nor02 U294 ( .Y(n275), .A0(n260), .A1(n262) );
  inv01 U295 ( .Y(n265), .A(n275) );
  nor02 U296 ( .Y(n276), .A0(n266), .A1(n267) );
  inv01 U297 ( .Y(n269), .A(n276) );
  inv01 U298 ( .Y(SUM[33]), .A(n277) );
  inv02 U299 ( .Y(carry_34_), .A(n278) );
  inv02 U300 ( .Y(n279), .A(B[33]) );
  inv02 U301 ( .Y(n280), .A(A[33]) );
  inv02 U302 ( .Y(n281), .A(carry_33_) );
  nor02 U303 ( .Y(n282), .A0(n279), .A1(n283) );
  nor02 U304 ( .Y(n284), .A0(n280), .A1(n285) );
  nor02 U305 ( .Y(n286), .A0(n281), .A1(n287) );
  nor02 U306 ( .Y(n288), .A0(n281), .A1(n289) );
  nor02 U307 ( .Y(n277), .A0(n290), .A1(n291) );
  nor02 U308 ( .Y(n292), .A0(n280), .A1(n281) );
  nor02 U309 ( .Y(n293), .A0(n279), .A1(n281) );
  nor02 U310 ( .Y(n294), .A0(n279), .A1(n280) );
  nor02 U311 ( .Y(n278), .A0(n294), .A1(n295) );
  nor02 U312 ( .Y(n296), .A0(A[33]), .A1(carry_33_) );
  inv01 U313 ( .Y(n283), .A(n296) );
  nor02 U314 ( .Y(n297), .A0(B[33]), .A1(carry_33_) );
  inv01 U315 ( .Y(n285), .A(n297) );
  nor02 U316 ( .Y(n298), .A0(B[33]), .A1(A[33]) );
  inv01 U317 ( .Y(n287), .A(n298) );
  nor02 U318 ( .Y(n299), .A0(n279), .A1(n280) );
  inv01 U319 ( .Y(n289), .A(n299) );
  nor02 U320 ( .Y(n300), .A0(n282), .A1(n284) );
  inv01 U321 ( .Y(n290), .A(n300) );
  nor02 U322 ( .Y(n301), .A0(n286), .A1(n288) );
  inv01 U323 ( .Y(n291), .A(n301) );
  nor02 U324 ( .Y(n302), .A0(n292), .A1(n293) );
  inv01 U325 ( .Y(n295), .A(n302) );
  inv01 U326 ( .Y(SUM[34]), .A(n303) );
  inv02 U327 ( .Y(carry_35_), .A(n304) );
  inv02 U328 ( .Y(n305), .A(B[34]) );
  inv02 U329 ( .Y(n306), .A(A[34]) );
  inv02 U330 ( .Y(n307), .A(carry_34_) );
  nor02 U331 ( .Y(n308), .A0(n305), .A1(n309) );
  nor02 U332 ( .Y(n310), .A0(n306), .A1(n311) );
  nor02 U333 ( .Y(n312), .A0(n307), .A1(n313) );
  nor02 U334 ( .Y(n314), .A0(n307), .A1(n315) );
  nor02 U335 ( .Y(n303), .A0(n316), .A1(n317) );
  nor02 U336 ( .Y(n318), .A0(n306), .A1(n307) );
  nor02 U337 ( .Y(n319), .A0(n305), .A1(n307) );
  nor02 U338 ( .Y(n320), .A0(n305), .A1(n306) );
  nor02 U339 ( .Y(n304), .A0(n320), .A1(n321) );
  nor02 U340 ( .Y(n322), .A0(A[34]), .A1(carry_34_) );
  inv01 U341 ( .Y(n309), .A(n322) );
  nor02 U342 ( .Y(n323), .A0(B[34]), .A1(carry_34_) );
  inv01 U343 ( .Y(n311), .A(n323) );
  nor02 U344 ( .Y(n324), .A0(B[34]), .A1(A[34]) );
  inv01 U345 ( .Y(n313), .A(n324) );
  nor02 U346 ( .Y(n325), .A0(n305), .A1(n306) );
  inv01 U347 ( .Y(n315), .A(n325) );
  nor02 U348 ( .Y(n326), .A0(n308), .A1(n310) );
  inv01 U349 ( .Y(n316), .A(n326) );
  nor02 U350 ( .Y(n327), .A0(n312), .A1(n314) );
  inv01 U351 ( .Y(n317), .A(n327) );
  nor02 U352 ( .Y(n328), .A0(n318), .A1(n319) );
  inv01 U353 ( .Y(n321), .A(n328) );
  inv01 U354 ( .Y(SUM[35]), .A(n329) );
  inv02 U355 ( .Y(carry_36_), .A(n330) );
  inv02 U356 ( .Y(n331), .A(B[35]) );
  inv02 U357 ( .Y(n332), .A(A[35]) );
  inv02 U358 ( .Y(n333), .A(carry_35_) );
  nor02 U359 ( .Y(n334), .A0(n331), .A1(n335) );
  nor02 U360 ( .Y(n336), .A0(n332), .A1(n337) );
  nor02 U361 ( .Y(n338), .A0(n333), .A1(n339) );
  nor02 U362 ( .Y(n340), .A0(n333), .A1(n341) );
  nor02 U363 ( .Y(n329), .A0(n342), .A1(n343) );
  nor02 U364 ( .Y(n344), .A0(n332), .A1(n333) );
  nor02 U365 ( .Y(n345), .A0(n331), .A1(n333) );
  nor02 U366 ( .Y(n346), .A0(n331), .A1(n332) );
  nor02 U367 ( .Y(n330), .A0(n346), .A1(n347) );
  nor02 U368 ( .Y(n348), .A0(A[35]), .A1(carry_35_) );
  inv01 U369 ( .Y(n335), .A(n348) );
  nor02 U370 ( .Y(n349), .A0(B[35]), .A1(carry_35_) );
  inv01 U371 ( .Y(n337), .A(n349) );
  nor02 U372 ( .Y(n350), .A0(B[35]), .A1(A[35]) );
  inv01 U373 ( .Y(n339), .A(n350) );
  nor02 U374 ( .Y(n351), .A0(n331), .A1(n332) );
  inv01 U375 ( .Y(n341), .A(n351) );
  nor02 U376 ( .Y(n352), .A0(n334), .A1(n336) );
  inv01 U377 ( .Y(n342), .A(n352) );
  nor02 U378 ( .Y(n353), .A0(n338), .A1(n340) );
  inv01 U379 ( .Y(n343), .A(n353) );
  nor02 U380 ( .Y(n354), .A0(n344), .A1(n345) );
  inv01 U381 ( .Y(n347), .A(n354) );
  inv01 U382 ( .Y(SUM[36]), .A(n355) );
  inv02 U383 ( .Y(carry_37_), .A(n356) );
  inv02 U384 ( .Y(n357), .A(B[36]) );
  inv02 U385 ( .Y(n358), .A(A[36]) );
  inv02 U386 ( .Y(n359), .A(carry_36_) );
  nor02 U387 ( .Y(n360), .A0(n357), .A1(n361) );
  nor02 U388 ( .Y(n362), .A0(n358), .A1(n363) );
  nor02 U389 ( .Y(n364), .A0(n359), .A1(n365) );
  nor02 U390 ( .Y(n366), .A0(n359), .A1(n367) );
  nor02 U391 ( .Y(n355), .A0(n368), .A1(n369) );
  nor02 U392 ( .Y(n370), .A0(n358), .A1(n359) );
  nor02 U393 ( .Y(n371), .A0(n357), .A1(n359) );
  nor02 U394 ( .Y(n372), .A0(n357), .A1(n358) );
  nor02 U395 ( .Y(n356), .A0(n372), .A1(n373) );
  nor02 U396 ( .Y(n374), .A0(A[36]), .A1(carry_36_) );
  inv01 U397 ( .Y(n361), .A(n374) );
  nor02 U398 ( .Y(n375), .A0(B[36]), .A1(carry_36_) );
  inv01 U399 ( .Y(n363), .A(n375) );
  nor02 U400 ( .Y(n376), .A0(B[36]), .A1(A[36]) );
  inv01 U401 ( .Y(n365), .A(n376) );
  nor02 U402 ( .Y(n377), .A0(n357), .A1(n358) );
  inv01 U403 ( .Y(n367), .A(n377) );
  nor02 U404 ( .Y(n378), .A0(n360), .A1(n362) );
  inv01 U405 ( .Y(n368), .A(n378) );
  nor02 U406 ( .Y(n379), .A0(n364), .A1(n366) );
  inv01 U407 ( .Y(n369), .A(n379) );
  nor02 U408 ( .Y(n380), .A0(n370), .A1(n371) );
  inv01 U409 ( .Y(n373), .A(n380) );
  xor2 U410 ( .Y(SUM[47]), .A0(A[47]), .A1(carry_47_) );
  and02 U411 ( .Y(carry_47_), .A0(n19), .A1(A[46]) );
  xor2 U412 ( .Y(SUM[46]), .A0(A[46]), .A1(n19) );
  xor2 U413 ( .Y(SUM[45]), .A0(A[45]), .A1(n29) );
  xor2 U414 ( .Y(SUM[44]), .A0(A[44]), .A1(n17) );
  xor2 U415 ( .Y(SUM[43]), .A0(A[43]), .A1(n25) );
  xor2 U416 ( .Y(SUM[42]), .A0(A[42]), .A1(n31) );
  xor2 U417 ( .Y(SUM[41]), .A0(A[41]), .A1(n15) );
  xor2 U418 ( .Y(SUM[40]), .A0(A[40]), .A1(n23) );
  xor2 U419 ( .Y(SUM[39]), .A0(A[39]), .A1(n27) );
  xor2 U420 ( .Y(SUM[38]), .A0(A[38]), .A1(n21) );
  xor2 U421 ( .Y(SUM[37]), .A0(A[37]), .A1(carry_37_) );
  xor2 U422 ( .Y(SUM[12]), .A0(B[12]), .A1(A[12]) );
  fadd1 U1_13 ( .S(n391), .CO(carry_14_), .A(A[13]), .B(B[13]), .CI(n13) );
  fadd1 U1_14 ( .S(n390), .CO(carry_15_), .A(A[14]), .B(B[14]), .CI(n41) );
  fadd1 U1_15 ( .S(n389), .CO(carry_16_), .A(A[15]), .B(B[15]), .CI(n40) );
  fadd1 U1_16 ( .S(n388), .CO(carry_17_), .A(A[16]), .B(B[16]), .CI(n39) );
  fadd1 U1_17 ( .S(n387), .CO(carry_18_), .A(A[17]), .B(B[17]), .CI(n38) );
  fadd1 U1_18 ( .S(n386), .CO(carry_19_), .A(A[18]), .B(B[18]), .CI(n37) );
  fadd1 U1_19 ( .S(n385), .CO(carry_20_), .A(A[19]), .B(B[19]), .CI(n36) );
  fadd1 U1_20 ( .S(n384), .CO(carry_21_), .A(A[20]), .B(B[20]), .CI(n35) );
  fadd1 U1_21 ( .S(n383), .CO(carry_22_), .A(A[21]), .B(B[21]), .CI(n34) );
  fadd1 U1_22 ( .S(n382), .CO(carry_23_), .A(A[22]), .B(B[22]), .CI(n33) );
  fadd1 U1_23 ( .S(n381), .CO(carry_24_), .A(A[23]), .B(B[23]), .CI(n32) );
endmodule


module mul_24_DW01_add_48_1 ( A, B, CI, SUM, CO );
  input [47:0] A;
  input [47:0] B;
  output [47:0] SUM;
  input CI;
  output CO;
  wire   carry_24_, carry_23_, carry_22_, carry_21_, carry_20_, carry_19_,
         carry_18_, carry_17_, carry_16_, carry_15_, carry_14_, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_, B_1_,
         B_0_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n26, n27, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325;
  assign SUM[11] = B_11_;
  assign B_11_ = B[11];
  assign SUM[10] = B_10_;
  assign B_10_ = B[10];
  assign SUM[9] = B_9_;
  assign B_9_ = B[9];
  assign SUM[8] = B_8_;
  assign B_8_ = B[8];
  assign SUM[7] = B_7_;
  assign B_7_ = B[7];
  assign SUM[6] = B_6_;
  assign B_6_ = B[6];
  assign SUM[5] = B_5_;
  assign B_5_ = B[5];
  assign SUM[4] = B_4_;
  assign B_4_ = B[4];
  assign SUM[3] = B_3_;
  assign B_3_ = B[3];
  assign SUM[2] = B_2_;
  assign B_2_ = B[2];
  assign SUM[1] = B_1_;
  assign B_1_ = B[1];
  assign SUM[0] = B_0_;
  assign B_0_ = B[0];

  nand02 U4 ( .Y(n1), .A0(n14), .A1(A[34]) );
  inv02 U5 ( .Y(n2), .A(n1) );
  nand02 U6 ( .Y(n3), .A0(n10), .A1(A[31]) );
  inv02 U7 ( .Y(n4), .A(n3) );
  nand02 U8 ( .Y(n5), .A0(n16), .A1(A[27]) );
  inv02 U9 ( .Y(n6), .A(n5) );
  nand02 U10 ( .Y(n7), .A0(carry_24_), .A1(A[24]) );
  inv02 U11 ( .Y(n8), .A(n7) );
  nand02 U12 ( .Y(n9), .A0(n20), .A1(A[30]) );
  inv02 U13 ( .Y(n10), .A(n9) );
  nand02 U14 ( .Y(n11), .A0(n8), .A1(A[25]) );
  inv02 U15 ( .Y(n12), .A(n11) );
  nand02 U16 ( .Y(n13), .A0(n22), .A1(A[33]) );
  inv02 U17 ( .Y(n14), .A(n13) );
  nand02 U18 ( .Y(n15), .A0(n12), .A1(A[26]) );
  inv02 U19 ( .Y(n16), .A(n15) );
  nand02 U20 ( .Y(n17), .A0(n6), .A1(A[28]) );
  inv02 U21 ( .Y(n18), .A(n17) );
  nand02 U22 ( .Y(n19), .A0(n18), .A1(A[29]) );
  inv02 U23 ( .Y(n20), .A(n19) );
  nand02 U24 ( .Y(n21), .A0(n4), .A1(A[32]) );
  inv02 U25 ( .Y(n22), .A(n21) );
  nand02 U26 ( .Y(n23), .A0(n2), .A1(A[35]) );
  inv02 U27 ( .Y(SUM[36]), .A(n23) );
  buf02 U28 ( .Y(SUM[12]), .A(n338) );
  nand02 U29 ( .Y(n26), .A0(A[12]), .A1(B[12]) );
  inv02 U30 ( .Y(n27), .A(n26) );
  buf02 U31 ( .Y(SUM[24]), .A(n337) );
  buf02 U32 ( .Y(SUM[29]), .A(n332) );
  buf02 U33 ( .Y(SUM[33]), .A(n328) );
  buf02 U34 ( .Y(SUM[32]), .A(n329) );
  buf02 U35 ( .Y(SUM[30]), .A(n331) );
  buf02 U36 ( .Y(SUM[25]), .A(n336) );
  buf02 U37 ( .Y(SUM[34]), .A(n327) );
  buf02 U38 ( .Y(SUM[35]), .A(n326) );
  buf02 U39 ( .Y(SUM[27]), .A(n334) );
  buf02 U40 ( .Y(SUM[31]), .A(n330) );
  buf02 U41 ( .Y(SUM[28]), .A(n333) );
  buf02 U42 ( .Y(SUM[26]), .A(n335) );
  inv02 U43 ( .Y(SUM[23]), .A(n40) );
  inv02 U44 ( .Y(carry_24_), .A(n41) );
  inv02 U45 ( .Y(n42), .A(B[23]) );
  inv02 U46 ( .Y(n43), .A(A[23]) );
  inv02 U47 ( .Y(n44), .A(carry_23_) );
  nor02 U48 ( .Y(n45), .A0(n42), .A1(n46) );
  nor02 U49 ( .Y(n47), .A0(n43), .A1(n48) );
  nor02 U50 ( .Y(n49), .A0(n44), .A1(n50) );
  nor02 U51 ( .Y(n51), .A0(n44), .A1(n52) );
  nor02 U52 ( .Y(n40), .A0(n53), .A1(n54) );
  nor02 U53 ( .Y(n55), .A0(n43), .A1(n44) );
  nor02 U54 ( .Y(n56), .A0(n42), .A1(n44) );
  nor02 U55 ( .Y(n57), .A0(n42), .A1(n43) );
  nor02 U56 ( .Y(n41), .A0(n57), .A1(n58) );
  nor02 U57 ( .Y(n59), .A0(A[23]), .A1(carry_23_) );
  inv01 U58 ( .Y(n46), .A(n59) );
  nor02 U59 ( .Y(n60), .A0(B[23]), .A1(carry_23_) );
  inv01 U60 ( .Y(n48), .A(n60) );
  nor02 U61 ( .Y(n61), .A0(B[23]), .A1(A[23]) );
  inv01 U62 ( .Y(n50), .A(n61) );
  nor02 U63 ( .Y(n62), .A0(n42), .A1(n43) );
  inv01 U64 ( .Y(n52), .A(n62) );
  nor02 U65 ( .Y(n63), .A0(n45), .A1(n47) );
  inv01 U66 ( .Y(n53), .A(n63) );
  nor02 U67 ( .Y(n64), .A0(n49), .A1(n51) );
  inv01 U68 ( .Y(n54), .A(n64) );
  nor02 U69 ( .Y(n65), .A0(n55), .A1(n56) );
  inv01 U70 ( .Y(n58), .A(n65) );
  inv02 U71 ( .Y(SUM[22]), .A(n66) );
  inv02 U72 ( .Y(carry_23_), .A(n67) );
  inv02 U73 ( .Y(n68), .A(B[22]) );
  inv02 U74 ( .Y(n69), .A(A[22]) );
  inv02 U75 ( .Y(n70), .A(carry_22_) );
  nor02 U76 ( .Y(n71), .A0(n68), .A1(n72) );
  nor02 U77 ( .Y(n73), .A0(n69), .A1(n74) );
  nor02 U78 ( .Y(n75), .A0(n70), .A1(n76) );
  nor02 U79 ( .Y(n77), .A0(n70), .A1(n78) );
  nor02 U80 ( .Y(n66), .A0(n79), .A1(n80) );
  nor02 U81 ( .Y(n81), .A0(n69), .A1(n70) );
  nor02 U82 ( .Y(n82), .A0(n68), .A1(n70) );
  nor02 U83 ( .Y(n83), .A0(n68), .A1(n69) );
  nor02 U84 ( .Y(n67), .A0(n83), .A1(n84) );
  nor02 U85 ( .Y(n85), .A0(A[22]), .A1(carry_22_) );
  inv01 U86 ( .Y(n72), .A(n85) );
  nor02 U87 ( .Y(n86), .A0(B[22]), .A1(carry_22_) );
  inv01 U88 ( .Y(n74), .A(n86) );
  nor02 U89 ( .Y(n87), .A0(B[22]), .A1(A[22]) );
  inv01 U90 ( .Y(n76), .A(n87) );
  nor02 U91 ( .Y(n88), .A0(n68), .A1(n69) );
  inv01 U92 ( .Y(n78), .A(n88) );
  nor02 U93 ( .Y(n89), .A0(n71), .A1(n73) );
  inv01 U94 ( .Y(n79), .A(n89) );
  nor02 U95 ( .Y(n90), .A0(n75), .A1(n77) );
  inv01 U96 ( .Y(n80), .A(n90) );
  nor02 U97 ( .Y(n91), .A0(n81), .A1(n82) );
  inv01 U98 ( .Y(n84), .A(n91) );
  inv02 U99 ( .Y(SUM[21]), .A(n92) );
  inv02 U100 ( .Y(carry_22_), .A(n93) );
  inv02 U101 ( .Y(n94), .A(B[21]) );
  inv02 U102 ( .Y(n95), .A(A[21]) );
  inv02 U103 ( .Y(n96), .A(carry_21_) );
  nor02 U104 ( .Y(n97), .A0(n94), .A1(n98) );
  nor02 U105 ( .Y(n99), .A0(n95), .A1(n100) );
  nor02 U106 ( .Y(n101), .A0(n96), .A1(n102) );
  nor02 U107 ( .Y(n103), .A0(n96), .A1(n104) );
  nor02 U108 ( .Y(n92), .A0(n105), .A1(n106) );
  nor02 U109 ( .Y(n107), .A0(n95), .A1(n96) );
  nor02 U110 ( .Y(n108), .A0(n94), .A1(n96) );
  nor02 U111 ( .Y(n109), .A0(n94), .A1(n95) );
  nor02 U112 ( .Y(n93), .A0(n109), .A1(n110) );
  nor02 U113 ( .Y(n111), .A0(A[21]), .A1(carry_21_) );
  inv01 U114 ( .Y(n98), .A(n111) );
  nor02 U115 ( .Y(n112), .A0(B[21]), .A1(carry_21_) );
  inv01 U116 ( .Y(n100), .A(n112) );
  nor02 U117 ( .Y(n113), .A0(B[21]), .A1(A[21]) );
  inv01 U118 ( .Y(n102), .A(n113) );
  nor02 U119 ( .Y(n114), .A0(n94), .A1(n95) );
  inv01 U120 ( .Y(n104), .A(n114) );
  nor02 U121 ( .Y(n115), .A0(n97), .A1(n99) );
  inv01 U122 ( .Y(n105), .A(n115) );
  nor02 U123 ( .Y(n116), .A0(n101), .A1(n103) );
  inv01 U124 ( .Y(n106), .A(n116) );
  nor02 U125 ( .Y(n117), .A0(n107), .A1(n108) );
  inv01 U126 ( .Y(n110), .A(n117) );
  inv02 U127 ( .Y(SUM[20]), .A(n118) );
  inv02 U128 ( .Y(carry_21_), .A(n119) );
  inv02 U129 ( .Y(n120), .A(B[20]) );
  inv02 U130 ( .Y(n121), .A(A[20]) );
  inv02 U131 ( .Y(n122), .A(carry_20_) );
  nor02 U132 ( .Y(n123), .A0(n120), .A1(n124) );
  nor02 U133 ( .Y(n125), .A0(n121), .A1(n126) );
  nor02 U134 ( .Y(n127), .A0(n122), .A1(n128) );
  nor02 U135 ( .Y(n129), .A0(n122), .A1(n130) );
  nor02 U136 ( .Y(n118), .A0(n131), .A1(n132) );
  nor02 U137 ( .Y(n133), .A0(n121), .A1(n122) );
  nor02 U138 ( .Y(n134), .A0(n120), .A1(n122) );
  nor02 U139 ( .Y(n135), .A0(n120), .A1(n121) );
  nor02 U140 ( .Y(n119), .A0(n135), .A1(n136) );
  nor02 U141 ( .Y(n137), .A0(A[20]), .A1(carry_20_) );
  inv01 U142 ( .Y(n124), .A(n137) );
  nor02 U143 ( .Y(n138), .A0(B[20]), .A1(carry_20_) );
  inv01 U144 ( .Y(n126), .A(n138) );
  nor02 U145 ( .Y(n139), .A0(B[20]), .A1(A[20]) );
  inv01 U146 ( .Y(n128), .A(n139) );
  nor02 U147 ( .Y(n140), .A0(n120), .A1(n121) );
  inv01 U148 ( .Y(n130), .A(n140) );
  nor02 U149 ( .Y(n141), .A0(n123), .A1(n125) );
  inv01 U150 ( .Y(n131), .A(n141) );
  nor02 U151 ( .Y(n142), .A0(n127), .A1(n129) );
  inv01 U152 ( .Y(n132), .A(n142) );
  nor02 U153 ( .Y(n143), .A0(n133), .A1(n134) );
  inv01 U154 ( .Y(n136), .A(n143) );
  inv02 U155 ( .Y(SUM[19]), .A(n144) );
  inv02 U156 ( .Y(carry_20_), .A(n145) );
  inv02 U157 ( .Y(n146), .A(B[19]) );
  inv02 U158 ( .Y(n147), .A(A[19]) );
  inv02 U159 ( .Y(n148), .A(carry_19_) );
  nor02 U160 ( .Y(n149), .A0(n146), .A1(n150) );
  nor02 U161 ( .Y(n151), .A0(n147), .A1(n152) );
  nor02 U162 ( .Y(n153), .A0(n148), .A1(n154) );
  nor02 U163 ( .Y(n155), .A0(n148), .A1(n156) );
  nor02 U164 ( .Y(n144), .A0(n157), .A1(n158) );
  nor02 U165 ( .Y(n159), .A0(n147), .A1(n148) );
  nor02 U166 ( .Y(n160), .A0(n146), .A1(n148) );
  nor02 U167 ( .Y(n161), .A0(n146), .A1(n147) );
  nor02 U168 ( .Y(n145), .A0(n161), .A1(n162) );
  nor02 U169 ( .Y(n163), .A0(A[19]), .A1(carry_19_) );
  inv01 U170 ( .Y(n150), .A(n163) );
  nor02 U171 ( .Y(n164), .A0(B[19]), .A1(carry_19_) );
  inv01 U172 ( .Y(n152), .A(n164) );
  nor02 U173 ( .Y(n165), .A0(B[19]), .A1(A[19]) );
  inv01 U174 ( .Y(n154), .A(n165) );
  nor02 U175 ( .Y(n166), .A0(n146), .A1(n147) );
  inv01 U176 ( .Y(n156), .A(n166) );
  nor02 U177 ( .Y(n167), .A0(n149), .A1(n151) );
  inv01 U178 ( .Y(n157), .A(n167) );
  nor02 U179 ( .Y(n168), .A0(n153), .A1(n155) );
  inv01 U180 ( .Y(n158), .A(n168) );
  nor02 U181 ( .Y(n169), .A0(n159), .A1(n160) );
  inv01 U182 ( .Y(n162), .A(n169) );
  inv02 U183 ( .Y(SUM[18]), .A(n170) );
  inv02 U184 ( .Y(carry_19_), .A(n171) );
  inv02 U185 ( .Y(n172), .A(B[18]) );
  inv02 U186 ( .Y(n173), .A(A[18]) );
  inv02 U187 ( .Y(n174), .A(carry_18_) );
  nor02 U188 ( .Y(n175), .A0(n172), .A1(n176) );
  nor02 U189 ( .Y(n177), .A0(n173), .A1(n178) );
  nor02 U190 ( .Y(n179), .A0(n174), .A1(n180) );
  nor02 U191 ( .Y(n181), .A0(n174), .A1(n182) );
  nor02 U192 ( .Y(n170), .A0(n183), .A1(n184) );
  nor02 U193 ( .Y(n185), .A0(n173), .A1(n174) );
  nor02 U194 ( .Y(n186), .A0(n172), .A1(n174) );
  nor02 U195 ( .Y(n187), .A0(n172), .A1(n173) );
  nor02 U196 ( .Y(n171), .A0(n187), .A1(n188) );
  nor02 U197 ( .Y(n189), .A0(A[18]), .A1(carry_18_) );
  inv01 U198 ( .Y(n176), .A(n189) );
  nor02 U199 ( .Y(n190), .A0(B[18]), .A1(carry_18_) );
  inv01 U200 ( .Y(n178), .A(n190) );
  nor02 U201 ( .Y(n191), .A0(B[18]), .A1(A[18]) );
  inv01 U202 ( .Y(n180), .A(n191) );
  nor02 U203 ( .Y(n192), .A0(n172), .A1(n173) );
  inv01 U204 ( .Y(n182), .A(n192) );
  nor02 U205 ( .Y(n193), .A0(n175), .A1(n177) );
  inv01 U206 ( .Y(n183), .A(n193) );
  nor02 U207 ( .Y(n194), .A0(n179), .A1(n181) );
  inv01 U208 ( .Y(n184), .A(n194) );
  nor02 U209 ( .Y(n195), .A0(n185), .A1(n186) );
  inv01 U210 ( .Y(n188), .A(n195) );
  inv02 U211 ( .Y(SUM[17]), .A(n196) );
  inv02 U212 ( .Y(carry_18_), .A(n197) );
  inv02 U213 ( .Y(n198), .A(B[17]) );
  inv02 U214 ( .Y(n199), .A(A[17]) );
  inv02 U215 ( .Y(n200), .A(carry_17_) );
  nor02 U216 ( .Y(n201), .A0(n198), .A1(n202) );
  nor02 U217 ( .Y(n203), .A0(n199), .A1(n204) );
  nor02 U218 ( .Y(n205), .A0(n200), .A1(n206) );
  nor02 U219 ( .Y(n207), .A0(n200), .A1(n208) );
  nor02 U220 ( .Y(n196), .A0(n209), .A1(n210) );
  nor02 U221 ( .Y(n211), .A0(n199), .A1(n200) );
  nor02 U222 ( .Y(n212), .A0(n198), .A1(n200) );
  nor02 U223 ( .Y(n213), .A0(n198), .A1(n199) );
  nor02 U224 ( .Y(n197), .A0(n213), .A1(n214) );
  nor02 U225 ( .Y(n215), .A0(A[17]), .A1(carry_17_) );
  inv01 U226 ( .Y(n202), .A(n215) );
  nor02 U227 ( .Y(n216), .A0(B[17]), .A1(carry_17_) );
  inv01 U228 ( .Y(n204), .A(n216) );
  nor02 U229 ( .Y(n217), .A0(B[17]), .A1(A[17]) );
  inv01 U230 ( .Y(n206), .A(n217) );
  nor02 U231 ( .Y(n218), .A0(n198), .A1(n199) );
  inv01 U232 ( .Y(n208), .A(n218) );
  nor02 U233 ( .Y(n219), .A0(n201), .A1(n203) );
  inv01 U234 ( .Y(n209), .A(n219) );
  nor02 U235 ( .Y(n220), .A0(n205), .A1(n207) );
  inv01 U236 ( .Y(n210), .A(n220) );
  nor02 U237 ( .Y(n221), .A0(n211), .A1(n212) );
  inv01 U238 ( .Y(n214), .A(n221) );
  inv02 U239 ( .Y(SUM[16]), .A(n222) );
  inv02 U240 ( .Y(carry_17_), .A(n223) );
  inv02 U241 ( .Y(n224), .A(B[16]) );
  inv02 U242 ( .Y(n225), .A(A[16]) );
  inv02 U243 ( .Y(n226), .A(carry_16_) );
  nor02 U244 ( .Y(n227), .A0(n224), .A1(n228) );
  nor02 U245 ( .Y(n229), .A0(n225), .A1(n230) );
  nor02 U246 ( .Y(n231), .A0(n226), .A1(n232) );
  nor02 U247 ( .Y(n233), .A0(n226), .A1(n234) );
  nor02 U248 ( .Y(n222), .A0(n235), .A1(n236) );
  nor02 U249 ( .Y(n237), .A0(n225), .A1(n226) );
  nor02 U250 ( .Y(n238), .A0(n224), .A1(n226) );
  nor02 U251 ( .Y(n239), .A0(n224), .A1(n225) );
  nor02 U252 ( .Y(n223), .A0(n239), .A1(n240) );
  nor02 U253 ( .Y(n241), .A0(A[16]), .A1(carry_16_) );
  inv01 U254 ( .Y(n228), .A(n241) );
  nor02 U255 ( .Y(n242), .A0(B[16]), .A1(carry_16_) );
  inv01 U256 ( .Y(n230), .A(n242) );
  nor02 U257 ( .Y(n243), .A0(B[16]), .A1(A[16]) );
  inv01 U258 ( .Y(n232), .A(n243) );
  nor02 U259 ( .Y(n244), .A0(n224), .A1(n225) );
  inv01 U260 ( .Y(n234), .A(n244) );
  nor02 U261 ( .Y(n245), .A0(n227), .A1(n229) );
  inv01 U262 ( .Y(n235), .A(n245) );
  nor02 U263 ( .Y(n246), .A0(n231), .A1(n233) );
  inv01 U264 ( .Y(n236), .A(n246) );
  nor02 U265 ( .Y(n247), .A0(n237), .A1(n238) );
  inv01 U266 ( .Y(n240), .A(n247) );
  inv02 U267 ( .Y(SUM[15]), .A(n248) );
  inv02 U268 ( .Y(carry_16_), .A(n249) );
  inv02 U269 ( .Y(n250), .A(B[15]) );
  inv02 U270 ( .Y(n251), .A(A[15]) );
  inv02 U271 ( .Y(n252), .A(carry_15_) );
  nor02 U272 ( .Y(n253), .A0(n250), .A1(n254) );
  nor02 U273 ( .Y(n255), .A0(n251), .A1(n256) );
  nor02 U274 ( .Y(n257), .A0(n252), .A1(n258) );
  nor02 U275 ( .Y(n259), .A0(n252), .A1(n260) );
  nor02 U276 ( .Y(n248), .A0(n261), .A1(n262) );
  nor02 U277 ( .Y(n263), .A0(n251), .A1(n252) );
  nor02 U278 ( .Y(n264), .A0(n250), .A1(n252) );
  nor02 U279 ( .Y(n265), .A0(n250), .A1(n251) );
  nor02 U280 ( .Y(n249), .A0(n265), .A1(n266) );
  nor02 U281 ( .Y(n267), .A0(A[15]), .A1(carry_15_) );
  inv01 U282 ( .Y(n254), .A(n267) );
  nor02 U283 ( .Y(n268), .A0(B[15]), .A1(carry_15_) );
  inv01 U284 ( .Y(n256), .A(n268) );
  nor02 U285 ( .Y(n269), .A0(B[15]), .A1(A[15]) );
  inv01 U286 ( .Y(n258), .A(n269) );
  nor02 U287 ( .Y(n270), .A0(n250), .A1(n251) );
  inv01 U288 ( .Y(n260), .A(n270) );
  nor02 U289 ( .Y(n271), .A0(n253), .A1(n255) );
  inv01 U290 ( .Y(n261), .A(n271) );
  nor02 U291 ( .Y(n272), .A0(n257), .A1(n259) );
  inv01 U292 ( .Y(n262), .A(n272) );
  nor02 U293 ( .Y(n273), .A0(n263), .A1(n264) );
  inv01 U294 ( .Y(n266), .A(n273) );
  inv02 U295 ( .Y(SUM[14]), .A(n274) );
  inv02 U296 ( .Y(carry_15_), .A(n275) );
  inv02 U297 ( .Y(n276), .A(B[14]) );
  inv02 U298 ( .Y(n277), .A(A[14]) );
  inv02 U299 ( .Y(n278), .A(carry_14_) );
  nor02 U300 ( .Y(n279), .A0(n276), .A1(n280) );
  nor02 U301 ( .Y(n281), .A0(n277), .A1(n282) );
  nor02 U302 ( .Y(n283), .A0(n278), .A1(n284) );
  nor02 U303 ( .Y(n285), .A0(n278), .A1(n286) );
  nor02 U304 ( .Y(n274), .A0(n287), .A1(n288) );
  nor02 U305 ( .Y(n289), .A0(n277), .A1(n278) );
  nor02 U306 ( .Y(n290), .A0(n276), .A1(n278) );
  nor02 U307 ( .Y(n291), .A0(n276), .A1(n277) );
  nor02 U308 ( .Y(n275), .A0(n291), .A1(n292) );
  nor02 U309 ( .Y(n293), .A0(A[14]), .A1(carry_14_) );
  inv01 U310 ( .Y(n280), .A(n293) );
  nor02 U311 ( .Y(n294), .A0(B[14]), .A1(carry_14_) );
  inv01 U312 ( .Y(n282), .A(n294) );
  nor02 U313 ( .Y(n295), .A0(B[14]), .A1(A[14]) );
  inv01 U314 ( .Y(n284), .A(n295) );
  nor02 U315 ( .Y(n296), .A0(n276), .A1(n277) );
  inv01 U316 ( .Y(n286), .A(n296) );
  nor02 U317 ( .Y(n297), .A0(n279), .A1(n281) );
  inv01 U318 ( .Y(n287), .A(n297) );
  nor02 U319 ( .Y(n298), .A0(n283), .A1(n285) );
  inv01 U320 ( .Y(n288), .A(n298) );
  nor02 U321 ( .Y(n299), .A0(n289), .A1(n290) );
  inv01 U322 ( .Y(n292), .A(n299) );
  inv02 U323 ( .Y(SUM[13]), .A(n300) );
  inv02 U324 ( .Y(carry_14_), .A(n301) );
  inv02 U325 ( .Y(n302), .A(B[13]) );
  inv02 U326 ( .Y(n303), .A(A[13]) );
  inv02 U327 ( .Y(n304), .A(n27) );
  nor02 U328 ( .Y(n305), .A0(n302), .A1(n306) );
  nor02 U329 ( .Y(n307), .A0(n303), .A1(n308) );
  nor02 U330 ( .Y(n309), .A0(n304), .A1(n310) );
  nor02 U331 ( .Y(n311), .A0(n304), .A1(n312) );
  nor02 U332 ( .Y(n300), .A0(n313), .A1(n314) );
  nor02 U333 ( .Y(n315), .A0(n303), .A1(n304) );
  nor02 U334 ( .Y(n316), .A0(n302), .A1(n304) );
  nor02 U335 ( .Y(n317), .A0(n302), .A1(n303) );
  nor02 U336 ( .Y(n301), .A0(n317), .A1(n318) );
  nor02 U337 ( .Y(n319), .A0(A[13]), .A1(n27) );
  inv01 U338 ( .Y(n306), .A(n319) );
  nor02 U339 ( .Y(n320), .A0(B[13]), .A1(n27) );
  inv01 U340 ( .Y(n308), .A(n320) );
  nor02 U341 ( .Y(n321), .A0(B[13]), .A1(A[13]) );
  inv01 U342 ( .Y(n310), .A(n321) );
  nor02 U343 ( .Y(n322), .A0(n302), .A1(n303) );
  inv01 U344 ( .Y(n312), .A(n322) );
  nor02 U345 ( .Y(n323), .A0(n305), .A1(n307) );
  inv01 U346 ( .Y(n313), .A(n323) );
  nor02 U347 ( .Y(n324), .A0(n309), .A1(n311) );
  inv01 U348 ( .Y(n314), .A(n324) );
  nor02 U349 ( .Y(n325), .A0(n315), .A1(n316) );
  inv01 U350 ( .Y(n318), .A(n325) );
  xor2 U351 ( .Y(n326), .A0(A[35]), .A1(n2) );
  xor2 U352 ( .Y(n327), .A0(A[34]), .A1(n14) );
  xor2 U353 ( .Y(n328), .A0(A[33]), .A1(n22) );
  xor2 U354 ( .Y(n329), .A0(A[32]), .A1(n4) );
  xor2 U355 ( .Y(n330), .A0(A[31]), .A1(n10) );
  xor2 U356 ( .Y(n331), .A0(A[30]), .A1(n20) );
  xor2 U357 ( .Y(n332), .A0(A[29]), .A1(n18) );
  xor2 U358 ( .Y(n333), .A0(A[28]), .A1(n6) );
  xor2 U359 ( .Y(n334), .A0(A[27]), .A1(n16) );
  xor2 U360 ( .Y(n335), .A0(A[26]), .A1(n12) );
  xor2 U361 ( .Y(n336), .A0(A[25]), .A1(n8) );
  xor2 U362 ( .Y(n337), .A0(A[24]), .A1(carry_24_) );
  xor2 U363 ( .Y(n338), .A0(B[12]), .A1(A[12]) );
endmodule


module mul_24_DW01_add_48_0 ( A, B, CI, SUM, CO );
  input [47:0] A;
  input [47:0] B;
  output [47:0] SUM;
  input CI;
  output CO;
  wire   carry_47_, carry_36_, carry_35_, carry_34_, carry_33_, carry_32_,
         carry_31_, carry_30_, carry_29_, carry_28_, carry_27_, carry_26_,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_,
         B_14_, B_13_, B_12_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n25, n27,
         n29, n31, n34, n36, n38, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328;
  assign SUM[23] = B_23_;
  assign B_23_ = B[23];
  assign SUM[22] = B_22_;
  assign B_22_ = B[22];
  assign SUM[21] = B_21_;
  assign B_21_ = B[21];
  assign SUM[20] = B_20_;
  assign B_20_ = B[20];
  assign SUM[19] = B_19_;
  assign B_19_ = B[19];
  assign SUM[18] = B_18_;
  assign B_18_ = B[18];
  assign SUM[17] = B_17_;
  assign B_17_ = B[17];
  assign SUM[16] = B_16_;
  assign B_16_ = B[16];
  assign SUM[15] = B_15_;
  assign B_15_ = B[15];
  assign SUM[14] = B_14_;
  assign B_14_ = B[14];
  assign SUM[13] = B_13_;
  assign B_13_ = B[13];
  assign SUM[12] = B_12_;
  assign B_12_ = B[12];

  nand02 U4 ( .Y(n1), .A0(A[24]), .A1(B[24]) );
  inv02 U5 ( .Y(n2), .A(n1) );
  nand02 U6 ( .Y(n3), .A0(n14), .A1(A[42]) );
  inv02 U7 ( .Y(n4), .A(n3) );
  nand02 U8 ( .Y(n5), .A0(n16), .A1(A[44]) );
  inv02 U9 ( .Y(n6), .A(n5) );
  nand02 U10 ( .Y(n7), .A0(carry_36_), .A1(A[36]) );
  inv02 U11 ( .Y(n8), .A(n7) );
  nand02 U12 ( .Y(n9), .A0(n20), .A1(A[39]) );
  inv02 U13 ( .Y(n10), .A(n9) );
  nand02 U14 ( .Y(n11), .A0(n10), .A1(A[40]) );
  inv02 U15 ( .Y(n12), .A(n11) );
  nand02 U16 ( .Y(n13), .A0(n12), .A1(A[41]) );
  inv02 U17 ( .Y(n14), .A(n13) );
  nand02 U18 ( .Y(n15), .A0(n4), .A1(A[43]) );
  inv02 U19 ( .Y(n16), .A(n15) );
  nand02 U20 ( .Y(n17), .A0(n6), .A1(A[45]) );
  inv02 U21 ( .Y(n18), .A(n17) );
  nand02 U22 ( .Y(n19), .A0(n22), .A1(A[38]) );
  inv02 U23 ( .Y(n20), .A(n19) );
  nand02 U24 ( .Y(n21), .A0(n8), .A1(A[37]) );
  inv02 U25 ( .Y(n22), .A(n21) );
  inv01 U26 ( .Y(n23), .A(n330) );
  inv02 U27 ( .Y(SUM[45]), .A(n23) );
  inv01 U28 ( .Y(n25), .A(n336) );
  inv02 U29 ( .Y(SUM[39]), .A(n25) );
  inv01 U30 ( .Y(n27), .A(n333) );
  inv02 U31 ( .Y(SUM[42]), .A(n27) );
  inv01 U32 ( .Y(n29), .A(n335) );
  inv02 U33 ( .Y(SUM[40]), .A(n29) );
  inv01 U34 ( .Y(n31), .A(n338) );
  inv02 U35 ( .Y(SUM[37]), .A(n31) );
  buf02 U36 ( .Y(SUM[46]), .A(n329) );
  inv01 U37 ( .Y(n34), .A(n332) );
  inv02 U38 ( .Y(SUM[43]), .A(n34) );
  inv01 U39 ( .Y(n36), .A(n334) );
  inv02 U40 ( .Y(SUM[41]), .A(n36) );
  inv01 U41 ( .Y(n38), .A(n337) );
  inv02 U42 ( .Y(SUM[38]), .A(n38) );
  buf02 U43 ( .Y(SUM[44]), .A(n331) );
  buf02 U44 ( .Y(SUM[36]), .A(n339) );
  buf02 U45 ( .Y(SUM[24]), .A(n340) );
  inv02 U46 ( .Y(SUM[34]), .A(n43) );
  inv02 U47 ( .Y(carry_35_), .A(n44) );
  inv02 U48 ( .Y(n45), .A(B[34]) );
  inv02 U49 ( .Y(n46), .A(A[34]) );
  inv02 U50 ( .Y(n47), .A(carry_34_) );
  nor02 U51 ( .Y(n48), .A0(n45), .A1(n49) );
  nor02 U52 ( .Y(n50), .A0(n46), .A1(n51) );
  nor02 U53 ( .Y(n52), .A0(n47), .A1(n53) );
  nor02 U54 ( .Y(n54), .A0(n47), .A1(n55) );
  nor02 U55 ( .Y(n43), .A0(n56), .A1(n57) );
  nor02 U56 ( .Y(n58), .A0(n46), .A1(n47) );
  nor02 U57 ( .Y(n59), .A0(n45), .A1(n47) );
  nor02 U58 ( .Y(n60), .A0(n45), .A1(n46) );
  nor02 U59 ( .Y(n44), .A0(n60), .A1(n61) );
  nor02 U60 ( .Y(n62), .A0(A[34]), .A1(carry_34_) );
  inv01 U61 ( .Y(n49), .A(n62) );
  nor02 U62 ( .Y(n63), .A0(B[34]), .A1(carry_34_) );
  inv01 U63 ( .Y(n51), .A(n63) );
  nor02 U64 ( .Y(n64), .A0(B[34]), .A1(A[34]) );
  inv01 U65 ( .Y(n53), .A(n64) );
  nor02 U66 ( .Y(n65), .A0(n45), .A1(n46) );
  inv01 U67 ( .Y(n55), .A(n65) );
  nor02 U68 ( .Y(n66), .A0(n48), .A1(n50) );
  inv01 U69 ( .Y(n56), .A(n66) );
  nor02 U70 ( .Y(n67), .A0(n52), .A1(n54) );
  inv01 U71 ( .Y(n57), .A(n67) );
  nor02 U72 ( .Y(n68), .A0(n58), .A1(n59) );
  inv01 U73 ( .Y(n61), .A(n68) );
  inv02 U74 ( .Y(SUM[35]), .A(n69) );
  inv02 U75 ( .Y(carry_36_), .A(n70) );
  inv02 U76 ( .Y(n71), .A(B[35]) );
  inv02 U77 ( .Y(n72), .A(A[35]) );
  inv02 U78 ( .Y(n73), .A(carry_35_) );
  nor02 U79 ( .Y(n74), .A0(n71), .A1(n75) );
  nor02 U80 ( .Y(n76), .A0(n72), .A1(n77) );
  nor02 U81 ( .Y(n78), .A0(n73), .A1(n79) );
  nor02 U82 ( .Y(n80), .A0(n73), .A1(n81) );
  nor02 U83 ( .Y(n69), .A0(n82), .A1(n83) );
  nor02 U84 ( .Y(n84), .A0(n72), .A1(n73) );
  nor02 U85 ( .Y(n85), .A0(n71), .A1(n73) );
  nor02 U86 ( .Y(n86), .A0(n71), .A1(n72) );
  nor02 U87 ( .Y(n70), .A0(n86), .A1(n87) );
  nor02 U88 ( .Y(n88), .A0(A[35]), .A1(carry_35_) );
  inv01 U89 ( .Y(n75), .A(n88) );
  nor02 U90 ( .Y(n89), .A0(B[35]), .A1(carry_35_) );
  inv01 U91 ( .Y(n77), .A(n89) );
  nor02 U92 ( .Y(n90), .A0(B[35]), .A1(A[35]) );
  inv01 U93 ( .Y(n79), .A(n90) );
  nor02 U94 ( .Y(n91), .A0(n71), .A1(n72) );
  inv01 U95 ( .Y(n81), .A(n91) );
  nor02 U96 ( .Y(n92), .A0(n74), .A1(n76) );
  inv01 U97 ( .Y(n82), .A(n92) );
  nor02 U98 ( .Y(n93), .A0(n78), .A1(n80) );
  inv01 U99 ( .Y(n83), .A(n93) );
  nor02 U100 ( .Y(n94), .A0(n84), .A1(n85) );
  inv01 U101 ( .Y(n87), .A(n94) );
  inv02 U102 ( .Y(SUM[33]), .A(n95) );
  inv02 U103 ( .Y(carry_34_), .A(n96) );
  inv02 U104 ( .Y(n97), .A(B[33]) );
  inv02 U105 ( .Y(n98), .A(A[33]) );
  inv02 U106 ( .Y(n99), .A(carry_33_) );
  nor02 U107 ( .Y(n100), .A0(n97), .A1(n101) );
  nor02 U108 ( .Y(n102), .A0(n98), .A1(n103) );
  nor02 U109 ( .Y(n104), .A0(n99), .A1(n105) );
  nor02 U110 ( .Y(n106), .A0(n99), .A1(n107) );
  nor02 U111 ( .Y(n95), .A0(n108), .A1(n109) );
  nor02 U112 ( .Y(n110), .A0(n98), .A1(n99) );
  nor02 U113 ( .Y(n111), .A0(n97), .A1(n99) );
  nor02 U114 ( .Y(n112), .A0(n97), .A1(n98) );
  nor02 U115 ( .Y(n96), .A0(n112), .A1(n113) );
  nor02 U116 ( .Y(n114), .A0(A[33]), .A1(carry_33_) );
  inv01 U117 ( .Y(n101), .A(n114) );
  nor02 U118 ( .Y(n115), .A0(B[33]), .A1(carry_33_) );
  inv01 U119 ( .Y(n103), .A(n115) );
  nor02 U120 ( .Y(n116), .A0(B[33]), .A1(A[33]) );
  inv01 U121 ( .Y(n105), .A(n116) );
  nor02 U122 ( .Y(n117), .A0(n97), .A1(n98) );
  inv01 U123 ( .Y(n107), .A(n117) );
  nor02 U124 ( .Y(n118), .A0(n100), .A1(n102) );
  inv01 U125 ( .Y(n108), .A(n118) );
  nor02 U126 ( .Y(n119), .A0(n104), .A1(n106) );
  inv01 U127 ( .Y(n109), .A(n119) );
  nor02 U128 ( .Y(n120), .A0(n110), .A1(n111) );
  inv01 U129 ( .Y(n113), .A(n120) );
  inv02 U130 ( .Y(SUM[32]), .A(n121) );
  inv02 U131 ( .Y(carry_33_), .A(n122) );
  inv02 U132 ( .Y(n123), .A(B[32]) );
  inv02 U133 ( .Y(n124), .A(A[32]) );
  inv02 U134 ( .Y(n125), .A(carry_32_) );
  nor02 U135 ( .Y(n126), .A0(n123), .A1(n127) );
  nor02 U136 ( .Y(n128), .A0(n124), .A1(n129) );
  nor02 U137 ( .Y(n130), .A0(n125), .A1(n131) );
  nor02 U138 ( .Y(n132), .A0(n125), .A1(n133) );
  nor02 U139 ( .Y(n121), .A0(n134), .A1(n135) );
  nor02 U140 ( .Y(n136), .A0(n124), .A1(n125) );
  nor02 U141 ( .Y(n137), .A0(n123), .A1(n125) );
  nor02 U142 ( .Y(n138), .A0(n123), .A1(n124) );
  nor02 U143 ( .Y(n122), .A0(n138), .A1(n139) );
  nor02 U144 ( .Y(n140), .A0(A[32]), .A1(carry_32_) );
  inv01 U145 ( .Y(n127), .A(n140) );
  nor02 U146 ( .Y(n141), .A0(B[32]), .A1(carry_32_) );
  inv01 U147 ( .Y(n129), .A(n141) );
  nor02 U148 ( .Y(n142), .A0(B[32]), .A1(A[32]) );
  inv01 U149 ( .Y(n131), .A(n142) );
  nor02 U150 ( .Y(n143), .A0(n123), .A1(n124) );
  inv01 U151 ( .Y(n133), .A(n143) );
  nor02 U152 ( .Y(n144), .A0(n126), .A1(n128) );
  inv01 U153 ( .Y(n134), .A(n144) );
  nor02 U154 ( .Y(n145), .A0(n130), .A1(n132) );
  inv01 U155 ( .Y(n135), .A(n145) );
  nor02 U156 ( .Y(n146), .A0(n136), .A1(n137) );
  inv01 U157 ( .Y(n139), .A(n146) );
  inv02 U158 ( .Y(SUM[31]), .A(n147) );
  inv02 U159 ( .Y(carry_32_), .A(n148) );
  inv02 U160 ( .Y(n149), .A(B[31]) );
  inv02 U161 ( .Y(n150), .A(A[31]) );
  inv02 U162 ( .Y(n151), .A(carry_31_) );
  nor02 U163 ( .Y(n152), .A0(n149), .A1(n153) );
  nor02 U164 ( .Y(n154), .A0(n150), .A1(n155) );
  nor02 U165 ( .Y(n156), .A0(n151), .A1(n157) );
  nor02 U166 ( .Y(n158), .A0(n151), .A1(n159) );
  nor02 U167 ( .Y(n147), .A0(n160), .A1(n161) );
  nor02 U168 ( .Y(n162), .A0(n150), .A1(n151) );
  nor02 U169 ( .Y(n163), .A0(n149), .A1(n151) );
  nor02 U170 ( .Y(n164), .A0(n149), .A1(n150) );
  nor02 U171 ( .Y(n148), .A0(n164), .A1(n165) );
  nor02 U172 ( .Y(n166), .A0(A[31]), .A1(carry_31_) );
  inv01 U173 ( .Y(n153), .A(n166) );
  nor02 U174 ( .Y(n167), .A0(B[31]), .A1(carry_31_) );
  inv01 U175 ( .Y(n155), .A(n167) );
  nor02 U176 ( .Y(n168), .A0(B[31]), .A1(A[31]) );
  inv01 U177 ( .Y(n157), .A(n168) );
  nor02 U178 ( .Y(n169), .A0(n149), .A1(n150) );
  inv01 U179 ( .Y(n159), .A(n169) );
  nor02 U180 ( .Y(n170), .A0(n152), .A1(n154) );
  inv01 U181 ( .Y(n160), .A(n170) );
  nor02 U182 ( .Y(n171), .A0(n156), .A1(n158) );
  inv01 U183 ( .Y(n161), .A(n171) );
  nor02 U184 ( .Y(n172), .A0(n162), .A1(n163) );
  inv01 U185 ( .Y(n165), .A(n172) );
  inv02 U186 ( .Y(SUM[30]), .A(n173) );
  inv02 U187 ( .Y(carry_31_), .A(n174) );
  inv02 U188 ( .Y(n175), .A(B[30]) );
  inv02 U189 ( .Y(n176), .A(A[30]) );
  inv02 U190 ( .Y(n177), .A(carry_30_) );
  nor02 U191 ( .Y(n178), .A0(n175), .A1(n179) );
  nor02 U192 ( .Y(n180), .A0(n176), .A1(n181) );
  nor02 U193 ( .Y(n182), .A0(n177), .A1(n183) );
  nor02 U194 ( .Y(n184), .A0(n177), .A1(n185) );
  nor02 U195 ( .Y(n173), .A0(n186), .A1(n187) );
  nor02 U196 ( .Y(n188), .A0(n176), .A1(n177) );
  nor02 U197 ( .Y(n189), .A0(n175), .A1(n177) );
  nor02 U198 ( .Y(n190), .A0(n175), .A1(n176) );
  nor02 U199 ( .Y(n174), .A0(n190), .A1(n191) );
  nor02 U200 ( .Y(n192), .A0(A[30]), .A1(carry_30_) );
  inv01 U201 ( .Y(n179), .A(n192) );
  nor02 U202 ( .Y(n193), .A0(B[30]), .A1(carry_30_) );
  inv01 U203 ( .Y(n181), .A(n193) );
  nor02 U204 ( .Y(n194), .A0(B[30]), .A1(A[30]) );
  inv01 U205 ( .Y(n183), .A(n194) );
  nor02 U206 ( .Y(n195), .A0(n175), .A1(n176) );
  inv01 U207 ( .Y(n185), .A(n195) );
  nor02 U208 ( .Y(n196), .A0(n178), .A1(n180) );
  inv01 U209 ( .Y(n186), .A(n196) );
  nor02 U210 ( .Y(n197), .A0(n182), .A1(n184) );
  inv01 U211 ( .Y(n187), .A(n197) );
  nor02 U212 ( .Y(n198), .A0(n188), .A1(n189) );
  inv01 U213 ( .Y(n191), .A(n198) );
  inv02 U214 ( .Y(SUM[29]), .A(n199) );
  inv02 U215 ( .Y(carry_30_), .A(n200) );
  inv02 U216 ( .Y(n201), .A(B[29]) );
  inv02 U217 ( .Y(n202), .A(A[29]) );
  inv02 U218 ( .Y(n203), .A(carry_29_) );
  nor02 U219 ( .Y(n204), .A0(n201), .A1(n205) );
  nor02 U220 ( .Y(n206), .A0(n202), .A1(n207) );
  nor02 U221 ( .Y(n208), .A0(n203), .A1(n209) );
  nor02 U222 ( .Y(n210), .A0(n203), .A1(n211) );
  nor02 U223 ( .Y(n199), .A0(n212), .A1(n213) );
  nor02 U224 ( .Y(n214), .A0(n202), .A1(n203) );
  nor02 U225 ( .Y(n215), .A0(n201), .A1(n203) );
  nor02 U226 ( .Y(n216), .A0(n201), .A1(n202) );
  nor02 U227 ( .Y(n200), .A0(n216), .A1(n217) );
  nor02 U228 ( .Y(n218), .A0(A[29]), .A1(carry_29_) );
  inv01 U229 ( .Y(n205), .A(n218) );
  nor02 U230 ( .Y(n219), .A0(B[29]), .A1(carry_29_) );
  inv01 U231 ( .Y(n207), .A(n219) );
  nor02 U232 ( .Y(n220), .A0(B[29]), .A1(A[29]) );
  inv01 U233 ( .Y(n209), .A(n220) );
  nor02 U234 ( .Y(n221), .A0(n201), .A1(n202) );
  inv01 U235 ( .Y(n211), .A(n221) );
  nor02 U236 ( .Y(n222), .A0(n204), .A1(n206) );
  inv01 U237 ( .Y(n212), .A(n222) );
  nor02 U238 ( .Y(n223), .A0(n208), .A1(n210) );
  inv01 U239 ( .Y(n213), .A(n223) );
  nor02 U240 ( .Y(n224), .A0(n214), .A1(n215) );
  inv01 U241 ( .Y(n217), .A(n224) );
  inv02 U242 ( .Y(SUM[28]), .A(n225) );
  inv02 U243 ( .Y(carry_29_), .A(n226) );
  inv02 U244 ( .Y(n227), .A(B[28]) );
  inv02 U245 ( .Y(n228), .A(A[28]) );
  inv02 U246 ( .Y(n229), .A(carry_28_) );
  nor02 U247 ( .Y(n230), .A0(n227), .A1(n231) );
  nor02 U248 ( .Y(n232), .A0(n228), .A1(n233) );
  nor02 U249 ( .Y(n234), .A0(n229), .A1(n235) );
  nor02 U250 ( .Y(n236), .A0(n229), .A1(n237) );
  nor02 U251 ( .Y(n225), .A0(n238), .A1(n239) );
  nor02 U252 ( .Y(n240), .A0(n228), .A1(n229) );
  nor02 U253 ( .Y(n241), .A0(n227), .A1(n229) );
  nor02 U254 ( .Y(n242), .A0(n227), .A1(n228) );
  nor02 U255 ( .Y(n226), .A0(n242), .A1(n243) );
  nor02 U256 ( .Y(n244), .A0(A[28]), .A1(carry_28_) );
  inv01 U257 ( .Y(n231), .A(n244) );
  nor02 U258 ( .Y(n245), .A0(B[28]), .A1(carry_28_) );
  inv01 U259 ( .Y(n233), .A(n245) );
  nor02 U260 ( .Y(n246), .A0(B[28]), .A1(A[28]) );
  inv01 U261 ( .Y(n235), .A(n246) );
  nor02 U262 ( .Y(n247), .A0(n227), .A1(n228) );
  inv01 U263 ( .Y(n237), .A(n247) );
  nor02 U264 ( .Y(n248), .A0(n230), .A1(n232) );
  inv01 U265 ( .Y(n238), .A(n248) );
  nor02 U266 ( .Y(n249), .A0(n234), .A1(n236) );
  inv01 U267 ( .Y(n239), .A(n249) );
  nor02 U268 ( .Y(n250), .A0(n240), .A1(n241) );
  inv01 U269 ( .Y(n243), .A(n250) );
  inv02 U270 ( .Y(SUM[27]), .A(n251) );
  inv02 U271 ( .Y(carry_28_), .A(n252) );
  inv02 U272 ( .Y(n253), .A(B[27]) );
  inv02 U273 ( .Y(n254), .A(A[27]) );
  inv02 U274 ( .Y(n255), .A(carry_27_) );
  nor02 U275 ( .Y(n256), .A0(n253), .A1(n257) );
  nor02 U276 ( .Y(n258), .A0(n254), .A1(n259) );
  nor02 U277 ( .Y(n260), .A0(n255), .A1(n261) );
  nor02 U278 ( .Y(n262), .A0(n255), .A1(n263) );
  nor02 U279 ( .Y(n251), .A0(n264), .A1(n265) );
  nor02 U280 ( .Y(n266), .A0(n254), .A1(n255) );
  nor02 U281 ( .Y(n267), .A0(n253), .A1(n255) );
  nor02 U282 ( .Y(n268), .A0(n253), .A1(n254) );
  nor02 U283 ( .Y(n252), .A0(n268), .A1(n269) );
  nor02 U284 ( .Y(n270), .A0(A[27]), .A1(carry_27_) );
  inv01 U285 ( .Y(n257), .A(n270) );
  nor02 U286 ( .Y(n271), .A0(B[27]), .A1(carry_27_) );
  inv01 U287 ( .Y(n259), .A(n271) );
  nor02 U288 ( .Y(n272), .A0(B[27]), .A1(A[27]) );
  inv01 U289 ( .Y(n261), .A(n272) );
  nor02 U290 ( .Y(n273), .A0(n253), .A1(n254) );
  inv01 U291 ( .Y(n263), .A(n273) );
  nor02 U292 ( .Y(n274), .A0(n256), .A1(n258) );
  inv01 U293 ( .Y(n264), .A(n274) );
  nor02 U294 ( .Y(n275), .A0(n260), .A1(n262) );
  inv01 U295 ( .Y(n265), .A(n275) );
  nor02 U296 ( .Y(n276), .A0(n266), .A1(n267) );
  inv01 U297 ( .Y(n269), .A(n276) );
  inv02 U298 ( .Y(SUM[26]), .A(n277) );
  inv02 U299 ( .Y(carry_27_), .A(n278) );
  inv02 U300 ( .Y(n279), .A(B[26]) );
  inv02 U301 ( .Y(n280), .A(A[26]) );
  inv02 U302 ( .Y(n281), .A(carry_26_) );
  nor02 U303 ( .Y(n282), .A0(n279), .A1(n283) );
  nor02 U304 ( .Y(n284), .A0(n280), .A1(n285) );
  nor02 U305 ( .Y(n286), .A0(n281), .A1(n287) );
  nor02 U306 ( .Y(n288), .A0(n281), .A1(n289) );
  nor02 U307 ( .Y(n277), .A0(n290), .A1(n291) );
  nor02 U308 ( .Y(n292), .A0(n280), .A1(n281) );
  nor02 U309 ( .Y(n293), .A0(n279), .A1(n281) );
  nor02 U310 ( .Y(n294), .A0(n279), .A1(n280) );
  nor02 U311 ( .Y(n278), .A0(n294), .A1(n295) );
  nor02 U312 ( .Y(n296), .A0(A[26]), .A1(carry_26_) );
  inv01 U313 ( .Y(n283), .A(n296) );
  nor02 U314 ( .Y(n297), .A0(B[26]), .A1(carry_26_) );
  inv01 U315 ( .Y(n285), .A(n297) );
  nor02 U316 ( .Y(n298), .A0(B[26]), .A1(A[26]) );
  inv01 U317 ( .Y(n287), .A(n298) );
  nor02 U318 ( .Y(n299), .A0(n279), .A1(n280) );
  inv01 U319 ( .Y(n289), .A(n299) );
  nor02 U320 ( .Y(n300), .A0(n282), .A1(n284) );
  inv01 U321 ( .Y(n290), .A(n300) );
  nor02 U322 ( .Y(n301), .A0(n286), .A1(n288) );
  inv01 U323 ( .Y(n291), .A(n301) );
  nor02 U324 ( .Y(n302), .A0(n292), .A1(n293) );
  inv01 U325 ( .Y(n295), .A(n302) );
  inv02 U326 ( .Y(SUM[25]), .A(n303) );
  inv02 U327 ( .Y(carry_26_), .A(n304) );
  inv02 U328 ( .Y(n305), .A(B[25]) );
  inv02 U329 ( .Y(n306), .A(A[25]) );
  inv02 U330 ( .Y(n307), .A(n2) );
  nor02 U331 ( .Y(n308), .A0(n305), .A1(n309) );
  nor02 U332 ( .Y(n310), .A0(n306), .A1(n311) );
  nor02 U333 ( .Y(n312), .A0(n307), .A1(n313) );
  nor02 U334 ( .Y(n314), .A0(n307), .A1(n315) );
  nor02 U335 ( .Y(n303), .A0(n316), .A1(n317) );
  nor02 U336 ( .Y(n318), .A0(n306), .A1(n307) );
  nor02 U337 ( .Y(n319), .A0(n305), .A1(n307) );
  nor02 U338 ( .Y(n320), .A0(n305), .A1(n306) );
  nor02 U339 ( .Y(n304), .A0(n320), .A1(n321) );
  nor02 U340 ( .Y(n322), .A0(A[25]), .A1(n2) );
  inv01 U341 ( .Y(n309), .A(n322) );
  nor02 U342 ( .Y(n323), .A0(B[25]), .A1(n2) );
  inv01 U343 ( .Y(n311), .A(n323) );
  nor02 U344 ( .Y(n324), .A0(B[25]), .A1(A[25]) );
  inv01 U345 ( .Y(n313), .A(n324) );
  nor02 U346 ( .Y(n325), .A0(n305), .A1(n306) );
  inv01 U347 ( .Y(n315), .A(n325) );
  nor02 U348 ( .Y(n326), .A0(n308), .A1(n310) );
  inv01 U349 ( .Y(n316), .A(n326) );
  nor02 U350 ( .Y(n327), .A0(n312), .A1(n314) );
  inv01 U351 ( .Y(n317), .A(n327) );
  nor02 U352 ( .Y(n328), .A0(n318), .A1(n319) );
  inv01 U353 ( .Y(n321), .A(n328) );
  xor2 U354 ( .Y(SUM[47]), .A0(A[47]), .A1(carry_47_) );
  and02 U355 ( .Y(carry_47_), .A0(n18), .A1(A[46]) );
  xor2 U356 ( .Y(n329), .A0(A[46]), .A1(n18) );
  xor2 U357 ( .Y(n330), .A0(A[45]), .A1(n6) );
  xor2 U358 ( .Y(n331), .A0(A[44]), .A1(n16) );
  xor2 U359 ( .Y(n332), .A0(A[43]), .A1(n4) );
  xor2 U360 ( .Y(n333), .A0(A[42]), .A1(n14) );
  xor2 U361 ( .Y(n334), .A0(A[41]), .A1(n12) );
  xor2 U362 ( .Y(n335), .A0(A[40]), .A1(n10) );
  xor2 U363 ( .Y(n336), .A0(A[39]), .A1(n20) );
  xor2 U364 ( .Y(n337), .A0(A[38]), .A1(n22) );
  xor2 U365 ( .Y(n338), .A0(A[37]), .A1(n8) );
  xor2 U366 ( .Y(n339), .A0(A[36]), .A1(carry_36_) );
  xor2 U367 ( .Y(n340), .A0(B[24]), .A1(A[24]) );
endmodule


module mul_24_DW01_add_24_2 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   carry_23_, carry_22_, carry_21_, carry_20_, carry_19_, carry_18_,
         carry_17_, carry_16_, carry_15_, carry_14_, carry_13_, carry_12_,
         carry_11_, carry_10_, carry_9_, carry_8_, carry_7_, carry_6_,
         carry_5_, carry_4_, carry_3_, carry_2_, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549;

  nand02 U4 ( .Y(n1), .A0(A[0]), .A1(B[0]) );
  inv02 U5 ( .Y(n2), .A(n1) );
  buf02 U6 ( .Y(n3), .A(carry_23_) );
  inv01 U7 ( .Y(SUM[21]), .A(n4) );
  inv02 U8 ( .Y(carry_22_), .A(n5) );
  inv02 U9 ( .Y(n6), .A(B[21]) );
  inv02 U10 ( .Y(n7), .A(A[21]) );
  inv02 U11 ( .Y(n8), .A(carry_21_) );
  nor02 U12 ( .Y(n9), .A0(n6), .A1(n10) );
  nor02 U13 ( .Y(n11), .A0(n7), .A1(n12) );
  nor02 U14 ( .Y(n13), .A0(n8), .A1(n14) );
  nor02 U15 ( .Y(n15), .A0(n8), .A1(n16) );
  nor02 U16 ( .Y(n4), .A0(n17), .A1(n18) );
  nor02 U17 ( .Y(n19), .A0(n7), .A1(n8) );
  nor02 U18 ( .Y(n20), .A0(n6), .A1(n8) );
  nor02 U19 ( .Y(n21), .A0(n6), .A1(n7) );
  nor02 U20 ( .Y(n5), .A0(n21), .A1(n22) );
  nor02 U21 ( .Y(n23), .A0(A[21]), .A1(carry_21_) );
  inv01 U22 ( .Y(n10), .A(n23) );
  nor02 U23 ( .Y(n24), .A0(B[21]), .A1(carry_21_) );
  inv01 U24 ( .Y(n12), .A(n24) );
  nor02 U25 ( .Y(n25), .A0(B[21]), .A1(A[21]) );
  inv01 U26 ( .Y(n14), .A(n25) );
  nor02 U27 ( .Y(n26), .A0(n6), .A1(n7) );
  inv01 U28 ( .Y(n16), .A(n26) );
  nor02 U29 ( .Y(n27), .A0(n9), .A1(n11) );
  inv01 U30 ( .Y(n17), .A(n27) );
  nor02 U31 ( .Y(n28), .A0(n13), .A1(n15) );
  inv01 U32 ( .Y(n18), .A(n28) );
  nor02 U33 ( .Y(n29), .A0(n19), .A1(n20) );
  inv01 U34 ( .Y(n22), .A(n29) );
  inv01 U35 ( .Y(SUM[20]), .A(n30) );
  inv02 U36 ( .Y(carry_21_), .A(n31) );
  inv02 U37 ( .Y(n32), .A(B[20]) );
  inv02 U38 ( .Y(n33), .A(A[20]) );
  inv02 U39 ( .Y(n34), .A(carry_20_) );
  nor02 U40 ( .Y(n35), .A0(n32), .A1(n36) );
  nor02 U41 ( .Y(n37), .A0(n33), .A1(n38) );
  nor02 U42 ( .Y(n39), .A0(n34), .A1(n40) );
  nor02 U43 ( .Y(n41), .A0(n34), .A1(n42) );
  nor02 U44 ( .Y(n30), .A0(n43), .A1(n44) );
  nor02 U45 ( .Y(n45), .A0(n33), .A1(n34) );
  nor02 U46 ( .Y(n46), .A0(n32), .A1(n34) );
  nor02 U47 ( .Y(n47), .A0(n32), .A1(n33) );
  nor02 U48 ( .Y(n31), .A0(n47), .A1(n48) );
  nor02 U49 ( .Y(n49), .A0(A[20]), .A1(carry_20_) );
  inv01 U50 ( .Y(n36), .A(n49) );
  nor02 U51 ( .Y(n50), .A0(B[20]), .A1(carry_20_) );
  inv01 U52 ( .Y(n38), .A(n50) );
  nor02 U53 ( .Y(n51), .A0(B[20]), .A1(A[20]) );
  inv01 U54 ( .Y(n40), .A(n51) );
  nor02 U55 ( .Y(n52), .A0(n32), .A1(n33) );
  inv01 U56 ( .Y(n42), .A(n52) );
  nor02 U57 ( .Y(n53), .A0(n35), .A1(n37) );
  inv01 U58 ( .Y(n43), .A(n53) );
  nor02 U59 ( .Y(n54), .A0(n39), .A1(n41) );
  inv01 U60 ( .Y(n44), .A(n54) );
  nor02 U61 ( .Y(n55), .A0(n45), .A1(n46) );
  inv01 U62 ( .Y(n48), .A(n55) );
  inv01 U63 ( .Y(SUM[19]), .A(n56) );
  inv02 U64 ( .Y(carry_20_), .A(n57) );
  inv02 U65 ( .Y(n58), .A(B[19]) );
  inv02 U66 ( .Y(n59), .A(A[19]) );
  inv02 U67 ( .Y(n60), .A(carry_19_) );
  nor02 U68 ( .Y(n61), .A0(n58), .A1(n62) );
  nor02 U69 ( .Y(n63), .A0(n59), .A1(n64) );
  nor02 U70 ( .Y(n65), .A0(n60), .A1(n66) );
  nor02 U71 ( .Y(n67), .A0(n60), .A1(n68) );
  nor02 U72 ( .Y(n56), .A0(n69), .A1(n70) );
  nor02 U73 ( .Y(n71), .A0(n59), .A1(n60) );
  nor02 U74 ( .Y(n72), .A0(n58), .A1(n60) );
  nor02 U75 ( .Y(n73), .A0(n58), .A1(n59) );
  nor02 U76 ( .Y(n57), .A0(n73), .A1(n74) );
  nor02 U77 ( .Y(n75), .A0(A[19]), .A1(carry_19_) );
  inv01 U78 ( .Y(n62), .A(n75) );
  nor02 U79 ( .Y(n76), .A0(B[19]), .A1(carry_19_) );
  inv01 U80 ( .Y(n64), .A(n76) );
  nor02 U81 ( .Y(n77), .A0(B[19]), .A1(A[19]) );
  inv01 U82 ( .Y(n66), .A(n77) );
  nor02 U83 ( .Y(n78), .A0(n58), .A1(n59) );
  inv01 U84 ( .Y(n68), .A(n78) );
  nor02 U85 ( .Y(n79), .A0(n61), .A1(n63) );
  inv01 U86 ( .Y(n69), .A(n79) );
  nor02 U87 ( .Y(n80), .A0(n65), .A1(n67) );
  inv01 U88 ( .Y(n70), .A(n80) );
  nor02 U89 ( .Y(n81), .A0(n71), .A1(n72) );
  inv01 U90 ( .Y(n74), .A(n81) );
  inv01 U91 ( .Y(SUM[18]), .A(n82) );
  inv02 U92 ( .Y(carry_19_), .A(n83) );
  inv02 U93 ( .Y(n84), .A(B[18]) );
  inv02 U94 ( .Y(n85), .A(A[18]) );
  inv02 U95 ( .Y(n86), .A(carry_18_) );
  nor02 U96 ( .Y(n87), .A0(n84), .A1(n88) );
  nor02 U97 ( .Y(n89), .A0(n85), .A1(n90) );
  nor02 U98 ( .Y(n91), .A0(n86), .A1(n92) );
  nor02 U99 ( .Y(n93), .A0(n86), .A1(n94) );
  nor02 U100 ( .Y(n82), .A0(n95), .A1(n96) );
  nor02 U101 ( .Y(n97), .A0(n85), .A1(n86) );
  nor02 U102 ( .Y(n98), .A0(n84), .A1(n86) );
  nor02 U103 ( .Y(n99), .A0(n84), .A1(n85) );
  nor02 U104 ( .Y(n83), .A0(n99), .A1(n100) );
  nor02 U105 ( .Y(n101), .A0(A[18]), .A1(carry_18_) );
  inv01 U106 ( .Y(n88), .A(n101) );
  nor02 U107 ( .Y(n102), .A0(B[18]), .A1(carry_18_) );
  inv01 U108 ( .Y(n90), .A(n102) );
  nor02 U109 ( .Y(n103), .A0(B[18]), .A1(A[18]) );
  inv01 U110 ( .Y(n92), .A(n103) );
  nor02 U111 ( .Y(n104), .A0(n84), .A1(n85) );
  inv01 U112 ( .Y(n94), .A(n104) );
  nor02 U113 ( .Y(n105), .A0(n87), .A1(n89) );
  inv01 U114 ( .Y(n95), .A(n105) );
  nor02 U115 ( .Y(n106), .A0(n91), .A1(n93) );
  inv01 U116 ( .Y(n96), .A(n106) );
  nor02 U117 ( .Y(n107), .A0(n97), .A1(n98) );
  inv01 U118 ( .Y(n100), .A(n107) );
  inv01 U119 ( .Y(SUM[17]), .A(n108) );
  inv02 U120 ( .Y(carry_18_), .A(n109) );
  inv02 U121 ( .Y(n110), .A(B[17]) );
  inv02 U122 ( .Y(n111), .A(A[17]) );
  inv02 U123 ( .Y(n112), .A(carry_17_) );
  nor02 U124 ( .Y(n113), .A0(n110), .A1(n114) );
  nor02 U125 ( .Y(n115), .A0(n111), .A1(n116) );
  nor02 U126 ( .Y(n117), .A0(n112), .A1(n118) );
  nor02 U127 ( .Y(n119), .A0(n112), .A1(n120) );
  nor02 U128 ( .Y(n108), .A0(n121), .A1(n122) );
  nor02 U129 ( .Y(n123), .A0(n111), .A1(n112) );
  nor02 U130 ( .Y(n124), .A0(n110), .A1(n112) );
  nor02 U131 ( .Y(n125), .A0(n110), .A1(n111) );
  nor02 U132 ( .Y(n109), .A0(n125), .A1(n126) );
  nor02 U133 ( .Y(n127), .A0(A[17]), .A1(carry_17_) );
  inv01 U134 ( .Y(n114), .A(n127) );
  nor02 U135 ( .Y(n128), .A0(B[17]), .A1(carry_17_) );
  inv01 U136 ( .Y(n116), .A(n128) );
  nor02 U137 ( .Y(n129), .A0(B[17]), .A1(A[17]) );
  inv01 U138 ( .Y(n118), .A(n129) );
  nor02 U139 ( .Y(n130), .A0(n110), .A1(n111) );
  inv01 U140 ( .Y(n120), .A(n130) );
  nor02 U141 ( .Y(n131), .A0(n113), .A1(n115) );
  inv01 U142 ( .Y(n121), .A(n131) );
  nor02 U143 ( .Y(n132), .A0(n117), .A1(n119) );
  inv01 U144 ( .Y(n122), .A(n132) );
  nor02 U145 ( .Y(n133), .A0(n123), .A1(n124) );
  inv01 U146 ( .Y(n126), .A(n133) );
  inv01 U147 ( .Y(SUM[16]), .A(n134) );
  inv02 U148 ( .Y(carry_17_), .A(n135) );
  inv02 U149 ( .Y(n136), .A(B[16]) );
  inv02 U150 ( .Y(n137), .A(A[16]) );
  inv02 U151 ( .Y(n138), .A(carry_16_) );
  nor02 U152 ( .Y(n139), .A0(n136), .A1(n140) );
  nor02 U153 ( .Y(n141), .A0(n137), .A1(n142) );
  nor02 U154 ( .Y(n143), .A0(n138), .A1(n144) );
  nor02 U155 ( .Y(n145), .A0(n138), .A1(n146) );
  nor02 U156 ( .Y(n134), .A0(n147), .A1(n148) );
  nor02 U157 ( .Y(n149), .A0(n137), .A1(n138) );
  nor02 U158 ( .Y(n150), .A0(n136), .A1(n138) );
  nor02 U159 ( .Y(n151), .A0(n136), .A1(n137) );
  nor02 U160 ( .Y(n135), .A0(n151), .A1(n152) );
  nor02 U161 ( .Y(n153), .A0(A[16]), .A1(carry_16_) );
  inv01 U162 ( .Y(n140), .A(n153) );
  nor02 U163 ( .Y(n154), .A0(B[16]), .A1(carry_16_) );
  inv01 U164 ( .Y(n142), .A(n154) );
  nor02 U165 ( .Y(n155), .A0(B[16]), .A1(A[16]) );
  inv01 U166 ( .Y(n144), .A(n155) );
  nor02 U167 ( .Y(n156), .A0(n136), .A1(n137) );
  inv01 U168 ( .Y(n146), .A(n156) );
  nor02 U169 ( .Y(n157), .A0(n139), .A1(n141) );
  inv01 U170 ( .Y(n147), .A(n157) );
  nor02 U171 ( .Y(n158), .A0(n143), .A1(n145) );
  inv01 U172 ( .Y(n148), .A(n158) );
  nor02 U173 ( .Y(n159), .A0(n149), .A1(n150) );
  inv01 U174 ( .Y(n152), .A(n159) );
  inv01 U175 ( .Y(SUM[15]), .A(n160) );
  inv02 U176 ( .Y(carry_16_), .A(n161) );
  inv02 U177 ( .Y(n162), .A(B[15]) );
  inv02 U178 ( .Y(n163), .A(A[15]) );
  inv02 U179 ( .Y(n164), .A(carry_15_) );
  nor02 U180 ( .Y(n165), .A0(n162), .A1(n166) );
  nor02 U181 ( .Y(n167), .A0(n163), .A1(n168) );
  nor02 U182 ( .Y(n169), .A0(n164), .A1(n170) );
  nor02 U183 ( .Y(n171), .A0(n164), .A1(n172) );
  nor02 U184 ( .Y(n160), .A0(n173), .A1(n174) );
  nor02 U185 ( .Y(n175), .A0(n163), .A1(n164) );
  nor02 U186 ( .Y(n176), .A0(n162), .A1(n164) );
  nor02 U187 ( .Y(n177), .A0(n162), .A1(n163) );
  nor02 U188 ( .Y(n161), .A0(n177), .A1(n178) );
  nor02 U189 ( .Y(n179), .A0(A[15]), .A1(carry_15_) );
  inv01 U190 ( .Y(n166), .A(n179) );
  nor02 U191 ( .Y(n180), .A0(B[15]), .A1(carry_15_) );
  inv01 U192 ( .Y(n168), .A(n180) );
  nor02 U193 ( .Y(n181), .A0(B[15]), .A1(A[15]) );
  inv01 U194 ( .Y(n170), .A(n181) );
  nor02 U195 ( .Y(n182), .A0(n162), .A1(n163) );
  inv01 U196 ( .Y(n172), .A(n182) );
  nor02 U197 ( .Y(n183), .A0(n165), .A1(n167) );
  inv01 U198 ( .Y(n173), .A(n183) );
  nor02 U199 ( .Y(n184), .A0(n169), .A1(n171) );
  inv01 U200 ( .Y(n174), .A(n184) );
  nor02 U201 ( .Y(n185), .A0(n175), .A1(n176) );
  inv01 U202 ( .Y(n178), .A(n185) );
  inv01 U203 ( .Y(SUM[14]), .A(n186) );
  inv02 U204 ( .Y(carry_15_), .A(n187) );
  inv02 U205 ( .Y(n188), .A(B[14]) );
  inv02 U206 ( .Y(n189), .A(A[14]) );
  inv02 U207 ( .Y(n190), .A(carry_14_) );
  nor02 U208 ( .Y(n191), .A0(n188), .A1(n192) );
  nor02 U209 ( .Y(n193), .A0(n189), .A1(n194) );
  nor02 U210 ( .Y(n195), .A0(n190), .A1(n196) );
  nor02 U211 ( .Y(n197), .A0(n190), .A1(n198) );
  nor02 U212 ( .Y(n186), .A0(n199), .A1(n200) );
  nor02 U213 ( .Y(n201), .A0(n189), .A1(n190) );
  nor02 U214 ( .Y(n202), .A0(n188), .A1(n190) );
  nor02 U215 ( .Y(n203), .A0(n188), .A1(n189) );
  nor02 U216 ( .Y(n187), .A0(n203), .A1(n204) );
  nor02 U217 ( .Y(n205), .A0(A[14]), .A1(carry_14_) );
  inv01 U218 ( .Y(n192), .A(n205) );
  nor02 U219 ( .Y(n206), .A0(B[14]), .A1(carry_14_) );
  inv01 U220 ( .Y(n194), .A(n206) );
  nor02 U221 ( .Y(n207), .A0(B[14]), .A1(A[14]) );
  inv01 U222 ( .Y(n196), .A(n207) );
  nor02 U223 ( .Y(n208), .A0(n188), .A1(n189) );
  inv01 U224 ( .Y(n198), .A(n208) );
  nor02 U225 ( .Y(n209), .A0(n191), .A1(n193) );
  inv01 U226 ( .Y(n199), .A(n209) );
  nor02 U227 ( .Y(n210), .A0(n195), .A1(n197) );
  inv01 U228 ( .Y(n200), .A(n210) );
  nor02 U229 ( .Y(n211), .A0(n201), .A1(n202) );
  inv01 U230 ( .Y(n204), .A(n211) );
  inv01 U231 ( .Y(SUM[13]), .A(n212) );
  inv02 U232 ( .Y(carry_14_), .A(n213) );
  inv02 U233 ( .Y(n214), .A(B[13]) );
  inv02 U234 ( .Y(n215), .A(A[13]) );
  inv02 U235 ( .Y(n216), .A(carry_13_) );
  nor02 U236 ( .Y(n217), .A0(n214), .A1(n218) );
  nor02 U237 ( .Y(n219), .A0(n215), .A1(n220) );
  nor02 U238 ( .Y(n221), .A0(n216), .A1(n222) );
  nor02 U239 ( .Y(n223), .A0(n216), .A1(n224) );
  nor02 U240 ( .Y(n212), .A0(n225), .A1(n226) );
  nor02 U241 ( .Y(n227), .A0(n215), .A1(n216) );
  nor02 U242 ( .Y(n228), .A0(n214), .A1(n216) );
  nor02 U243 ( .Y(n229), .A0(n214), .A1(n215) );
  nor02 U244 ( .Y(n213), .A0(n229), .A1(n230) );
  nor02 U245 ( .Y(n231), .A0(A[13]), .A1(carry_13_) );
  inv01 U246 ( .Y(n218), .A(n231) );
  nor02 U247 ( .Y(n232), .A0(B[13]), .A1(carry_13_) );
  inv01 U248 ( .Y(n220), .A(n232) );
  nor02 U249 ( .Y(n233), .A0(B[13]), .A1(A[13]) );
  inv01 U250 ( .Y(n222), .A(n233) );
  nor02 U251 ( .Y(n234), .A0(n214), .A1(n215) );
  inv01 U252 ( .Y(n224), .A(n234) );
  nor02 U253 ( .Y(n235), .A0(n217), .A1(n219) );
  inv01 U254 ( .Y(n225), .A(n235) );
  nor02 U255 ( .Y(n236), .A0(n221), .A1(n223) );
  inv01 U256 ( .Y(n226), .A(n236) );
  nor02 U257 ( .Y(n237), .A0(n227), .A1(n228) );
  inv01 U258 ( .Y(n230), .A(n237) );
  inv01 U259 ( .Y(SUM[12]), .A(n238) );
  inv02 U260 ( .Y(carry_13_), .A(n239) );
  inv02 U261 ( .Y(n240), .A(B[12]) );
  inv02 U262 ( .Y(n241), .A(A[12]) );
  inv02 U263 ( .Y(n242), .A(carry_12_) );
  nor02 U264 ( .Y(n243), .A0(n240), .A1(n244) );
  nor02 U265 ( .Y(n245), .A0(n241), .A1(n246) );
  nor02 U266 ( .Y(n247), .A0(n242), .A1(n248) );
  nor02 U267 ( .Y(n249), .A0(n242), .A1(n250) );
  nor02 U268 ( .Y(n238), .A0(n251), .A1(n252) );
  nor02 U269 ( .Y(n253), .A0(n241), .A1(n242) );
  nor02 U270 ( .Y(n254), .A0(n240), .A1(n242) );
  nor02 U271 ( .Y(n255), .A0(n240), .A1(n241) );
  nor02 U272 ( .Y(n239), .A0(n255), .A1(n256) );
  nor02 U273 ( .Y(n257), .A0(A[12]), .A1(carry_12_) );
  inv01 U274 ( .Y(n244), .A(n257) );
  nor02 U275 ( .Y(n258), .A0(B[12]), .A1(carry_12_) );
  inv01 U276 ( .Y(n246), .A(n258) );
  nor02 U277 ( .Y(n259), .A0(B[12]), .A1(A[12]) );
  inv01 U278 ( .Y(n248), .A(n259) );
  nor02 U279 ( .Y(n260), .A0(n240), .A1(n241) );
  inv01 U280 ( .Y(n250), .A(n260) );
  nor02 U281 ( .Y(n261), .A0(n243), .A1(n245) );
  inv01 U282 ( .Y(n251), .A(n261) );
  nor02 U283 ( .Y(n262), .A0(n247), .A1(n249) );
  inv01 U284 ( .Y(n252), .A(n262) );
  nor02 U285 ( .Y(n263), .A0(n253), .A1(n254) );
  inv01 U286 ( .Y(n256), .A(n263) );
  inv01 U287 ( .Y(SUM[11]), .A(n264) );
  inv02 U288 ( .Y(carry_12_), .A(n265) );
  inv02 U289 ( .Y(n266), .A(B[11]) );
  inv02 U290 ( .Y(n267), .A(A[11]) );
  inv02 U291 ( .Y(n268), .A(carry_11_) );
  nor02 U292 ( .Y(n269), .A0(n266), .A1(n270) );
  nor02 U293 ( .Y(n271), .A0(n267), .A1(n272) );
  nor02 U294 ( .Y(n273), .A0(n268), .A1(n274) );
  nor02 U295 ( .Y(n275), .A0(n268), .A1(n276) );
  nor02 U296 ( .Y(n264), .A0(n277), .A1(n278) );
  nor02 U297 ( .Y(n279), .A0(n267), .A1(n268) );
  nor02 U298 ( .Y(n280), .A0(n266), .A1(n268) );
  nor02 U299 ( .Y(n281), .A0(n266), .A1(n267) );
  nor02 U300 ( .Y(n265), .A0(n281), .A1(n282) );
  nor02 U301 ( .Y(n283), .A0(A[11]), .A1(carry_11_) );
  inv01 U302 ( .Y(n270), .A(n283) );
  nor02 U303 ( .Y(n284), .A0(B[11]), .A1(carry_11_) );
  inv01 U304 ( .Y(n272), .A(n284) );
  nor02 U305 ( .Y(n285), .A0(B[11]), .A1(A[11]) );
  inv01 U306 ( .Y(n274), .A(n285) );
  nor02 U307 ( .Y(n286), .A0(n266), .A1(n267) );
  inv01 U308 ( .Y(n276), .A(n286) );
  nor02 U309 ( .Y(n287), .A0(n269), .A1(n271) );
  inv01 U310 ( .Y(n277), .A(n287) );
  nor02 U311 ( .Y(n288), .A0(n273), .A1(n275) );
  inv01 U312 ( .Y(n278), .A(n288) );
  nor02 U313 ( .Y(n289), .A0(n279), .A1(n280) );
  inv01 U314 ( .Y(n282), .A(n289) );
  inv01 U315 ( .Y(SUM[10]), .A(n290) );
  inv02 U316 ( .Y(carry_11_), .A(n291) );
  inv02 U317 ( .Y(n292), .A(B[10]) );
  inv02 U318 ( .Y(n293), .A(A[10]) );
  inv02 U319 ( .Y(n294), .A(carry_10_) );
  nor02 U320 ( .Y(n295), .A0(n292), .A1(n296) );
  nor02 U321 ( .Y(n297), .A0(n293), .A1(n298) );
  nor02 U322 ( .Y(n299), .A0(n294), .A1(n300) );
  nor02 U323 ( .Y(n301), .A0(n294), .A1(n302) );
  nor02 U324 ( .Y(n290), .A0(n303), .A1(n304) );
  nor02 U325 ( .Y(n305), .A0(n293), .A1(n294) );
  nor02 U326 ( .Y(n306), .A0(n292), .A1(n294) );
  nor02 U327 ( .Y(n307), .A0(n292), .A1(n293) );
  nor02 U328 ( .Y(n291), .A0(n307), .A1(n308) );
  nor02 U329 ( .Y(n309), .A0(A[10]), .A1(carry_10_) );
  inv01 U330 ( .Y(n296), .A(n309) );
  nor02 U331 ( .Y(n310), .A0(B[10]), .A1(carry_10_) );
  inv01 U332 ( .Y(n298), .A(n310) );
  nor02 U333 ( .Y(n311), .A0(B[10]), .A1(A[10]) );
  inv01 U334 ( .Y(n300), .A(n311) );
  nor02 U335 ( .Y(n312), .A0(n292), .A1(n293) );
  inv01 U336 ( .Y(n302), .A(n312) );
  nor02 U337 ( .Y(n313), .A0(n295), .A1(n297) );
  inv01 U338 ( .Y(n303), .A(n313) );
  nor02 U339 ( .Y(n314), .A0(n299), .A1(n301) );
  inv01 U340 ( .Y(n304), .A(n314) );
  nor02 U341 ( .Y(n315), .A0(n305), .A1(n306) );
  inv01 U342 ( .Y(n308), .A(n315) );
  inv01 U343 ( .Y(SUM[9]), .A(n316) );
  inv02 U344 ( .Y(carry_10_), .A(n317) );
  inv02 U345 ( .Y(n318), .A(B[9]) );
  inv02 U346 ( .Y(n319), .A(A[9]) );
  inv02 U347 ( .Y(n320), .A(carry_9_) );
  nor02 U348 ( .Y(n321), .A0(n318), .A1(n322) );
  nor02 U349 ( .Y(n323), .A0(n319), .A1(n324) );
  nor02 U350 ( .Y(n325), .A0(n320), .A1(n326) );
  nor02 U351 ( .Y(n327), .A0(n320), .A1(n328) );
  nor02 U352 ( .Y(n316), .A0(n329), .A1(n330) );
  nor02 U353 ( .Y(n331), .A0(n319), .A1(n320) );
  nor02 U354 ( .Y(n332), .A0(n318), .A1(n320) );
  nor02 U355 ( .Y(n333), .A0(n318), .A1(n319) );
  nor02 U356 ( .Y(n317), .A0(n333), .A1(n334) );
  nor02 U357 ( .Y(n335), .A0(A[9]), .A1(carry_9_) );
  inv01 U358 ( .Y(n322), .A(n335) );
  nor02 U359 ( .Y(n336), .A0(B[9]), .A1(carry_9_) );
  inv01 U360 ( .Y(n324), .A(n336) );
  nor02 U361 ( .Y(n337), .A0(B[9]), .A1(A[9]) );
  inv01 U362 ( .Y(n326), .A(n337) );
  nor02 U363 ( .Y(n338), .A0(n318), .A1(n319) );
  inv01 U364 ( .Y(n328), .A(n338) );
  nor02 U365 ( .Y(n339), .A0(n321), .A1(n323) );
  inv01 U366 ( .Y(n329), .A(n339) );
  nor02 U367 ( .Y(n340), .A0(n325), .A1(n327) );
  inv01 U368 ( .Y(n330), .A(n340) );
  nor02 U369 ( .Y(n341), .A0(n331), .A1(n332) );
  inv01 U370 ( .Y(n334), .A(n341) );
  inv01 U371 ( .Y(SUM[8]), .A(n342) );
  inv02 U372 ( .Y(carry_9_), .A(n343) );
  inv02 U373 ( .Y(n344), .A(B[8]) );
  inv02 U374 ( .Y(n345), .A(A[8]) );
  inv02 U375 ( .Y(n346), .A(carry_8_) );
  nor02 U376 ( .Y(n347), .A0(n344), .A1(n348) );
  nor02 U377 ( .Y(n349), .A0(n345), .A1(n350) );
  nor02 U378 ( .Y(n351), .A0(n346), .A1(n352) );
  nor02 U379 ( .Y(n353), .A0(n346), .A1(n354) );
  nor02 U380 ( .Y(n342), .A0(n355), .A1(n356) );
  nor02 U381 ( .Y(n357), .A0(n345), .A1(n346) );
  nor02 U382 ( .Y(n358), .A0(n344), .A1(n346) );
  nor02 U383 ( .Y(n359), .A0(n344), .A1(n345) );
  nor02 U384 ( .Y(n343), .A0(n359), .A1(n360) );
  nor02 U385 ( .Y(n361), .A0(A[8]), .A1(carry_8_) );
  inv01 U386 ( .Y(n348), .A(n361) );
  nor02 U387 ( .Y(n362), .A0(B[8]), .A1(carry_8_) );
  inv01 U388 ( .Y(n350), .A(n362) );
  nor02 U389 ( .Y(n363), .A0(B[8]), .A1(A[8]) );
  inv01 U390 ( .Y(n352), .A(n363) );
  nor02 U391 ( .Y(n364), .A0(n344), .A1(n345) );
  inv01 U392 ( .Y(n354), .A(n364) );
  nor02 U393 ( .Y(n365), .A0(n347), .A1(n349) );
  inv01 U394 ( .Y(n355), .A(n365) );
  nor02 U395 ( .Y(n366), .A0(n351), .A1(n353) );
  inv01 U396 ( .Y(n356), .A(n366) );
  nor02 U397 ( .Y(n367), .A0(n357), .A1(n358) );
  inv01 U398 ( .Y(n360), .A(n367) );
  inv01 U399 ( .Y(SUM[7]), .A(n368) );
  inv02 U400 ( .Y(carry_8_), .A(n369) );
  inv02 U401 ( .Y(n370), .A(B[7]) );
  inv02 U402 ( .Y(n371), .A(A[7]) );
  inv02 U403 ( .Y(n372), .A(carry_7_) );
  nor02 U404 ( .Y(n373), .A0(n370), .A1(n374) );
  nor02 U405 ( .Y(n375), .A0(n371), .A1(n376) );
  nor02 U406 ( .Y(n377), .A0(n372), .A1(n378) );
  nor02 U407 ( .Y(n379), .A0(n372), .A1(n380) );
  nor02 U408 ( .Y(n368), .A0(n381), .A1(n382) );
  nor02 U409 ( .Y(n383), .A0(n371), .A1(n372) );
  nor02 U410 ( .Y(n384), .A0(n370), .A1(n372) );
  nor02 U411 ( .Y(n385), .A0(n370), .A1(n371) );
  nor02 U412 ( .Y(n369), .A0(n385), .A1(n386) );
  nor02 U413 ( .Y(n387), .A0(A[7]), .A1(carry_7_) );
  inv01 U414 ( .Y(n374), .A(n387) );
  nor02 U415 ( .Y(n388), .A0(B[7]), .A1(carry_7_) );
  inv01 U416 ( .Y(n376), .A(n388) );
  nor02 U417 ( .Y(n389), .A0(B[7]), .A1(A[7]) );
  inv01 U418 ( .Y(n378), .A(n389) );
  nor02 U419 ( .Y(n390), .A0(n370), .A1(n371) );
  inv01 U420 ( .Y(n380), .A(n390) );
  nor02 U421 ( .Y(n391), .A0(n373), .A1(n375) );
  inv01 U422 ( .Y(n381), .A(n391) );
  nor02 U423 ( .Y(n392), .A0(n377), .A1(n379) );
  inv01 U424 ( .Y(n382), .A(n392) );
  nor02 U425 ( .Y(n393), .A0(n383), .A1(n384) );
  inv01 U426 ( .Y(n386), .A(n393) );
  inv01 U427 ( .Y(SUM[6]), .A(n394) );
  inv02 U428 ( .Y(carry_7_), .A(n395) );
  inv02 U429 ( .Y(n396), .A(B[6]) );
  inv02 U430 ( .Y(n397), .A(A[6]) );
  inv02 U431 ( .Y(n398), .A(carry_6_) );
  nor02 U432 ( .Y(n399), .A0(n396), .A1(n400) );
  nor02 U433 ( .Y(n401), .A0(n397), .A1(n402) );
  nor02 U434 ( .Y(n403), .A0(n398), .A1(n404) );
  nor02 U435 ( .Y(n405), .A0(n398), .A1(n406) );
  nor02 U436 ( .Y(n394), .A0(n407), .A1(n408) );
  nor02 U437 ( .Y(n409), .A0(n397), .A1(n398) );
  nor02 U438 ( .Y(n410), .A0(n396), .A1(n398) );
  nor02 U439 ( .Y(n411), .A0(n396), .A1(n397) );
  nor02 U440 ( .Y(n395), .A0(n411), .A1(n412) );
  nor02 U441 ( .Y(n413), .A0(A[6]), .A1(carry_6_) );
  inv01 U442 ( .Y(n400), .A(n413) );
  nor02 U443 ( .Y(n414), .A0(B[6]), .A1(carry_6_) );
  inv01 U444 ( .Y(n402), .A(n414) );
  nor02 U445 ( .Y(n415), .A0(B[6]), .A1(A[6]) );
  inv01 U446 ( .Y(n404), .A(n415) );
  nor02 U447 ( .Y(n416), .A0(n396), .A1(n397) );
  inv01 U448 ( .Y(n406), .A(n416) );
  nor02 U449 ( .Y(n417), .A0(n399), .A1(n401) );
  inv01 U450 ( .Y(n407), .A(n417) );
  nor02 U451 ( .Y(n418), .A0(n403), .A1(n405) );
  inv01 U452 ( .Y(n408), .A(n418) );
  nor02 U453 ( .Y(n419), .A0(n409), .A1(n410) );
  inv01 U454 ( .Y(n412), .A(n419) );
  inv01 U455 ( .Y(SUM[5]), .A(n420) );
  inv02 U456 ( .Y(carry_6_), .A(n421) );
  inv02 U457 ( .Y(n422), .A(B[5]) );
  inv02 U458 ( .Y(n423), .A(A[5]) );
  inv02 U459 ( .Y(n424), .A(carry_5_) );
  nor02 U460 ( .Y(n425), .A0(n422), .A1(n426) );
  nor02 U461 ( .Y(n427), .A0(n423), .A1(n428) );
  nor02 U462 ( .Y(n429), .A0(n424), .A1(n430) );
  nor02 U463 ( .Y(n431), .A0(n424), .A1(n432) );
  nor02 U464 ( .Y(n420), .A0(n433), .A1(n434) );
  nor02 U465 ( .Y(n435), .A0(n423), .A1(n424) );
  nor02 U466 ( .Y(n436), .A0(n422), .A1(n424) );
  nor02 U467 ( .Y(n437), .A0(n422), .A1(n423) );
  nor02 U468 ( .Y(n421), .A0(n437), .A1(n438) );
  nor02 U469 ( .Y(n439), .A0(A[5]), .A1(carry_5_) );
  inv01 U470 ( .Y(n426), .A(n439) );
  nor02 U471 ( .Y(n440), .A0(B[5]), .A1(carry_5_) );
  inv01 U472 ( .Y(n428), .A(n440) );
  nor02 U473 ( .Y(n441), .A0(B[5]), .A1(A[5]) );
  inv01 U474 ( .Y(n430), .A(n441) );
  nor02 U475 ( .Y(n442), .A0(n422), .A1(n423) );
  inv01 U476 ( .Y(n432), .A(n442) );
  nor02 U477 ( .Y(n443), .A0(n425), .A1(n427) );
  inv01 U478 ( .Y(n433), .A(n443) );
  nor02 U479 ( .Y(n444), .A0(n429), .A1(n431) );
  inv01 U480 ( .Y(n434), .A(n444) );
  nor02 U481 ( .Y(n445), .A0(n435), .A1(n436) );
  inv01 U482 ( .Y(n438), .A(n445) );
  inv01 U483 ( .Y(SUM[4]), .A(n446) );
  inv02 U484 ( .Y(carry_5_), .A(n447) );
  inv02 U485 ( .Y(n448), .A(B[4]) );
  inv02 U486 ( .Y(n449), .A(A[4]) );
  inv02 U487 ( .Y(n450), .A(carry_4_) );
  nor02 U488 ( .Y(n451), .A0(n448), .A1(n452) );
  nor02 U489 ( .Y(n453), .A0(n449), .A1(n454) );
  nor02 U490 ( .Y(n455), .A0(n450), .A1(n456) );
  nor02 U491 ( .Y(n457), .A0(n450), .A1(n458) );
  nor02 U492 ( .Y(n446), .A0(n459), .A1(n460) );
  nor02 U493 ( .Y(n461), .A0(n449), .A1(n450) );
  nor02 U494 ( .Y(n462), .A0(n448), .A1(n450) );
  nor02 U495 ( .Y(n463), .A0(n448), .A1(n449) );
  nor02 U496 ( .Y(n447), .A0(n463), .A1(n464) );
  nor02 U497 ( .Y(n465), .A0(A[4]), .A1(carry_4_) );
  inv01 U498 ( .Y(n452), .A(n465) );
  nor02 U499 ( .Y(n466), .A0(B[4]), .A1(carry_4_) );
  inv01 U500 ( .Y(n454), .A(n466) );
  nor02 U501 ( .Y(n467), .A0(B[4]), .A1(A[4]) );
  inv01 U502 ( .Y(n456), .A(n467) );
  nor02 U503 ( .Y(n468), .A0(n448), .A1(n449) );
  inv01 U504 ( .Y(n458), .A(n468) );
  nor02 U505 ( .Y(n469), .A0(n451), .A1(n453) );
  inv01 U506 ( .Y(n459), .A(n469) );
  nor02 U507 ( .Y(n470), .A0(n455), .A1(n457) );
  inv01 U508 ( .Y(n460), .A(n470) );
  nor02 U509 ( .Y(n471), .A0(n461), .A1(n462) );
  inv01 U510 ( .Y(n464), .A(n471) );
  inv01 U511 ( .Y(SUM[3]), .A(n472) );
  inv02 U512 ( .Y(carry_4_), .A(n473) );
  inv02 U513 ( .Y(n474), .A(B[3]) );
  inv02 U514 ( .Y(n475), .A(A[3]) );
  inv02 U515 ( .Y(n476), .A(carry_3_) );
  nor02 U516 ( .Y(n477), .A0(n474), .A1(n478) );
  nor02 U517 ( .Y(n479), .A0(n475), .A1(n480) );
  nor02 U518 ( .Y(n481), .A0(n476), .A1(n482) );
  nor02 U519 ( .Y(n483), .A0(n476), .A1(n484) );
  nor02 U520 ( .Y(n472), .A0(n485), .A1(n486) );
  nor02 U521 ( .Y(n487), .A0(n475), .A1(n476) );
  nor02 U522 ( .Y(n488), .A0(n474), .A1(n476) );
  nor02 U523 ( .Y(n489), .A0(n474), .A1(n475) );
  nor02 U524 ( .Y(n473), .A0(n489), .A1(n490) );
  nor02 U525 ( .Y(n491), .A0(A[3]), .A1(carry_3_) );
  inv01 U526 ( .Y(n478), .A(n491) );
  nor02 U527 ( .Y(n492), .A0(B[3]), .A1(carry_3_) );
  inv01 U528 ( .Y(n480), .A(n492) );
  nor02 U529 ( .Y(n493), .A0(B[3]), .A1(A[3]) );
  inv01 U530 ( .Y(n482), .A(n493) );
  nor02 U531 ( .Y(n494), .A0(n474), .A1(n475) );
  inv01 U532 ( .Y(n484), .A(n494) );
  nor02 U533 ( .Y(n495), .A0(n477), .A1(n479) );
  inv01 U534 ( .Y(n485), .A(n495) );
  nor02 U535 ( .Y(n496), .A0(n481), .A1(n483) );
  inv01 U536 ( .Y(n486), .A(n496) );
  nor02 U537 ( .Y(n497), .A0(n487), .A1(n488) );
  inv01 U538 ( .Y(n490), .A(n497) );
  inv01 U539 ( .Y(SUM[2]), .A(n498) );
  inv02 U540 ( .Y(carry_3_), .A(n499) );
  inv02 U541 ( .Y(n500), .A(B[2]) );
  inv02 U542 ( .Y(n501), .A(A[2]) );
  inv02 U543 ( .Y(n502), .A(carry_2_) );
  nor02 U544 ( .Y(n503), .A0(n500), .A1(n504) );
  nor02 U545 ( .Y(n505), .A0(n501), .A1(n506) );
  nor02 U546 ( .Y(n507), .A0(n502), .A1(n508) );
  nor02 U547 ( .Y(n509), .A0(n502), .A1(n510) );
  nor02 U548 ( .Y(n498), .A0(n511), .A1(n512) );
  nor02 U549 ( .Y(n513), .A0(n501), .A1(n502) );
  nor02 U550 ( .Y(n514), .A0(n500), .A1(n502) );
  nor02 U551 ( .Y(n515), .A0(n500), .A1(n501) );
  nor02 U552 ( .Y(n499), .A0(n515), .A1(n516) );
  nor02 U553 ( .Y(n517), .A0(A[2]), .A1(carry_2_) );
  inv01 U554 ( .Y(n504), .A(n517) );
  nor02 U555 ( .Y(n518), .A0(B[2]), .A1(carry_2_) );
  inv01 U556 ( .Y(n506), .A(n518) );
  nor02 U557 ( .Y(n519), .A0(B[2]), .A1(A[2]) );
  inv01 U558 ( .Y(n508), .A(n519) );
  nor02 U559 ( .Y(n520), .A0(n500), .A1(n501) );
  inv01 U560 ( .Y(n510), .A(n520) );
  nor02 U561 ( .Y(n521), .A0(n503), .A1(n505) );
  inv01 U562 ( .Y(n511), .A(n521) );
  nor02 U563 ( .Y(n522), .A0(n507), .A1(n509) );
  inv01 U564 ( .Y(n512), .A(n522) );
  nor02 U565 ( .Y(n523), .A0(n513), .A1(n514) );
  inv01 U566 ( .Y(n516), .A(n523) );
  inv01 U567 ( .Y(SUM[1]), .A(n524) );
  inv02 U568 ( .Y(carry_2_), .A(n525) );
  inv02 U569 ( .Y(n526), .A(B[1]) );
  inv02 U570 ( .Y(n527), .A(A[1]) );
  inv02 U571 ( .Y(n528), .A(n2) );
  nor02 U572 ( .Y(n529), .A0(n526), .A1(n530) );
  nor02 U573 ( .Y(n531), .A0(n527), .A1(n532) );
  nor02 U574 ( .Y(n533), .A0(n528), .A1(n534) );
  nor02 U575 ( .Y(n535), .A0(n528), .A1(n536) );
  nor02 U576 ( .Y(n524), .A0(n537), .A1(n538) );
  nor02 U577 ( .Y(n539), .A0(n527), .A1(n528) );
  nor02 U578 ( .Y(n540), .A0(n526), .A1(n528) );
  nor02 U579 ( .Y(n541), .A0(n526), .A1(n527) );
  nor02 U580 ( .Y(n525), .A0(n541), .A1(n542) );
  nor02 U581 ( .Y(n543), .A0(A[1]), .A1(n2) );
  inv01 U582 ( .Y(n530), .A(n543) );
  nor02 U583 ( .Y(n544), .A0(B[1]), .A1(n2) );
  inv01 U584 ( .Y(n532), .A(n544) );
  nor02 U585 ( .Y(n545), .A0(B[1]), .A1(A[1]) );
  inv01 U586 ( .Y(n534), .A(n545) );
  nor02 U587 ( .Y(n546), .A0(n526), .A1(n527) );
  inv01 U588 ( .Y(n536), .A(n546) );
  nor02 U589 ( .Y(n547), .A0(n529), .A1(n531) );
  inv01 U590 ( .Y(n537), .A(n547) );
  nor02 U591 ( .Y(n548), .A0(n533), .A1(n535) );
  inv01 U592 ( .Y(n538), .A(n548) );
  nor02 U593 ( .Y(n549), .A0(n539), .A1(n540) );
  inv01 U594 ( .Y(n542), .A(n549) );
  xor2 U595 ( .Y(SUM[0]), .A0(B[0]), .A1(A[0]) );
  fadd1 U1_22 ( .S(SUM[22]), .CO(carry_23_), .A(A[22]), .B(B[22]), .CI(
        carry_22_) );
  fadd1 U1_23 ( .S(SUM[23]), .A(A[23]), .B(B[23]), .CI(n3) );
endmodule


module mul_24_DW01_add_24_1 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   carry_23_, carry_22_, carry_21_, carry_20_, carry_19_, carry_18_,
         carry_17_, carry_16_, carry_15_, carry_14_, carry_13_, carry_12_,
         carry_11_, carry_10_, carry_9_, carry_8_, carry_7_, carry_6_,
         carry_5_, carry_4_, carry_3_, carry_2_, n577, n578, n2, n3, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576;

  buf02 U4 ( .Y(SUM[0]), .A(n578) );
  nand02 U5 ( .Y(n2), .A0(A[0]), .A1(B[0]) );
  inv02 U6 ( .Y(n3), .A(n2) );
  buf02 U7 ( .Y(SUM[23]), .A(n577) );
  inv02 U8 ( .Y(SUM[21]), .A(n5) );
  inv02 U9 ( .Y(carry_22_), .A(n6) );
  inv02 U10 ( .Y(n7), .A(B[21]) );
  inv02 U11 ( .Y(n8), .A(A[21]) );
  inv02 U12 ( .Y(n9), .A(carry_21_) );
  nor02 U13 ( .Y(n10), .A0(n7), .A1(n11) );
  nor02 U14 ( .Y(n12), .A0(n8), .A1(n13) );
  nor02 U15 ( .Y(n14), .A0(n9), .A1(n15) );
  nor02 U16 ( .Y(n16), .A0(n9), .A1(n17) );
  nor02 U17 ( .Y(n5), .A0(n18), .A1(n19) );
  nor02 U18 ( .Y(n20), .A0(n8), .A1(n9) );
  nor02 U19 ( .Y(n21), .A0(n7), .A1(n9) );
  nor02 U20 ( .Y(n22), .A0(n7), .A1(n8) );
  nor02 U21 ( .Y(n6), .A0(n22), .A1(n23) );
  nor02 U22 ( .Y(n24), .A0(A[21]), .A1(carry_21_) );
  inv01 U23 ( .Y(n11), .A(n24) );
  nor02 U24 ( .Y(n25), .A0(B[21]), .A1(carry_21_) );
  inv01 U25 ( .Y(n13), .A(n25) );
  nor02 U26 ( .Y(n26), .A0(B[21]), .A1(A[21]) );
  inv01 U27 ( .Y(n15), .A(n26) );
  nor02 U28 ( .Y(n27), .A0(n7), .A1(n8) );
  inv01 U29 ( .Y(n17), .A(n27) );
  nor02 U30 ( .Y(n28), .A0(n10), .A1(n12) );
  inv01 U31 ( .Y(n18), .A(n28) );
  nor02 U32 ( .Y(n29), .A0(n14), .A1(n16) );
  inv01 U33 ( .Y(n19), .A(n29) );
  nor02 U34 ( .Y(n30), .A0(n20), .A1(n21) );
  inv01 U35 ( .Y(n23), .A(n30) );
  inv02 U36 ( .Y(SUM[22]), .A(n31) );
  inv02 U37 ( .Y(carry_23_), .A(n32) );
  inv02 U38 ( .Y(n33), .A(B[22]) );
  inv02 U39 ( .Y(n34), .A(A[22]) );
  inv02 U40 ( .Y(n35), .A(carry_22_) );
  nor02 U41 ( .Y(n36), .A0(n33), .A1(n37) );
  nor02 U42 ( .Y(n38), .A0(n34), .A1(n39) );
  nor02 U43 ( .Y(n40), .A0(n35), .A1(n41) );
  nor02 U44 ( .Y(n42), .A0(n35), .A1(n43) );
  nor02 U45 ( .Y(n31), .A0(n44), .A1(n45) );
  nor02 U46 ( .Y(n46), .A0(n34), .A1(n35) );
  nor02 U47 ( .Y(n47), .A0(n33), .A1(n35) );
  nor02 U48 ( .Y(n48), .A0(n33), .A1(n34) );
  nor02 U49 ( .Y(n32), .A0(n48), .A1(n49) );
  nor02 U50 ( .Y(n50), .A0(A[22]), .A1(carry_22_) );
  inv01 U51 ( .Y(n37), .A(n50) );
  nor02 U52 ( .Y(n51), .A0(B[22]), .A1(carry_22_) );
  inv01 U53 ( .Y(n39), .A(n51) );
  nor02 U54 ( .Y(n52), .A0(B[22]), .A1(A[22]) );
  inv01 U55 ( .Y(n41), .A(n52) );
  nor02 U56 ( .Y(n53), .A0(n33), .A1(n34) );
  inv01 U57 ( .Y(n43), .A(n53) );
  nor02 U58 ( .Y(n54), .A0(n36), .A1(n38) );
  inv01 U59 ( .Y(n44), .A(n54) );
  nor02 U60 ( .Y(n55), .A0(n40), .A1(n42) );
  inv01 U61 ( .Y(n45), .A(n55) );
  nor02 U62 ( .Y(n56), .A0(n46), .A1(n47) );
  inv01 U63 ( .Y(n49), .A(n56) );
  inv02 U64 ( .Y(SUM[19]), .A(n57) );
  inv02 U65 ( .Y(carry_20_), .A(n58) );
  inv02 U66 ( .Y(n59), .A(B[19]) );
  inv02 U67 ( .Y(n60), .A(A[19]) );
  inv02 U68 ( .Y(n61), .A(carry_19_) );
  nor02 U69 ( .Y(n62), .A0(n59), .A1(n63) );
  nor02 U70 ( .Y(n64), .A0(n60), .A1(n65) );
  nor02 U71 ( .Y(n66), .A0(n61), .A1(n67) );
  nor02 U72 ( .Y(n68), .A0(n61), .A1(n69) );
  nor02 U73 ( .Y(n57), .A0(n70), .A1(n71) );
  nor02 U74 ( .Y(n72), .A0(n60), .A1(n61) );
  nor02 U75 ( .Y(n73), .A0(n59), .A1(n61) );
  nor02 U76 ( .Y(n74), .A0(n59), .A1(n60) );
  nor02 U77 ( .Y(n58), .A0(n74), .A1(n75) );
  nor02 U78 ( .Y(n76), .A0(A[19]), .A1(carry_19_) );
  inv01 U79 ( .Y(n63), .A(n76) );
  nor02 U80 ( .Y(n77), .A0(B[19]), .A1(carry_19_) );
  inv01 U81 ( .Y(n65), .A(n77) );
  nor02 U82 ( .Y(n78), .A0(B[19]), .A1(A[19]) );
  inv01 U83 ( .Y(n67), .A(n78) );
  nor02 U84 ( .Y(n79), .A0(n59), .A1(n60) );
  inv01 U85 ( .Y(n69), .A(n79) );
  nor02 U86 ( .Y(n80), .A0(n62), .A1(n64) );
  inv01 U87 ( .Y(n70), .A(n80) );
  nor02 U88 ( .Y(n81), .A0(n66), .A1(n68) );
  inv01 U89 ( .Y(n71), .A(n81) );
  nor02 U90 ( .Y(n82), .A0(n72), .A1(n73) );
  inv01 U91 ( .Y(n75), .A(n82) );
  inv02 U92 ( .Y(SUM[20]), .A(n83) );
  inv02 U93 ( .Y(carry_21_), .A(n84) );
  inv02 U94 ( .Y(n85), .A(B[20]) );
  inv02 U95 ( .Y(n86), .A(A[20]) );
  inv02 U96 ( .Y(n87), .A(carry_20_) );
  nor02 U97 ( .Y(n88), .A0(n85), .A1(n89) );
  nor02 U98 ( .Y(n90), .A0(n86), .A1(n91) );
  nor02 U99 ( .Y(n92), .A0(n87), .A1(n93) );
  nor02 U100 ( .Y(n94), .A0(n87), .A1(n95) );
  nor02 U101 ( .Y(n83), .A0(n96), .A1(n97) );
  nor02 U102 ( .Y(n98), .A0(n86), .A1(n87) );
  nor02 U103 ( .Y(n99), .A0(n85), .A1(n87) );
  nor02 U104 ( .Y(n100), .A0(n85), .A1(n86) );
  nor02 U105 ( .Y(n84), .A0(n100), .A1(n101) );
  nor02 U106 ( .Y(n102), .A0(A[20]), .A1(carry_20_) );
  inv01 U107 ( .Y(n89), .A(n102) );
  nor02 U108 ( .Y(n103), .A0(B[20]), .A1(carry_20_) );
  inv01 U109 ( .Y(n91), .A(n103) );
  nor02 U110 ( .Y(n104), .A0(B[20]), .A1(A[20]) );
  inv01 U111 ( .Y(n93), .A(n104) );
  nor02 U112 ( .Y(n105), .A0(n85), .A1(n86) );
  inv01 U113 ( .Y(n95), .A(n105) );
  nor02 U114 ( .Y(n106), .A0(n88), .A1(n90) );
  inv01 U115 ( .Y(n96), .A(n106) );
  nor02 U116 ( .Y(n107), .A0(n92), .A1(n94) );
  inv01 U117 ( .Y(n97), .A(n107) );
  nor02 U118 ( .Y(n108), .A0(n98), .A1(n99) );
  inv01 U119 ( .Y(n101), .A(n108) );
  inv02 U120 ( .Y(SUM[17]), .A(n109) );
  inv02 U121 ( .Y(carry_18_), .A(n110) );
  inv02 U122 ( .Y(n111), .A(B[17]) );
  inv02 U123 ( .Y(n112), .A(A[17]) );
  inv02 U124 ( .Y(n113), .A(carry_17_) );
  nor02 U125 ( .Y(n114), .A0(n111), .A1(n115) );
  nor02 U126 ( .Y(n116), .A0(n112), .A1(n117) );
  nor02 U127 ( .Y(n118), .A0(n113), .A1(n119) );
  nor02 U128 ( .Y(n120), .A0(n113), .A1(n121) );
  nor02 U129 ( .Y(n109), .A0(n122), .A1(n123) );
  nor02 U130 ( .Y(n124), .A0(n112), .A1(n113) );
  nor02 U131 ( .Y(n125), .A0(n111), .A1(n113) );
  nor02 U132 ( .Y(n126), .A0(n111), .A1(n112) );
  nor02 U133 ( .Y(n110), .A0(n126), .A1(n127) );
  nor02 U134 ( .Y(n128), .A0(A[17]), .A1(carry_17_) );
  inv01 U135 ( .Y(n115), .A(n128) );
  nor02 U136 ( .Y(n129), .A0(B[17]), .A1(carry_17_) );
  inv01 U137 ( .Y(n117), .A(n129) );
  nor02 U138 ( .Y(n130), .A0(B[17]), .A1(A[17]) );
  inv01 U139 ( .Y(n119), .A(n130) );
  nor02 U140 ( .Y(n131), .A0(n111), .A1(n112) );
  inv01 U141 ( .Y(n121), .A(n131) );
  nor02 U142 ( .Y(n132), .A0(n114), .A1(n116) );
  inv01 U143 ( .Y(n122), .A(n132) );
  nor02 U144 ( .Y(n133), .A0(n118), .A1(n120) );
  inv01 U145 ( .Y(n123), .A(n133) );
  nor02 U146 ( .Y(n134), .A0(n124), .A1(n125) );
  inv01 U147 ( .Y(n127), .A(n134) );
  inv02 U148 ( .Y(SUM[18]), .A(n135) );
  inv02 U149 ( .Y(carry_19_), .A(n136) );
  inv02 U150 ( .Y(n137), .A(B[18]) );
  inv02 U151 ( .Y(n138), .A(A[18]) );
  inv02 U152 ( .Y(n139), .A(carry_18_) );
  nor02 U153 ( .Y(n140), .A0(n137), .A1(n141) );
  nor02 U154 ( .Y(n142), .A0(n138), .A1(n143) );
  nor02 U155 ( .Y(n144), .A0(n139), .A1(n145) );
  nor02 U156 ( .Y(n146), .A0(n139), .A1(n147) );
  nor02 U157 ( .Y(n135), .A0(n148), .A1(n149) );
  nor02 U158 ( .Y(n150), .A0(n138), .A1(n139) );
  nor02 U159 ( .Y(n151), .A0(n137), .A1(n139) );
  nor02 U160 ( .Y(n152), .A0(n137), .A1(n138) );
  nor02 U161 ( .Y(n136), .A0(n152), .A1(n153) );
  nor02 U162 ( .Y(n154), .A0(A[18]), .A1(carry_18_) );
  inv01 U163 ( .Y(n141), .A(n154) );
  nor02 U164 ( .Y(n155), .A0(B[18]), .A1(carry_18_) );
  inv01 U165 ( .Y(n143), .A(n155) );
  nor02 U166 ( .Y(n156), .A0(B[18]), .A1(A[18]) );
  inv01 U167 ( .Y(n145), .A(n156) );
  nor02 U168 ( .Y(n157), .A0(n137), .A1(n138) );
  inv01 U169 ( .Y(n147), .A(n157) );
  nor02 U170 ( .Y(n158), .A0(n140), .A1(n142) );
  inv01 U171 ( .Y(n148), .A(n158) );
  nor02 U172 ( .Y(n159), .A0(n144), .A1(n146) );
  inv01 U173 ( .Y(n149), .A(n159) );
  nor02 U174 ( .Y(n160), .A0(n150), .A1(n151) );
  inv01 U175 ( .Y(n153), .A(n160) );
  inv02 U176 ( .Y(SUM[15]), .A(n161) );
  inv02 U177 ( .Y(carry_16_), .A(n162) );
  inv02 U178 ( .Y(n163), .A(B[15]) );
  inv02 U179 ( .Y(n164), .A(A[15]) );
  inv02 U180 ( .Y(n165), .A(carry_15_) );
  nor02 U181 ( .Y(n166), .A0(n163), .A1(n167) );
  nor02 U182 ( .Y(n168), .A0(n164), .A1(n169) );
  nor02 U183 ( .Y(n170), .A0(n165), .A1(n171) );
  nor02 U184 ( .Y(n172), .A0(n165), .A1(n173) );
  nor02 U185 ( .Y(n161), .A0(n174), .A1(n175) );
  nor02 U186 ( .Y(n176), .A0(n164), .A1(n165) );
  nor02 U187 ( .Y(n177), .A0(n163), .A1(n165) );
  nor02 U188 ( .Y(n178), .A0(n163), .A1(n164) );
  nor02 U189 ( .Y(n162), .A0(n178), .A1(n179) );
  nor02 U190 ( .Y(n180), .A0(A[15]), .A1(carry_15_) );
  inv01 U191 ( .Y(n167), .A(n180) );
  nor02 U192 ( .Y(n181), .A0(B[15]), .A1(carry_15_) );
  inv01 U193 ( .Y(n169), .A(n181) );
  nor02 U194 ( .Y(n182), .A0(B[15]), .A1(A[15]) );
  inv01 U195 ( .Y(n171), .A(n182) );
  nor02 U196 ( .Y(n183), .A0(n163), .A1(n164) );
  inv01 U197 ( .Y(n173), .A(n183) );
  nor02 U198 ( .Y(n184), .A0(n166), .A1(n168) );
  inv01 U199 ( .Y(n174), .A(n184) );
  nor02 U200 ( .Y(n185), .A0(n170), .A1(n172) );
  inv01 U201 ( .Y(n175), .A(n185) );
  nor02 U202 ( .Y(n186), .A0(n176), .A1(n177) );
  inv01 U203 ( .Y(n179), .A(n186) );
  inv02 U204 ( .Y(SUM[16]), .A(n187) );
  inv02 U205 ( .Y(carry_17_), .A(n188) );
  inv02 U206 ( .Y(n189), .A(B[16]) );
  inv02 U207 ( .Y(n190), .A(A[16]) );
  inv02 U208 ( .Y(n191), .A(carry_16_) );
  nor02 U209 ( .Y(n192), .A0(n189), .A1(n193) );
  nor02 U210 ( .Y(n194), .A0(n190), .A1(n195) );
  nor02 U211 ( .Y(n196), .A0(n191), .A1(n197) );
  nor02 U212 ( .Y(n198), .A0(n191), .A1(n199) );
  nor02 U213 ( .Y(n187), .A0(n200), .A1(n201) );
  nor02 U214 ( .Y(n202), .A0(n190), .A1(n191) );
  nor02 U215 ( .Y(n203), .A0(n189), .A1(n191) );
  nor02 U216 ( .Y(n204), .A0(n189), .A1(n190) );
  nor02 U217 ( .Y(n188), .A0(n204), .A1(n205) );
  nor02 U218 ( .Y(n206), .A0(A[16]), .A1(carry_16_) );
  inv01 U219 ( .Y(n193), .A(n206) );
  nor02 U220 ( .Y(n207), .A0(B[16]), .A1(carry_16_) );
  inv01 U221 ( .Y(n195), .A(n207) );
  nor02 U222 ( .Y(n208), .A0(B[16]), .A1(A[16]) );
  inv01 U223 ( .Y(n197), .A(n208) );
  nor02 U224 ( .Y(n209), .A0(n189), .A1(n190) );
  inv01 U225 ( .Y(n199), .A(n209) );
  nor02 U226 ( .Y(n210), .A0(n192), .A1(n194) );
  inv01 U227 ( .Y(n200), .A(n210) );
  nor02 U228 ( .Y(n211), .A0(n196), .A1(n198) );
  inv01 U229 ( .Y(n201), .A(n211) );
  nor02 U230 ( .Y(n212), .A0(n202), .A1(n203) );
  inv01 U231 ( .Y(n205), .A(n212) );
  inv02 U232 ( .Y(SUM[13]), .A(n213) );
  inv02 U233 ( .Y(carry_14_), .A(n214) );
  inv02 U234 ( .Y(n215), .A(B[13]) );
  inv02 U235 ( .Y(n216), .A(A[13]) );
  inv02 U236 ( .Y(n217), .A(carry_13_) );
  nor02 U237 ( .Y(n218), .A0(n215), .A1(n219) );
  nor02 U238 ( .Y(n220), .A0(n216), .A1(n221) );
  nor02 U239 ( .Y(n222), .A0(n217), .A1(n223) );
  nor02 U240 ( .Y(n224), .A0(n217), .A1(n225) );
  nor02 U241 ( .Y(n213), .A0(n226), .A1(n227) );
  nor02 U242 ( .Y(n228), .A0(n216), .A1(n217) );
  nor02 U243 ( .Y(n229), .A0(n215), .A1(n217) );
  nor02 U244 ( .Y(n230), .A0(n215), .A1(n216) );
  nor02 U245 ( .Y(n214), .A0(n230), .A1(n231) );
  nor02 U246 ( .Y(n232), .A0(A[13]), .A1(carry_13_) );
  inv01 U247 ( .Y(n219), .A(n232) );
  nor02 U248 ( .Y(n233), .A0(B[13]), .A1(carry_13_) );
  inv01 U249 ( .Y(n221), .A(n233) );
  nor02 U250 ( .Y(n234), .A0(B[13]), .A1(A[13]) );
  inv01 U251 ( .Y(n223), .A(n234) );
  nor02 U252 ( .Y(n235), .A0(n215), .A1(n216) );
  inv01 U253 ( .Y(n225), .A(n235) );
  nor02 U254 ( .Y(n236), .A0(n218), .A1(n220) );
  inv01 U255 ( .Y(n226), .A(n236) );
  nor02 U256 ( .Y(n237), .A0(n222), .A1(n224) );
  inv01 U257 ( .Y(n227), .A(n237) );
  nor02 U258 ( .Y(n238), .A0(n228), .A1(n229) );
  inv01 U259 ( .Y(n231), .A(n238) );
  inv02 U260 ( .Y(SUM[14]), .A(n239) );
  inv02 U261 ( .Y(carry_15_), .A(n240) );
  inv02 U262 ( .Y(n241), .A(B[14]) );
  inv02 U263 ( .Y(n242), .A(A[14]) );
  inv02 U264 ( .Y(n243), .A(carry_14_) );
  nor02 U265 ( .Y(n244), .A0(n241), .A1(n245) );
  nor02 U266 ( .Y(n246), .A0(n242), .A1(n247) );
  nor02 U267 ( .Y(n248), .A0(n243), .A1(n249) );
  nor02 U268 ( .Y(n250), .A0(n243), .A1(n251) );
  nor02 U269 ( .Y(n239), .A0(n252), .A1(n253) );
  nor02 U270 ( .Y(n254), .A0(n242), .A1(n243) );
  nor02 U271 ( .Y(n255), .A0(n241), .A1(n243) );
  nor02 U272 ( .Y(n256), .A0(n241), .A1(n242) );
  nor02 U273 ( .Y(n240), .A0(n256), .A1(n257) );
  nor02 U274 ( .Y(n258), .A0(A[14]), .A1(carry_14_) );
  inv01 U275 ( .Y(n245), .A(n258) );
  nor02 U276 ( .Y(n259), .A0(B[14]), .A1(carry_14_) );
  inv01 U277 ( .Y(n247), .A(n259) );
  nor02 U278 ( .Y(n260), .A0(B[14]), .A1(A[14]) );
  inv01 U279 ( .Y(n249), .A(n260) );
  nor02 U280 ( .Y(n261), .A0(n241), .A1(n242) );
  inv01 U281 ( .Y(n251), .A(n261) );
  nor02 U282 ( .Y(n262), .A0(n244), .A1(n246) );
  inv01 U283 ( .Y(n252), .A(n262) );
  nor02 U284 ( .Y(n263), .A0(n248), .A1(n250) );
  inv01 U285 ( .Y(n253), .A(n263) );
  nor02 U286 ( .Y(n264), .A0(n254), .A1(n255) );
  inv01 U287 ( .Y(n257), .A(n264) );
  inv02 U288 ( .Y(SUM[11]), .A(n265) );
  inv02 U289 ( .Y(carry_12_), .A(n266) );
  inv02 U290 ( .Y(n267), .A(B[11]) );
  inv02 U291 ( .Y(n268), .A(A[11]) );
  inv02 U292 ( .Y(n269), .A(carry_11_) );
  nor02 U293 ( .Y(n270), .A0(n267), .A1(n271) );
  nor02 U294 ( .Y(n272), .A0(n268), .A1(n273) );
  nor02 U295 ( .Y(n274), .A0(n269), .A1(n275) );
  nor02 U296 ( .Y(n276), .A0(n269), .A1(n277) );
  nor02 U297 ( .Y(n265), .A0(n278), .A1(n279) );
  nor02 U298 ( .Y(n280), .A0(n268), .A1(n269) );
  nor02 U299 ( .Y(n281), .A0(n267), .A1(n269) );
  nor02 U300 ( .Y(n282), .A0(n267), .A1(n268) );
  nor02 U301 ( .Y(n266), .A0(n282), .A1(n283) );
  nor02 U302 ( .Y(n284), .A0(A[11]), .A1(carry_11_) );
  inv01 U303 ( .Y(n271), .A(n284) );
  nor02 U304 ( .Y(n285), .A0(B[11]), .A1(carry_11_) );
  inv01 U305 ( .Y(n273), .A(n285) );
  nor02 U306 ( .Y(n286), .A0(B[11]), .A1(A[11]) );
  inv01 U307 ( .Y(n275), .A(n286) );
  nor02 U308 ( .Y(n287), .A0(n267), .A1(n268) );
  inv01 U309 ( .Y(n277), .A(n287) );
  nor02 U310 ( .Y(n288), .A0(n270), .A1(n272) );
  inv01 U311 ( .Y(n278), .A(n288) );
  nor02 U312 ( .Y(n289), .A0(n274), .A1(n276) );
  inv01 U313 ( .Y(n279), .A(n289) );
  nor02 U314 ( .Y(n290), .A0(n280), .A1(n281) );
  inv01 U315 ( .Y(n283), .A(n290) );
  inv02 U316 ( .Y(SUM[12]), .A(n291) );
  inv02 U317 ( .Y(carry_13_), .A(n292) );
  inv02 U318 ( .Y(n293), .A(B[12]) );
  inv02 U319 ( .Y(n294), .A(A[12]) );
  inv02 U320 ( .Y(n295), .A(carry_12_) );
  nor02 U321 ( .Y(n296), .A0(n293), .A1(n297) );
  nor02 U322 ( .Y(n298), .A0(n294), .A1(n299) );
  nor02 U323 ( .Y(n300), .A0(n295), .A1(n301) );
  nor02 U324 ( .Y(n302), .A0(n295), .A1(n303) );
  nor02 U325 ( .Y(n291), .A0(n304), .A1(n305) );
  nor02 U326 ( .Y(n306), .A0(n294), .A1(n295) );
  nor02 U327 ( .Y(n307), .A0(n293), .A1(n295) );
  nor02 U328 ( .Y(n308), .A0(n293), .A1(n294) );
  nor02 U329 ( .Y(n292), .A0(n308), .A1(n309) );
  nor02 U330 ( .Y(n310), .A0(A[12]), .A1(carry_12_) );
  inv01 U331 ( .Y(n297), .A(n310) );
  nor02 U332 ( .Y(n311), .A0(B[12]), .A1(carry_12_) );
  inv01 U333 ( .Y(n299), .A(n311) );
  nor02 U334 ( .Y(n312), .A0(B[12]), .A1(A[12]) );
  inv01 U335 ( .Y(n301), .A(n312) );
  nor02 U336 ( .Y(n313), .A0(n293), .A1(n294) );
  inv01 U337 ( .Y(n303), .A(n313) );
  nor02 U338 ( .Y(n314), .A0(n296), .A1(n298) );
  inv01 U339 ( .Y(n304), .A(n314) );
  nor02 U340 ( .Y(n315), .A0(n300), .A1(n302) );
  inv01 U341 ( .Y(n305), .A(n315) );
  nor02 U342 ( .Y(n316), .A0(n306), .A1(n307) );
  inv01 U343 ( .Y(n309), .A(n316) );
  inv02 U344 ( .Y(SUM[10]), .A(n317) );
  inv02 U345 ( .Y(carry_11_), .A(n318) );
  inv02 U346 ( .Y(n319), .A(B[10]) );
  inv02 U347 ( .Y(n320), .A(A[10]) );
  inv02 U348 ( .Y(n321), .A(carry_10_) );
  nor02 U349 ( .Y(n322), .A0(n319), .A1(n323) );
  nor02 U350 ( .Y(n324), .A0(n320), .A1(n325) );
  nor02 U351 ( .Y(n326), .A0(n321), .A1(n327) );
  nor02 U352 ( .Y(n328), .A0(n321), .A1(n329) );
  nor02 U353 ( .Y(n317), .A0(n330), .A1(n331) );
  nor02 U354 ( .Y(n332), .A0(n320), .A1(n321) );
  nor02 U355 ( .Y(n333), .A0(n319), .A1(n321) );
  nor02 U356 ( .Y(n334), .A0(n319), .A1(n320) );
  nor02 U357 ( .Y(n318), .A0(n334), .A1(n335) );
  nor02 U358 ( .Y(n336), .A0(A[10]), .A1(carry_10_) );
  inv01 U359 ( .Y(n323), .A(n336) );
  nor02 U360 ( .Y(n337), .A0(B[10]), .A1(carry_10_) );
  inv01 U361 ( .Y(n325), .A(n337) );
  nor02 U362 ( .Y(n338), .A0(B[10]), .A1(A[10]) );
  inv01 U363 ( .Y(n327), .A(n338) );
  nor02 U364 ( .Y(n339), .A0(n319), .A1(n320) );
  inv01 U365 ( .Y(n329), .A(n339) );
  nor02 U366 ( .Y(n340), .A0(n322), .A1(n324) );
  inv01 U367 ( .Y(n330), .A(n340) );
  nor02 U368 ( .Y(n341), .A0(n326), .A1(n328) );
  inv01 U369 ( .Y(n331), .A(n341) );
  nor02 U370 ( .Y(n342), .A0(n332), .A1(n333) );
  inv01 U371 ( .Y(n335), .A(n342) );
  inv02 U372 ( .Y(SUM[9]), .A(n343) );
  inv02 U373 ( .Y(carry_10_), .A(n344) );
  inv02 U374 ( .Y(n345), .A(B[9]) );
  inv02 U375 ( .Y(n346), .A(A[9]) );
  inv02 U376 ( .Y(n347), .A(carry_9_) );
  nor02 U377 ( .Y(n348), .A0(n345), .A1(n349) );
  nor02 U378 ( .Y(n350), .A0(n346), .A1(n351) );
  nor02 U379 ( .Y(n352), .A0(n347), .A1(n353) );
  nor02 U380 ( .Y(n354), .A0(n347), .A1(n355) );
  nor02 U381 ( .Y(n343), .A0(n356), .A1(n357) );
  nor02 U382 ( .Y(n358), .A0(n346), .A1(n347) );
  nor02 U383 ( .Y(n359), .A0(n345), .A1(n347) );
  nor02 U384 ( .Y(n360), .A0(n345), .A1(n346) );
  nor02 U385 ( .Y(n344), .A0(n360), .A1(n361) );
  nor02 U386 ( .Y(n362), .A0(A[9]), .A1(carry_9_) );
  inv01 U387 ( .Y(n349), .A(n362) );
  nor02 U388 ( .Y(n363), .A0(B[9]), .A1(carry_9_) );
  inv01 U389 ( .Y(n351), .A(n363) );
  nor02 U390 ( .Y(n364), .A0(B[9]), .A1(A[9]) );
  inv01 U391 ( .Y(n353), .A(n364) );
  nor02 U392 ( .Y(n365), .A0(n345), .A1(n346) );
  inv01 U393 ( .Y(n355), .A(n365) );
  nor02 U394 ( .Y(n366), .A0(n348), .A1(n350) );
  inv01 U395 ( .Y(n356), .A(n366) );
  nor02 U396 ( .Y(n367), .A0(n352), .A1(n354) );
  inv01 U397 ( .Y(n357), .A(n367) );
  nor02 U398 ( .Y(n368), .A0(n358), .A1(n359) );
  inv01 U399 ( .Y(n361), .A(n368) );
  inv02 U400 ( .Y(SUM[8]), .A(n369) );
  inv02 U401 ( .Y(carry_9_), .A(n370) );
  inv02 U402 ( .Y(n371), .A(B[8]) );
  inv02 U403 ( .Y(n372), .A(A[8]) );
  inv02 U404 ( .Y(n373), .A(carry_8_) );
  nor02 U405 ( .Y(n374), .A0(n371), .A1(n375) );
  nor02 U406 ( .Y(n376), .A0(n372), .A1(n377) );
  nor02 U407 ( .Y(n378), .A0(n373), .A1(n379) );
  nor02 U408 ( .Y(n380), .A0(n373), .A1(n381) );
  nor02 U409 ( .Y(n369), .A0(n382), .A1(n383) );
  nor02 U410 ( .Y(n384), .A0(n372), .A1(n373) );
  nor02 U411 ( .Y(n385), .A0(n371), .A1(n373) );
  nor02 U412 ( .Y(n386), .A0(n371), .A1(n372) );
  nor02 U413 ( .Y(n370), .A0(n386), .A1(n387) );
  nor02 U414 ( .Y(n388), .A0(A[8]), .A1(carry_8_) );
  inv01 U415 ( .Y(n375), .A(n388) );
  nor02 U416 ( .Y(n389), .A0(B[8]), .A1(carry_8_) );
  inv01 U417 ( .Y(n377), .A(n389) );
  nor02 U418 ( .Y(n390), .A0(B[8]), .A1(A[8]) );
  inv01 U419 ( .Y(n379), .A(n390) );
  nor02 U420 ( .Y(n391), .A0(n371), .A1(n372) );
  inv01 U421 ( .Y(n381), .A(n391) );
  nor02 U422 ( .Y(n392), .A0(n374), .A1(n376) );
  inv01 U423 ( .Y(n382), .A(n392) );
  nor02 U424 ( .Y(n393), .A0(n378), .A1(n380) );
  inv01 U425 ( .Y(n383), .A(n393) );
  nor02 U426 ( .Y(n394), .A0(n384), .A1(n385) );
  inv01 U427 ( .Y(n387), .A(n394) );
  inv02 U428 ( .Y(SUM[7]), .A(n395) );
  inv02 U429 ( .Y(carry_8_), .A(n396) );
  inv02 U430 ( .Y(n397), .A(B[7]) );
  inv02 U431 ( .Y(n398), .A(A[7]) );
  inv02 U432 ( .Y(n399), .A(carry_7_) );
  nor02 U433 ( .Y(n400), .A0(n397), .A1(n401) );
  nor02 U434 ( .Y(n402), .A0(n398), .A1(n403) );
  nor02 U435 ( .Y(n404), .A0(n399), .A1(n405) );
  nor02 U436 ( .Y(n406), .A0(n399), .A1(n407) );
  nor02 U437 ( .Y(n395), .A0(n408), .A1(n409) );
  nor02 U438 ( .Y(n410), .A0(n398), .A1(n399) );
  nor02 U439 ( .Y(n411), .A0(n397), .A1(n399) );
  nor02 U440 ( .Y(n412), .A0(n397), .A1(n398) );
  nor02 U441 ( .Y(n396), .A0(n412), .A1(n413) );
  nor02 U442 ( .Y(n414), .A0(A[7]), .A1(carry_7_) );
  inv01 U443 ( .Y(n401), .A(n414) );
  nor02 U444 ( .Y(n415), .A0(B[7]), .A1(carry_7_) );
  inv01 U445 ( .Y(n403), .A(n415) );
  nor02 U446 ( .Y(n416), .A0(B[7]), .A1(A[7]) );
  inv01 U447 ( .Y(n405), .A(n416) );
  nor02 U448 ( .Y(n417), .A0(n397), .A1(n398) );
  inv01 U449 ( .Y(n407), .A(n417) );
  nor02 U450 ( .Y(n418), .A0(n400), .A1(n402) );
  inv01 U451 ( .Y(n408), .A(n418) );
  nor02 U452 ( .Y(n419), .A0(n404), .A1(n406) );
  inv01 U453 ( .Y(n409), .A(n419) );
  nor02 U454 ( .Y(n420), .A0(n410), .A1(n411) );
  inv01 U455 ( .Y(n413), .A(n420) );
  inv02 U456 ( .Y(SUM[6]), .A(n421) );
  inv02 U457 ( .Y(carry_7_), .A(n422) );
  inv02 U458 ( .Y(n423), .A(B[6]) );
  inv02 U459 ( .Y(n424), .A(A[6]) );
  inv02 U460 ( .Y(n425), .A(carry_6_) );
  nor02 U461 ( .Y(n426), .A0(n423), .A1(n427) );
  nor02 U462 ( .Y(n428), .A0(n424), .A1(n429) );
  nor02 U463 ( .Y(n430), .A0(n425), .A1(n431) );
  nor02 U464 ( .Y(n432), .A0(n425), .A1(n433) );
  nor02 U465 ( .Y(n421), .A0(n434), .A1(n435) );
  nor02 U466 ( .Y(n436), .A0(n424), .A1(n425) );
  nor02 U467 ( .Y(n437), .A0(n423), .A1(n425) );
  nor02 U468 ( .Y(n438), .A0(n423), .A1(n424) );
  nor02 U469 ( .Y(n422), .A0(n438), .A1(n439) );
  nor02 U470 ( .Y(n440), .A0(A[6]), .A1(carry_6_) );
  inv01 U471 ( .Y(n427), .A(n440) );
  nor02 U472 ( .Y(n441), .A0(B[6]), .A1(carry_6_) );
  inv01 U473 ( .Y(n429), .A(n441) );
  nor02 U474 ( .Y(n442), .A0(B[6]), .A1(A[6]) );
  inv01 U475 ( .Y(n431), .A(n442) );
  nor02 U476 ( .Y(n443), .A0(n423), .A1(n424) );
  inv01 U477 ( .Y(n433), .A(n443) );
  nor02 U478 ( .Y(n444), .A0(n426), .A1(n428) );
  inv01 U479 ( .Y(n434), .A(n444) );
  nor02 U480 ( .Y(n445), .A0(n430), .A1(n432) );
  inv01 U481 ( .Y(n435), .A(n445) );
  nor02 U482 ( .Y(n446), .A0(n436), .A1(n437) );
  inv01 U483 ( .Y(n439), .A(n446) );
  inv02 U484 ( .Y(SUM[5]), .A(n447) );
  inv02 U485 ( .Y(carry_6_), .A(n448) );
  inv02 U486 ( .Y(n449), .A(B[5]) );
  inv02 U487 ( .Y(n450), .A(A[5]) );
  inv02 U488 ( .Y(n451), .A(carry_5_) );
  nor02 U489 ( .Y(n452), .A0(n449), .A1(n453) );
  nor02 U490 ( .Y(n454), .A0(n450), .A1(n455) );
  nor02 U491 ( .Y(n456), .A0(n451), .A1(n457) );
  nor02 U492 ( .Y(n458), .A0(n451), .A1(n459) );
  nor02 U493 ( .Y(n447), .A0(n460), .A1(n461) );
  nor02 U494 ( .Y(n462), .A0(n450), .A1(n451) );
  nor02 U495 ( .Y(n463), .A0(n449), .A1(n451) );
  nor02 U496 ( .Y(n464), .A0(n449), .A1(n450) );
  nor02 U497 ( .Y(n448), .A0(n464), .A1(n465) );
  nor02 U498 ( .Y(n466), .A0(A[5]), .A1(carry_5_) );
  inv01 U499 ( .Y(n453), .A(n466) );
  nor02 U500 ( .Y(n467), .A0(B[5]), .A1(carry_5_) );
  inv01 U501 ( .Y(n455), .A(n467) );
  nor02 U502 ( .Y(n468), .A0(B[5]), .A1(A[5]) );
  inv01 U503 ( .Y(n457), .A(n468) );
  nor02 U504 ( .Y(n469), .A0(n449), .A1(n450) );
  inv01 U505 ( .Y(n459), .A(n469) );
  nor02 U506 ( .Y(n470), .A0(n452), .A1(n454) );
  inv01 U507 ( .Y(n460), .A(n470) );
  nor02 U508 ( .Y(n471), .A0(n456), .A1(n458) );
  inv01 U509 ( .Y(n461), .A(n471) );
  nor02 U510 ( .Y(n472), .A0(n462), .A1(n463) );
  inv01 U511 ( .Y(n465), .A(n472) );
  inv02 U512 ( .Y(SUM[4]), .A(n473) );
  inv02 U513 ( .Y(carry_5_), .A(n474) );
  inv02 U514 ( .Y(n475), .A(B[4]) );
  inv02 U515 ( .Y(n476), .A(A[4]) );
  inv02 U516 ( .Y(n477), .A(carry_4_) );
  nor02 U517 ( .Y(n478), .A0(n475), .A1(n479) );
  nor02 U518 ( .Y(n480), .A0(n476), .A1(n481) );
  nor02 U519 ( .Y(n482), .A0(n477), .A1(n483) );
  nor02 U520 ( .Y(n484), .A0(n477), .A1(n485) );
  nor02 U521 ( .Y(n473), .A0(n486), .A1(n487) );
  nor02 U522 ( .Y(n488), .A0(n476), .A1(n477) );
  nor02 U523 ( .Y(n489), .A0(n475), .A1(n477) );
  nor02 U524 ( .Y(n490), .A0(n475), .A1(n476) );
  nor02 U525 ( .Y(n474), .A0(n490), .A1(n491) );
  nor02 U526 ( .Y(n492), .A0(A[4]), .A1(carry_4_) );
  inv01 U527 ( .Y(n479), .A(n492) );
  nor02 U528 ( .Y(n493), .A0(B[4]), .A1(carry_4_) );
  inv01 U529 ( .Y(n481), .A(n493) );
  nor02 U530 ( .Y(n494), .A0(B[4]), .A1(A[4]) );
  inv01 U531 ( .Y(n483), .A(n494) );
  nor02 U532 ( .Y(n495), .A0(n475), .A1(n476) );
  inv01 U533 ( .Y(n485), .A(n495) );
  nor02 U534 ( .Y(n496), .A0(n478), .A1(n480) );
  inv01 U535 ( .Y(n486), .A(n496) );
  nor02 U536 ( .Y(n497), .A0(n482), .A1(n484) );
  inv01 U537 ( .Y(n487), .A(n497) );
  nor02 U538 ( .Y(n498), .A0(n488), .A1(n489) );
  inv01 U539 ( .Y(n491), .A(n498) );
  inv02 U540 ( .Y(SUM[3]), .A(n499) );
  inv02 U541 ( .Y(carry_4_), .A(n500) );
  inv02 U542 ( .Y(n501), .A(B[3]) );
  inv02 U543 ( .Y(n502), .A(A[3]) );
  inv02 U544 ( .Y(n503), .A(carry_3_) );
  nor02 U545 ( .Y(n504), .A0(n501), .A1(n505) );
  nor02 U546 ( .Y(n506), .A0(n502), .A1(n507) );
  nor02 U547 ( .Y(n508), .A0(n503), .A1(n509) );
  nor02 U548 ( .Y(n510), .A0(n503), .A1(n511) );
  nor02 U549 ( .Y(n499), .A0(n512), .A1(n513) );
  nor02 U550 ( .Y(n514), .A0(n502), .A1(n503) );
  nor02 U551 ( .Y(n515), .A0(n501), .A1(n503) );
  nor02 U552 ( .Y(n516), .A0(n501), .A1(n502) );
  nor02 U553 ( .Y(n500), .A0(n516), .A1(n517) );
  nor02 U554 ( .Y(n518), .A0(A[3]), .A1(carry_3_) );
  inv01 U555 ( .Y(n505), .A(n518) );
  nor02 U556 ( .Y(n519), .A0(B[3]), .A1(carry_3_) );
  inv01 U557 ( .Y(n507), .A(n519) );
  nor02 U558 ( .Y(n520), .A0(B[3]), .A1(A[3]) );
  inv01 U559 ( .Y(n509), .A(n520) );
  nor02 U560 ( .Y(n521), .A0(n501), .A1(n502) );
  inv01 U561 ( .Y(n511), .A(n521) );
  nor02 U562 ( .Y(n522), .A0(n504), .A1(n506) );
  inv01 U563 ( .Y(n512), .A(n522) );
  nor02 U564 ( .Y(n523), .A0(n508), .A1(n510) );
  inv01 U565 ( .Y(n513), .A(n523) );
  nor02 U566 ( .Y(n524), .A0(n514), .A1(n515) );
  inv01 U567 ( .Y(n517), .A(n524) );
  inv02 U568 ( .Y(SUM[2]), .A(n525) );
  inv02 U569 ( .Y(carry_3_), .A(n526) );
  inv02 U570 ( .Y(n527), .A(B[2]) );
  inv02 U571 ( .Y(n528), .A(A[2]) );
  inv02 U572 ( .Y(n529), .A(carry_2_) );
  nor02 U573 ( .Y(n530), .A0(n527), .A1(n531) );
  nor02 U574 ( .Y(n532), .A0(n528), .A1(n533) );
  nor02 U575 ( .Y(n534), .A0(n529), .A1(n535) );
  nor02 U576 ( .Y(n536), .A0(n529), .A1(n537) );
  nor02 U577 ( .Y(n525), .A0(n538), .A1(n539) );
  nor02 U578 ( .Y(n540), .A0(n528), .A1(n529) );
  nor02 U579 ( .Y(n541), .A0(n527), .A1(n529) );
  nor02 U580 ( .Y(n542), .A0(n527), .A1(n528) );
  nor02 U581 ( .Y(n526), .A0(n542), .A1(n543) );
  nor02 U582 ( .Y(n544), .A0(A[2]), .A1(carry_2_) );
  inv01 U583 ( .Y(n531), .A(n544) );
  nor02 U584 ( .Y(n545), .A0(B[2]), .A1(carry_2_) );
  inv01 U585 ( .Y(n533), .A(n545) );
  nor02 U586 ( .Y(n546), .A0(B[2]), .A1(A[2]) );
  inv01 U587 ( .Y(n535), .A(n546) );
  nor02 U588 ( .Y(n547), .A0(n527), .A1(n528) );
  inv01 U589 ( .Y(n537), .A(n547) );
  nor02 U590 ( .Y(n548), .A0(n530), .A1(n532) );
  inv01 U591 ( .Y(n538), .A(n548) );
  nor02 U592 ( .Y(n549), .A0(n534), .A1(n536) );
  inv01 U593 ( .Y(n539), .A(n549) );
  nor02 U594 ( .Y(n550), .A0(n540), .A1(n541) );
  inv01 U595 ( .Y(n543), .A(n550) );
  inv02 U596 ( .Y(SUM[1]), .A(n551) );
  inv02 U597 ( .Y(carry_2_), .A(n552) );
  inv02 U598 ( .Y(n553), .A(B[1]) );
  inv02 U599 ( .Y(n554), .A(A[1]) );
  inv02 U600 ( .Y(n555), .A(n3) );
  nor02 U601 ( .Y(n556), .A0(n553), .A1(n557) );
  nor02 U602 ( .Y(n558), .A0(n554), .A1(n559) );
  nor02 U603 ( .Y(n560), .A0(n555), .A1(n561) );
  nor02 U604 ( .Y(n562), .A0(n555), .A1(n563) );
  nor02 U605 ( .Y(n551), .A0(n564), .A1(n565) );
  nor02 U606 ( .Y(n566), .A0(n554), .A1(n555) );
  nor02 U607 ( .Y(n567), .A0(n553), .A1(n555) );
  nor02 U608 ( .Y(n568), .A0(n553), .A1(n554) );
  nor02 U609 ( .Y(n552), .A0(n568), .A1(n569) );
  nor02 U610 ( .Y(n570), .A0(A[1]), .A1(n3) );
  inv01 U611 ( .Y(n557), .A(n570) );
  nor02 U612 ( .Y(n571), .A0(B[1]), .A1(n3) );
  inv01 U613 ( .Y(n559), .A(n571) );
  nor02 U614 ( .Y(n572), .A0(B[1]), .A1(A[1]) );
  inv01 U615 ( .Y(n561), .A(n572) );
  nor02 U616 ( .Y(n573), .A0(n553), .A1(n554) );
  inv01 U617 ( .Y(n563), .A(n573) );
  nor02 U618 ( .Y(n574), .A0(n556), .A1(n558) );
  inv01 U619 ( .Y(n564), .A(n574) );
  nor02 U620 ( .Y(n575), .A0(n560), .A1(n562) );
  inv01 U621 ( .Y(n565), .A(n575) );
  nor02 U622 ( .Y(n576), .A0(n566), .A1(n567) );
  inv01 U623 ( .Y(n569), .A(n576) );
  xor2 U624 ( .Y(n578), .A0(B[0]), .A1(A[0]) );
  fadd1 U1_23 ( .S(n577), .A(A[23]), .B(B[23]), .CI(carry_23_) );
endmodule


module mul_24_DW01_add_24_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   carry_23_, carry_22_, carry_21_, carry_20_, carry_19_, carry_18_,
         carry_17_, carry_16_, carry_15_, carry_14_, carry_13_, carry_12_,
         carry_11_, carry_10_, carry_9_, carry_8_, carry_7_, carry_6_,
         carry_5_, carry_4_, carry_3_, carry_2_, n554, n555, n556, n557, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553;

  buf02 U4 ( .Y(SUM[0]), .A(n557) );
  nand02 U5 ( .Y(n2), .A0(A[0]), .A1(B[0]) );
  inv02 U6 ( .Y(n3), .A(n2) );
  buf02 U7 ( .Y(n4), .A(carry_23_) );
  inv01 U8 ( .Y(n556), .A(n5) );
  inv02 U9 ( .Y(carry_22_), .A(n6) );
  inv02 U10 ( .Y(n7), .A(B[21]) );
  inv02 U11 ( .Y(n8), .A(A[21]) );
  inv02 U12 ( .Y(n9), .A(carry_21_) );
  nor02 U13 ( .Y(n10), .A0(n7), .A1(n11) );
  nor02 U14 ( .Y(n12), .A0(n8), .A1(n13) );
  nor02 U15 ( .Y(n14), .A0(n9), .A1(n15) );
  nor02 U16 ( .Y(n16), .A0(n9), .A1(n17) );
  nor02 U17 ( .Y(n5), .A0(n18), .A1(n19) );
  nor02 U18 ( .Y(n20), .A0(n8), .A1(n9) );
  nor02 U19 ( .Y(n21), .A0(n7), .A1(n9) );
  nor02 U20 ( .Y(n22), .A0(n7), .A1(n8) );
  nor02 U21 ( .Y(n6), .A0(n22), .A1(n23) );
  nor02 U22 ( .Y(n24), .A0(A[21]), .A1(carry_21_) );
  inv01 U23 ( .Y(n11), .A(n24) );
  nor02 U24 ( .Y(n25), .A0(B[21]), .A1(carry_21_) );
  inv01 U25 ( .Y(n13), .A(n25) );
  nor02 U26 ( .Y(n26), .A0(B[21]), .A1(A[21]) );
  inv01 U27 ( .Y(n15), .A(n26) );
  nor02 U28 ( .Y(n27), .A0(n7), .A1(n8) );
  inv01 U29 ( .Y(n17), .A(n27) );
  nor02 U30 ( .Y(n28), .A0(n10), .A1(n12) );
  inv01 U31 ( .Y(n18), .A(n28) );
  nor02 U32 ( .Y(n29), .A0(n14), .A1(n16) );
  inv01 U33 ( .Y(n19), .A(n29) );
  nor02 U34 ( .Y(n30), .A0(n20), .A1(n21) );
  inv01 U35 ( .Y(n23), .A(n30) );
  buf02 U36 ( .Y(SUM[23]), .A(n554) );
  inv02 U37 ( .Y(SUM[20]), .A(n32) );
  inv02 U38 ( .Y(carry_21_), .A(n33) );
  inv02 U39 ( .Y(n34), .A(B[20]) );
  inv02 U40 ( .Y(n35), .A(A[20]) );
  inv02 U41 ( .Y(n36), .A(carry_20_) );
  nor02 U42 ( .Y(n37), .A0(n34), .A1(n38) );
  nor02 U43 ( .Y(n39), .A0(n35), .A1(n40) );
  nor02 U44 ( .Y(n41), .A0(n36), .A1(n42) );
  nor02 U45 ( .Y(n43), .A0(n36), .A1(n44) );
  nor02 U46 ( .Y(n32), .A0(n45), .A1(n46) );
  nor02 U47 ( .Y(n47), .A0(n35), .A1(n36) );
  nor02 U48 ( .Y(n48), .A0(n34), .A1(n36) );
  nor02 U49 ( .Y(n49), .A0(n34), .A1(n35) );
  nor02 U50 ( .Y(n33), .A0(n49), .A1(n50) );
  nor02 U51 ( .Y(n51), .A0(A[20]), .A1(carry_20_) );
  inv01 U52 ( .Y(n38), .A(n51) );
  nor02 U53 ( .Y(n52), .A0(B[20]), .A1(carry_20_) );
  inv01 U54 ( .Y(n40), .A(n52) );
  nor02 U55 ( .Y(n53), .A0(B[20]), .A1(A[20]) );
  inv01 U56 ( .Y(n42), .A(n53) );
  nor02 U57 ( .Y(n54), .A0(n34), .A1(n35) );
  inv01 U58 ( .Y(n44), .A(n54) );
  nor02 U59 ( .Y(n55), .A0(n37), .A1(n39) );
  inv01 U60 ( .Y(n45), .A(n55) );
  nor02 U61 ( .Y(n56), .A0(n41), .A1(n43) );
  inv01 U62 ( .Y(n46), .A(n56) );
  nor02 U63 ( .Y(n57), .A0(n47), .A1(n48) );
  inv01 U64 ( .Y(n50), .A(n57) );
  buf02 U65 ( .Y(SUM[22]), .A(n555) );
  inv02 U66 ( .Y(SUM[18]), .A(n59) );
  inv02 U67 ( .Y(carry_19_), .A(n60) );
  inv02 U68 ( .Y(n61), .A(B[18]) );
  inv02 U69 ( .Y(n62), .A(A[18]) );
  inv02 U70 ( .Y(n63), .A(carry_18_) );
  nor02 U71 ( .Y(n64), .A0(n61), .A1(n65) );
  nor02 U72 ( .Y(n66), .A0(n62), .A1(n67) );
  nor02 U73 ( .Y(n68), .A0(n63), .A1(n69) );
  nor02 U74 ( .Y(n70), .A0(n63), .A1(n71) );
  nor02 U75 ( .Y(n59), .A0(n72), .A1(n73) );
  nor02 U76 ( .Y(n74), .A0(n62), .A1(n63) );
  nor02 U77 ( .Y(n75), .A0(n61), .A1(n63) );
  nor02 U78 ( .Y(n76), .A0(n61), .A1(n62) );
  nor02 U79 ( .Y(n60), .A0(n76), .A1(n77) );
  nor02 U80 ( .Y(n78), .A0(A[18]), .A1(carry_18_) );
  inv01 U81 ( .Y(n65), .A(n78) );
  nor02 U82 ( .Y(n79), .A0(B[18]), .A1(carry_18_) );
  inv01 U83 ( .Y(n67), .A(n79) );
  nor02 U84 ( .Y(n80), .A0(B[18]), .A1(A[18]) );
  inv01 U85 ( .Y(n69), .A(n80) );
  nor02 U86 ( .Y(n81), .A0(n61), .A1(n62) );
  inv01 U87 ( .Y(n71), .A(n81) );
  nor02 U88 ( .Y(n82), .A0(n64), .A1(n66) );
  inv01 U89 ( .Y(n72), .A(n82) );
  nor02 U90 ( .Y(n83), .A0(n68), .A1(n70) );
  inv01 U91 ( .Y(n73), .A(n83) );
  nor02 U92 ( .Y(n84), .A0(n74), .A1(n75) );
  inv01 U93 ( .Y(n77), .A(n84) );
  inv02 U94 ( .Y(SUM[19]), .A(n85) );
  inv02 U95 ( .Y(carry_20_), .A(n86) );
  inv02 U96 ( .Y(n87), .A(B[19]) );
  inv02 U97 ( .Y(n88), .A(A[19]) );
  inv02 U98 ( .Y(n89), .A(carry_19_) );
  nor02 U99 ( .Y(n90), .A0(n87), .A1(n91) );
  nor02 U100 ( .Y(n92), .A0(n88), .A1(n93) );
  nor02 U101 ( .Y(n94), .A0(n89), .A1(n95) );
  nor02 U102 ( .Y(n96), .A0(n89), .A1(n97) );
  nor02 U103 ( .Y(n85), .A0(n98), .A1(n99) );
  nor02 U104 ( .Y(n100), .A0(n88), .A1(n89) );
  nor02 U105 ( .Y(n101), .A0(n87), .A1(n89) );
  nor02 U106 ( .Y(n102), .A0(n87), .A1(n88) );
  nor02 U107 ( .Y(n86), .A0(n102), .A1(n103) );
  nor02 U108 ( .Y(n104), .A0(A[19]), .A1(carry_19_) );
  inv01 U109 ( .Y(n91), .A(n104) );
  nor02 U110 ( .Y(n105), .A0(B[19]), .A1(carry_19_) );
  inv01 U111 ( .Y(n93), .A(n105) );
  nor02 U112 ( .Y(n106), .A0(B[19]), .A1(A[19]) );
  inv01 U113 ( .Y(n95), .A(n106) );
  nor02 U114 ( .Y(n107), .A0(n87), .A1(n88) );
  inv01 U115 ( .Y(n97), .A(n107) );
  nor02 U116 ( .Y(n108), .A0(n90), .A1(n92) );
  inv01 U117 ( .Y(n98), .A(n108) );
  nor02 U118 ( .Y(n109), .A0(n94), .A1(n96) );
  inv01 U119 ( .Y(n99), .A(n109) );
  nor02 U120 ( .Y(n110), .A0(n100), .A1(n101) );
  inv01 U121 ( .Y(n103), .A(n110) );
  inv02 U122 ( .Y(SUM[16]), .A(n111) );
  inv02 U123 ( .Y(carry_17_), .A(n112) );
  inv02 U124 ( .Y(n113), .A(B[16]) );
  inv02 U125 ( .Y(n114), .A(A[16]) );
  inv02 U126 ( .Y(n115), .A(carry_16_) );
  nor02 U127 ( .Y(n116), .A0(n113), .A1(n117) );
  nor02 U128 ( .Y(n118), .A0(n114), .A1(n119) );
  nor02 U129 ( .Y(n120), .A0(n115), .A1(n121) );
  nor02 U130 ( .Y(n122), .A0(n115), .A1(n123) );
  nor02 U131 ( .Y(n111), .A0(n124), .A1(n125) );
  nor02 U132 ( .Y(n126), .A0(n114), .A1(n115) );
  nor02 U133 ( .Y(n127), .A0(n113), .A1(n115) );
  nor02 U134 ( .Y(n128), .A0(n113), .A1(n114) );
  nor02 U135 ( .Y(n112), .A0(n128), .A1(n129) );
  nor02 U136 ( .Y(n130), .A0(A[16]), .A1(carry_16_) );
  inv01 U137 ( .Y(n117), .A(n130) );
  nor02 U138 ( .Y(n131), .A0(B[16]), .A1(carry_16_) );
  inv01 U139 ( .Y(n119), .A(n131) );
  nor02 U140 ( .Y(n132), .A0(B[16]), .A1(A[16]) );
  inv01 U141 ( .Y(n121), .A(n132) );
  nor02 U142 ( .Y(n133), .A0(n113), .A1(n114) );
  inv01 U143 ( .Y(n123), .A(n133) );
  nor02 U144 ( .Y(n134), .A0(n116), .A1(n118) );
  inv01 U145 ( .Y(n124), .A(n134) );
  nor02 U146 ( .Y(n135), .A0(n120), .A1(n122) );
  inv01 U147 ( .Y(n125), .A(n135) );
  nor02 U148 ( .Y(n136), .A0(n126), .A1(n127) );
  inv01 U149 ( .Y(n129), .A(n136) );
  inv02 U150 ( .Y(SUM[17]), .A(n137) );
  inv02 U151 ( .Y(carry_18_), .A(n138) );
  inv02 U152 ( .Y(n139), .A(B[17]) );
  inv02 U153 ( .Y(n140), .A(A[17]) );
  inv02 U154 ( .Y(n141), .A(carry_17_) );
  nor02 U155 ( .Y(n142), .A0(n139), .A1(n143) );
  nor02 U156 ( .Y(n144), .A0(n140), .A1(n145) );
  nor02 U157 ( .Y(n146), .A0(n141), .A1(n147) );
  nor02 U158 ( .Y(n148), .A0(n141), .A1(n149) );
  nor02 U159 ( .Y(n137), .A0(n150), .A1(n151) );
  nor02 U160 ( .Y(n152), .A0(n140), .A1(n141) );
  nor02 U161 ( .Y(n153), .A0(n139), .A1(n141) );
  nor02 U162 ( .Y(n154), .A0(n139), .A1(n140) );
  nor02 U163 ( .Y(n138), .A0(n154), .A1(n155) );
  nor02 U164 ( .Y(n156), .A0(A[17]), .A1(carry_17_) );
  inv01 U165 ( .Y(n143), .A(n156) );
  nor02 U166 ( .Y(n157), .A0(B[17]), .A1(carry_17_) );
  inv01 U167 ( .Y(n145), .A(n157) );
  nor02 U168 ( .Y(n158), .A0(B[17]), .A1(A[17]) );
  inv01 U169 ( .Y(n147), .A(n158) );
  nor02 U170 ( .Y(n159), .A0(n139), .A1(n140) );
  inv01 U171 ( .Y(n149), .A(n159) );
  nor02 U172 ( .Y(n160), .A0(n142), .A1(n144) );
  inv01 U173 ( .Y(n150), .A(n160) );
  nor02 U174 ( .Y(n161), .A0(n146), .A1(n148) );
  inv01 U175 ( .Y(n151), .A(n161) );
  nor02 U176 ( .Y(n162), .A0(n152), .A1(n153) );
  inv01 U177 ( .Y(n155), .A(n162) );
  inv02 U178 ( .Y(SUM[14]), .A(n163) );
  inv02 U179 ( .Y(carry_15_), .A(n164) );
  inv02 U180 ( .Y(n165), .A(B[14]) );
  inv02 U181 ( .Y(n166), .A(A[14]) );
  inv02 U182 ( .Y(n167), .A(carry_14_) );
  nor02 U183 ( .Y(n168), .A0(n165), .A1(n169) );
  nor02 U184 ( .Y(n170), .A0(n166), .A1(n171) );
  nor02 U185 ( .Y(n172), .A0(n167), .A1(n173) );
  nor02 U186 ( .Y(n174), .A0(n167), .A1(n175) );
  nor02 U187 ( .Y(n163), .A0(n176), .A1(n177) );
  nor02 U188 ( .Y(n178), .A0(n166), .A1(n167) );
  nor02 U189 ( .Y(n179), .A0(n165), .A1(n167) );
  nor02 U190 ( .Y(n180), .A0(n165), .A1(n166) );
  nor02 U191 ( .Y(n164), .A0(n180), .A1(n181) );
  nor02 U192 ( .Y(n182), .A0(A[14]), .A1(carry_14_) );
  inv01 U193 ( .Y(n169), .A(n182) );
  nor02 U194 ( .Y(n183), .A0(B[14]), .A1(carry_14_) );
  inv01 U195 ( .Y(n171), .A(n183) );
  nor02 U196 ( .Y(n184), .A0(B[14]), .A1(A[14]) );
  inv01 U197 ( .Y(n173), .A(n184) );
  nor02 U198 ( .Y(n185), .A0(n165), .A1(n166) );
  inv01 U199 ( .Y(n175), .A(n185) );
  nor02 U200 ( .Y(n186), .A0(n168), .A1(n170) );
  inv01 U201 ( .Y(n176), .A(n186) );
  nor02 U202 ( .Y(n187), .A0(n172), .A1(n174) );
  inv01 U203 ( .Y(n177), .A(n187) );
  nor02 U204 ( .Y(n188), .A0(n178), .A1(n179) );
  inv01 U205 ( .Y(n181), .A(n188) );
  inv02 U206 ( .Y(SUM[15]), .A(n189) );
  inv02 U207 ( .Y(carry_16_), .A(n190) );
  inv02 U208 ( .Y(n191), .A(B[15]) );
  inv02 U209 ( .Y(n192), .A(A[15]) );
  inv02 U210 ( .Y(n193), .A(carry_15_) );
  nor02 U211 ( .Y(n194), .A0(n191), .A1(n195) );
  nor02 U212 ( .Y(n196), .A0(n192), .A1(n197) );
  nor02 U213 ( .Y(n198), .A0(n193), .A1(n199) );
  nor02 U214 ( .Y(n200), .A0(n193), .A1(n201) );
  nor02 U215 ( .Y(n189), .A0(n202), .A1(n203) );
  nor02 U216 ( .Y(n204), .A0(n192), .A1(n193) );
  nor02 U217 ( .Y(n205), .A0(n191), .A1(n193) );
  nor02 U218 ( .Y(n206), .A0(n191), .A1(n192) );
  nor02 U219 ( .Y(n190), .A0(n206), .A1(n207) );
  nor02 U220 ( .Y(n208), .A0(A[15]), .A1(carry_15_) );
  inv01 U221 ( .Y(n195), .A(n208) );
  nor02 U222 ( .Y(n209), .A0(B[15]), .A1(carry_15_) );
  inv01 U223 ( .Y(n197), .A(n209) );
  nor02 U224 ( .Y(n210), .A0(B[15]), .A1(A[15]) );
  inv01 U225 ( .Y(n199), .A(n210) );
  nor02 U226 ( .Y(n211), .A0(n191), .A1(n192) );
  inv01 U227 ( .Y(n201), .A(n211) );
  nor02 U228 ( .Y(n212), .A0(n194), .A1(n196) );
  inv01 U229 ( .Y(n202), .A(n212) );
  nor02 U230 ( .Y(n213), .A0(n198), .A1(n200) );
  inv01 U231 ( .Y(n203), .A(n213) );
  nor02 U232 ( .Y(n214), .A0(n204), .A1(n205) );
  inv01 U233 ( .Y(n207), .A(n214) );
  inv02 U234 ( .Y(SUM[12]), .A(n215) );
  inv02 U235 ( .Y(carry_13_), .A(n216) );
  inv02 U236 ( .Y(n217), .A(B[12]) );
  inv02 U237 ( .Y(n218), .A(A[12]) );
  inv02 U238 ( .Y(n219), .A(carry_12_) );
  nor02 U239 ( .Y(n220), .A0(n217), .A1(n221) );
  nor02 U240 ( .Y(n222), .A0(n218), .A1(n223) );
  nor02 U241 ( .Y(n224), .A0(n219), .A1(n225) );
  nor02 U242 ( .Y(n226), .A0(n219), .A1(n227) );
  nor02 U243 ( .Y(n215), .A0(n228), .A1(n229) );
  nor02 U244 ( .Y(n230), .A0(n218), .A1(n219) );
  nor02 U245 ( .Y(n231), .A0(n217), .A1(n219) );
  nor02 U246 ( .Y(n232), .A0(n217), .A1(n218) );
  nor02 U247 ( .Y(n216), .A0(n232), .A1(n233) );
  nor02 U248 ( .Y(n234), .A0(A[12]), .A1(carry_12_) );
  inv01 U249 ( .Y(n221), .A(n234) );
  nor02 U250 ( .Y(n235), .A0(B[12]), .A1(carry_12_) );
  inv01 U251 ( .Y(n223), .A(n235) );
  nor02 U252 ( .Y(n236), .A0(B[12]), .A1(A[12]) );
  inv01 U253 ( .Y(n225), .A(n236) );
  nor02 U254 ( .Y(n237), .A0(n217), .A1(n218) );
  inv01 U255 ( .Y(n227), .A(n237) );
  nor02 U256 ( .Y(n238), .A0(n220), .A1(n222) );
  inv01 U257 ( .Y(n228), .A(n238) );
  nor02 U258 ( .Y(n239), .A0(n224), .A1(n226) );
  inv01 U259 ( .Y(n229), .A(n239) );
  nor02 U260 ( .Y(n240), .A0(n230), .A1(n231) );
  inv01 U261 ( .Y(n233), .A(n240) );
  inv02 U262 ( .Y(SUM[13]), .A(n241) );
  inv02 U263 ( .Y(carry_14_), .A(n242) );
  inv02 U264 ( .Y(n243), .A(B[13]) );
  inv02 U265 ( .Y(n244), .A(A[13]) );
  inv02 U266 ( .Y(n245), .A(carry_13_) );
  nor02 U267 ( .Y(n246), .A0(n243), .A1(n247) );
  nor02 U268 ( .Y(n248), .A0(n244), .A1(n249) );
  nor02 U269 ( .Y(n250), .A0(n245), .A1(n251) );
  nor02 U270 ( .Y(n252), .A0(n245), .A1(n253) );
  nor02 U271 ( .Y(n241), .A0(n254), .A1(n255) );
  nor02 U272 ( .Y(n256), .A0(n244), .A1(n245) );
  nor02 U273 ( .Y(n257), .A0(n243), .A1(n245) );
  nor02 U274 ( .Y(n258), .A0(n243), .A1(n244) );
  nor02 U275 ( .Y(n242), .A0(n258), .A1(n259) );
  nor02 U276 ( .Y(n260), .A0(A[13]), .A1(carry_13_) );
  inv01 U277 ( .Y(n247), .A(n260) );
  nor02 U278 ( .Y(n261), .A0(B[13]), .A1(carry_13_) );
  inv01 U279 ( .Y(n249), .A(n261) );
  nor02 U280 ( .Y(n262), .A0(B[13]), .A1(A[13]) );
  inv01 U281 ( .Y(n251), .A(n262) );
  nor02 U282 ( .Y(n263), .A0(n243), .A1(n244) );
  inv01 U283 ( .Y(n253), .A(n263) );
  nor02 U284 ( .Y(n264), .A0(n246), .A1(n248) );
  inv01 U285 ( .Y(n254), .A(n264) );
  nor02 U286 ( .Y(n265), .A0(n250), .A1(n252) );
  inv01 U287 ( .Y(n255), .A(n265) );
  nor02 U288 ( .Y(n266), .A0(n256), .A1(n257) );
  inv01 U289 ( .Y(n259), .A(n266) );
  buf02 U290 ( .Y(SUM[21]), .A(n556) );
  inv02 U291 ( .Y(SUM[10]), .A(n268) );
  inv02 U292 ( .Y(carry_11_), .A(n269) );
  inv02 U293 ( .Y(n270), .A(B[10]) );
  inv02 U294 ( .Y(n271), .A(A[10]) );
  inv02 U295 ( .Y(n272), .A(carry_10_) );
  nor02 U296 ( .Y(n273), .A0(n270), .A1(n274) );
  nor02 U297 ( .Y(n275), .A0(n271), .A1(n276) );
  nor02 U298 ( .Y(n277), .A0(n272), .A1(n278) );
  nor02 U299 ( .Y(n279), .A0(n272), .A1(n280) );
  nor02 U300 ( .Y(n268), .A0(n281), .A1(n282) );
  nor02 U301 ( .Y(n283), .A0(n271), .A1(n272) );
  nor02 U302 ( .Y(n284), .A0(n270), .A1(n272) );
  nor02 U303 ( .Y(n285), .A0(n270), .A1(n271) );
  nor02 U304 ( .Y(n269), .A0(n285), .A1(n286) );
  nor02 U305 ( .Y(n287), .A0(A[10]), .A1(carry_10_) );
  inv01 U306 ( .Y(n274), .A(n287) );
  nor02 U307 ( .Y(n288), .A0(B[10]), .A1(carry_10_) );
  inv01 U308 ( .Y(n276), .A(n288) );
  nor02 U309 ( .Y(n289), .A0(B[10]), .A1(A[10]) );
  inv01 U310 ( .Y(n278), .A(n289) );
  nor02 U311 ( .Y(n290), .A0(n270), .A1(n271) );
  inv01 U312 ( .Y(n280), .A(n290) );
  nor02 U313 ( .Y(n291), .A0(n273), .A1(n275) );
  inv01 U314 ( .Y(n281), .A(n291) );
  nor02 U315 ( .Y(n292), .A0(n277), .A1(n279) );
  inv01 U316 ( .Y(n282), .A(n292) );
  nor02 U317 ( .Y(n293), .A0(n283), .A1(n284) );
  inv01 U318 ( .Y(n286), .A(n293) );
  inv02 U319 ( .Y(SUM[11]), .A(n294) );
  inv02 U320 ( .Y(carry_12_), .A(n295) );
  inv02 U321 ( .Y(n296), .A(B[11]) );
  inv02 U322 ( .Y(n297), .A(A[11]) );
  inv02 U323 ( .Y(n298), .A(carry_11_) );
  nor02 U324 ( .Y(n299), .A0(n296), .A1(n300) );
  nor02 U325 ( .Y(n301), .A0(n297), .A1(n302) );
  nor02 U326 ( .Y(n303), .A0(n298), .A1(n304) );
  nor02 U327 ( .Y(n305), .A0(n298), .A1(n306) );
  nor02 U328 ( .Y(n294), .A0(n307), .A1(n308) );
  nor02 U329 ( .Y(n309), .A0(n297), .A1(n298) );
  nor02 U330 ( .Y(n310), .A0(n296), .A1(n298) );
  nor02 U331 ( .Y(n311), .A0(n296), .A1(n297) );
  nor02 U332 ( .Y(n295), .A0(n311), .A1(n312) );
  nor02 U333 ( .Y(n313), .A0(A[11]), .A1(carry_11_) );
  inv01 U334 ( .Y(n300), .A(n313) );
  nor02 U335 ( .Y(n314), .A0(B[11]), .A1(carry_11_) );
  inv01 U336 ( .Y(n302), .A(n314) );
  nor02 U337 ( .Y(n315), .A0(B[11]), .A1(A[11]) );
  inv01 U338 ( .Y(n304), .A(n315) );
  nor02 U339 ( .Y(n316), .A0(n296), .A1(n297) );
  inv01 U340 ( .Y(n306), .A(n316) );
  nor02 U341 ( .Y(n317), .A0(n299), .A1(n301) );
  inv01 U342 ( .Y(n307), .A(n317) );
  nor02 U343 ( .Y(n318), .A0(n303), .A1(n305) );
  inv01 U344 ( .Y(n308), .A(n318) );
  nor02 U345 ( .Y(n319), .A0(n309), .A1(n310) );
  inv01 U346 ( .Y(n312), .A(n319) );
  inv02 U347 ( .Y(SUM[9]), .A(n320) );
  inv02 U348 ( .Y(carry_10_), .A(n321) );
  inv02 U349 ( .Y(n322), .A(B[9]) );
  inv02 U350 ( .Y(n323), .A(A[9]) );
  inv02 U351 ( .Y(n324), .A(carry_9_) );
  nor02 U352 ( .Y(n325), .A0(n322), .A1(n326) );
  nor02 U353 ( .Y(n327), .A0(n323), .A1(n328) );
  nor02 U354 ( .Y(n329), .A0(n324), .A1(n330) );
  nor02 U355 ( .Y(n331), .A0(n324), .A1(n332) );
  nor02 U356 ( .Y(n320), .A0(n333), .A1(n334) );
  nor02 U357 ( .Y(n335), .A0(n323), .A1(n324) );
  nor02 U358 ( .Y(n336), .A0(n322), .A1(n324) );
  nor02 U359 ( .Y(n337), .A0(n322), .A1(n323) );
  nor02 U360 ( .Y(n321), .A0(n337), .A1(n338) );
  nor02 U361 ( .Y(n339), .A0(A[9]), .A1(carry_9_) );
  inv01 U362 ( .Y(n326), .A(n339) );
  nor02 U363 ( .Y(n340), .A0(B[9]), .A1(carry_9_) );
  inv01 U364 ( .Y(n328), .A(n340) );
  nor02 U365 ( .Y(n341), .A0(B[9]), .A1(A[9]) );
  inv01 U366 ( .Y(n330), .A(n341) );
  nor02 U367 ( .Y(n342), .A0(n322), .A1(n323) );
  inv01 U368 ( .Y(n332), .A(n342) );
  nor02 U369 ( .Y(n343), .A0(n325), .A1(n327) );
  inv01 U370 ( .Y(n333), .A(n343) );
  nor02 U371 ( .Y(n344), .A0(n329), .A1(n331) );
  inv01 U372 ( .Y(n334), .A(n344) );
  nor02 U373 ( .Y(n345), .A0(n335), .A1(n336) );
  inv01 U374 ( .Y(n338), .A(n345) );
  inv02 U375 ( .Y(SUM[8]), .A(n346) );
  inv02 U376 ( .Y(carry_9_), .A(n347) );
  inv02 U377 ( .Y(n348), .A(B[8]) );
  inv02 U378 ( .Y(n349), .A(A[8]) );
  inv02 U379 ( .Y(n350), .A(carry_8_) );
  nor02 U380 ( .Y(n351), .A0(n348), .A1(n352) );
  nor02 U381 ( .Y(n353), .A0(n349), .A1(n354) );
  nor02 U382 ( .Y(n355), .A0(n350), .A1(n356) );
  nor02 U383 ( .Y(n357), .A0(n350), .A1(n358) );
  nor02 U384 ( .Y(n346), .A0(n359), .A1(n360) );
  nor02 U385 ( .Y(n361), .A0(n349), .A1(n350) );
  nor02 U386 ( .Y(n362), .A0(n348), .A1(n350) );
  nor02 U387 ( .Y(n363), .A0(n348), .A1(n349) );
  nor02 U388 ( .Y(n347), .A0(n363), .A1(n364) );
  nor02 U389 ( .Y(n365), .A0(A[8]), .A1(carry_8_) );
  inv01 U390 ( .Y(n352), .A(n365) );
  nor02 U391 ( .Y(n366), .A0(B[8]), .A1(carry_8_) );
  inv01 U392 ( .Y(n354), .A(n366) );
  nor02 U393 ( .Y(n367), .A0(B[8]), .A1(A[8]) );
  inv01 U394 ( .Y(n356), .A(n367) );
  nor02 U395 ( .Y(n368), .A0(n348), .A1(n349) );
  inv01 U396 ( .Y(n358), .A(n368) );
  nor02 U397 ( .Y(n369), .A0(n351), .A1(n353) );
  inv01 U398 ( .Y(n359), .A(n369) );
  nor02 U399 ( .Y(n370), .A0(n355), .A1(n357) );
  inv01 U400 ( .Y(n360), .A(n370) );
  nor02 U401 ( .Y(n371), .A0(n361), .A1(n362) );
  inv01 U402 ( .Y(n364), .A(n371) );
  inv02 U403 ( .Y(SUM[7]), .A(n372) );
  inv02 U404 ( .Y(carry_8_), .A(n373) );
  inv02 U405 ( .Y(n374), .A(B[7]) );
  inv02 U406 ( .Y(n375), .A(A[7]) );
  inv02 U407 ( .Y(n376), .A(carry_7_) );
  nor02 U408 ( .Y(n377), .A0(n374), .A1(n378) );
  nor02 U409 ( .Y(n379), .A0(n375), .A1(n380) );
  nor02 U410 ( .Y(n381), .A0(n376), .A1(n382) );
  nor02 U411 ( .Y(n383), .A0(n376), .A1(n384) );
  nor02 U412 ( .Y(n372), .A0(n385), .A1(n386) );
  nor02 U413 ( .Y(n387), .A0(n375), .A1(n376) );
  nor02 U414 ( .Y(n388), .A0(n374), .A1(n376) );
  nor02 U415 ( .Y(n389), .A0(n374), .A1(n375) );
  nor02 U416 ( .Y(n373), .A0(n389), .A1(n390) );
  nor02 U417 ( .Y(n391), .A0(A[7]), .A1(carry_7_) );
  inv01 U418 ( .Y(n378), .A(n391) );
  nor02 U419 ( .Y(n392), .A0(B[7]), .A1(carry_7_) );
  inv01 U420 ( .Y(n380), .A(n392) );
  nor02 U421 ( .Y(n393), .A0(B[7]), .A1(A[7]) );
  inv01 U422 ( .Y(n382), .A(n393) );
  nor02 U423 ( .Y(n394), .A0(n374), .A1(n375) );
  inv01 U424 ( .Y(n384), .A(n394) );
  nor02 U425 ( .Y(n395), .A0(n377), .A1(n379) );
  inv01 U426 ( .Y(n385), .A(n395) );
  nor02 U427 ( .Y(n396), .A0(n381), .A1(n383) );
  inv01 U428 ( .Y(n386), .A(n396) );
  nor02 U429 ( .Y(n397), .A0(n387), .A1(n388) );
  inv01 U430 ( .Y(n390), .A(n397) );
  inv02 U431 ( .Y(SUM[6]), .A(n398) );
  inv02 U432 ( .Y(carry_7_), .A(n399) );
  inv02 U433 ( .Y(n400), .A(B[6]) );
  inv02 U434 ( .Y(n401), .A(A[6]) );
  inv02 U435 ( .Y(n402), .A(carry_6_) );
  nor02 U436 ( .Y(n403), .A0(n400), .A1(n404) );
  nor02 U437 ( .Y(n405), .A0(n401), .A1(n406) );
  nor02 U438 ( .Y(n407), .A0(n402), .A1(n408) );
  nor02 U439 ( .Y(n409), .A0(n402), .A1(n410) );
  nor02 U440 ( .Y(n398), .A0(n411), .A1(n412) );
  nor02 U441 ( .Y(n413), .A0(n401), .A1(n402) );
  nor02 U442 ( .Y(n414), .A0(n400), .A1(n402) );
  nor02 U443 ( .Y(n415), .A0(n400), .A1(n401) );
  nor02 U444 ( .Y(n399), .A0(n415), .A1(n416) );
  nor02 U445 ( .Y(n417), .A0(A[6]), .A1(carry_6_) );
  inv01 U446 ( .Y(n404), .A(n417) );
  nor02 U447 ( .Y(n418), .A0(B[6]), .A1(carry_6_) );
  inv01 U448 ( .Y(n406), .A(n418) );
  nor02 U449 ( .Y(n419), .A0(B[6]), .A1(A[6]) );
  inv01 U450 ( .Y(n408), .A(n419) );
  nor02 U451 ( .Y(n420), .A0(n400), .A1(n401) );
  inv01 U452 ( .Y(n410), .A(n420) );
  nor02 U453 ( .Y(n421), .A0(n403), .A1(n405) );
  inv01 U454 ( .Y(n411), .A(n421) );
  nor02 U455 ( .Y(n422), .A0(n407), .A1(n409) );
  inv01 U456 ( .Y(n412), .A(n422) );
  nor02 U457 ( .Y(n423), .A0(n413), .A1(n414) );
  inv01 U458 ( .Y(n416), .A(n423) );
  inv02 U459 ( .Y(SUM[5]), .A(n424) );
  inv02 U460 ( .Y(carry_6_), .A(n425) );
  inv02 U461 ( .Y(n426), .A(B[5]) );
  inv02 U462 ( .Y(n427), .A(A[5]) );
  inv02 U463 ( .Y(n428), .A(carry_5_) );
  nor02 U464 ( .Y(n429), .A0(n426), .A1(n430) );
  nor02 U465 ( .Y(n431), .A0(n427), .A1(n432) );
  nor02 U466 ( .Y(n433), .A0(n428), .A1(n434) );
  nor02 U467 ( .Y(n435), .A0(n428), .A1(n436) );
  nor02 U468 ( .Y(n424), .A0(n437), .A1(n438) );
  nor02 U469 ( .Y(n439), .A0(n427), .A1(n428) );
  nor02 U470 ( .Y(n440), .A0(n426), .A1(n428) );
  nor02 U471 ( .Y(n441), .A0(n426), .A1(n427) );
  nor02 U472 ( .Y(n425), .A0(n441), .A1(n442) );
  nor02 U473 ( .Y(n443), .A0(A[5]), .A1(carry_5_) );
  inv01 U474 ( .Y(n430), .A(n443) );
  nor02 U475 ( .Y(n444), .A0(B[5]), .A1(carry_5_) );
  inv01 U476 ( .Y(n432), .A(n444) );
  nor02 U477 ( .Y(n445), .A0(B[5]), .A1(A[5]) );
  inv01 U478 ( .Y(n434), .A(n445) );
  nor02 U479 ( .Y(n446), .A0(n426), .A1(n427) );
  inv01 U480 ( .Y(n436), .A(n446) );
  nor02 U481 ( .Y(n447), .A0(n429), .A1(n431) );
  inv01 U482 ( .Y(n437), .A(n447) );
  nor02 U483 ( .Y(n448), .A0(n433), .A1(n435) );
  inv01 U484 ( .Y(n438), .A(n448) );
  nor02 U485 ( .Y(n449), .A0(n439), .A1(n440) );
  inv01 U486 ( .Y(n442), .A(n449) );
  inv02 U487 ( .Y(SUM[4]), .A(n450) );
  inv02 U488 ( .Y(carry_5_), .A(n451) );
  inv02 U489 ( .Y(n452), .A(B[4]) );
  inv02 U490 ( .Y(n453), .A(A[4]) );
  inv02 U491 ( .Y(n454), .A(carry_4_) );
  nor02 U492 ( .Y(n455), .A0(n452), .A1(n456) );
  nor02 U493 ( .Y(n457), .A0(n453), .A1(n458) );
  nor02 U494 ( .Y(n459), .A0(n454), .A1(n460) );
  nor02 U495 ( .Y(n461), .A0(n454), .A1(n462) );
  nor02 U496 ( .Y(n450), .A0(n463), .A1(n464) );
  nor02 U497 ( .Y(n465), .A0(n453), .A1(n454) );
  nor02 U498 ( .Y(n466), .A0(n452), .A1(n454) );
  nor02 U499 ( .Y(n467), .A0(n452), .A1(n453) );
  nor02 U500 ( .Y(n451), .A0(n467), .A1(n468) );
  nor02 U501 ( .Y(n469), .A0(A[4]), .A1(carry_4_) );
  inv01 U502 ( .Y(n456), .A(n469) );
  nor02 U503 ( .Y(n470), .A0(B[4]), .A1(carry_4_) );
  inv01 U504 ( .Y(n458), .A(n470) );
  nor02 U505 ( .Y(n471), .A0(B[4]), .A1(A[4]) );
  inv01 U506 ( .Y(n460), .A(n471) );
  nor02 U507 ( .Y(n472), .A0(n452), .A1(n453) );
  inv01 U508 ( .Y(n462), .A(n472) );
  nor02 U509 ( .Y(n473), .A0(n455), .A1(n457) );
  inv01 U510 ( .Y(n463), .A(n473) );
  nor02 U511 ( .Y(n474), .A0(n459), .A1(n461) );
  inv01 U512 ( .Y(n464), .A(n474) );
  nor02 U513 ( .Y(n475), .A0(n465), .A1(n466) );
  inv01 U514 ( .Y(n468), .A(n475) );
  inv02 U515 ( .Y(SUM[3]), .A(n476) );
  inv02 U516 ( .Y(carry_4_), .A(n477) );
  inv02 U517 ( .Y(n478), .A(B[3]) );
  inv02 U518 ( .Y(n479), .A(A[3]) );
  inv02 U519 ( .Y(n480), .A(carry_3_) );
  nor02 U520 ( .Y(n481), .A0(n478), .A1(n482) );
  nor02 U521 ( .Y(n483), .A0(n479), .A1(n484) );
  nor02 U522 ( .Y(n485), .A0(n480), .A1(n486) );
  nor02 U523 ( .Y(n487), .A0(n480), .A1(n488) );
  nor02 U524 ( .Y(n476), .A0(n489), .A1(n490) );
  nor02 U525 ( .Y(n491), .A0(n479), .A1(n480) );
  nor02 U526 ( .Y(n492), .A0(n478), .A1(n480) );
  nor02 U527 ( .Y(n493), .A0(n478), .A1(n479) );
  nor02 U528 ( .Y(n477), .A0(n493), .A1(n494) );
  nor02 U529 ( .Y(n495), .A0(A[3]), .A1(carry_3_) );
  inv01 U530 ( .Y(n482), .A(n495) );
  nor02 U531 ( .Y(n496), .A0(B[3]), .A1(carry_3_) );
  inv01 U532 ( .Y(n484), .A(n496) );
  nor02 U533 ( .Y(n497), .A0(B[3]), .A1(A[3]) );
  inv01 U534 ( .Y(n486), .A(n497) );
  nor02 U535 ( .Y(n498), .A0(n478), .A1(n479) );
  inv01 U536 ( .Y(n488), .A(n498) );
  nor02 U537 ( .Y(n499), .A0(n481), .A1(n483) );
  inv01 U538 ( .Y(n489), .A(n499) );
  nor02 U539 ( .Y(n500), .A0(n485), .A1(n487) );
  inv01 U540 ( .Y(n490), .A(n500) );
  nor02 U541 ( .Y(n501), .A0(n491), .A1(n492) );
  inv01 U542 ( .Y(n494), .A(n501) );
  inv02 U543 ( .Y(SUM[2]), .A(n502) );
  inv02 U544 ( .Y(carry_3_), .A(n503) );
  inv02 U545 ( .Y(n504), .A(B[2]) );
  inv02 U546 ( .Y(n505), .A(A[2]) );
  inv02 U547 ( .Y(n506), .A(carry_2_) );
  nor02 U548 ( .Y(n507), .A0(n504), .A1(n508) );
  nor02 U549 ( .Y(n509), .A0(n505), .A1(n510) );
  nor02 U550 ( .Y(n511), .A0(n506), .A1(n512) );
  nor02 U551 ( .Y(n513), .A0(n506), .A1(n514) );
  nor02 U552 ( .Y(n502), .A0(n515), .A1(n516) );
  nor02 U553 ( .Y(n517), .A0(n505), .A1(n506) );
  nor02 U554 ( .Y(n518), .A0(n504), .A1(n506) );
  nor02 U555 ( .Y(n519), .A0(n504), .A1(n505) );
  nor02 U556 ( .Y(n503), .A0(n519), .A1(n520) );
  nor02 U557 ( .Y(n521), .A0(A[2]), .A1(carry_2_) );
  inv01 U558 ( .Y(n508), .A(n521) );
  nor02 U559 ( .Y(n522), .A0(B[2]), .A1(carry_2_) );
  inv01 U560 ( .Y(n510), .A(n522) );
  nor02 U561 ( .Y(n523), .A0(B[2]), .A1(A[2]) );
  inv01 U562 ( .Y(n512), .A(n523) );
  nor02 U563 ( .Y(n524), .A0(n504), .A1(n505) );
  inv01 U564 ( .Y(n514), .A(n524) );
  nor02 U565 ( .Y(n525), .A0(n507), .A1(n509) );
  inv01 U566 ( .Y(n515), .A(n525) );
  nor02 U567 ( .Y(n526), .A0(n511), .A1(n513) );
  inv01 U568 ( .Y(n516), .A(n526) );
  nor02 U569 ( .Y(n527), .A0(n517), .A1(n518) );
  inv01 U570 ( .Y(n520), .A(n527) );
  inv02 U571 ( .Y(SUM[1]), .A(n528) );
  inv02 U572 ( .Y(carry_2_), .A(n529) );
  inv02 U573 ( .Y(n530), .A(B[1]) );
  inv02 U574 ( .Y(n531), .A(A[1]) );
  inv02 U575 ( .Y(n532), .A(n3) );
  nor02 U576 ( .Y(n533), .A0(n530), .A1(n534) );
  nor02 U577 ( .Y(n535), .A0(n531), .A1(n536) );
  nor02 U578 ( .Y(n537), .A0(n532), .A1(n538) );
  nor02 U579 ( .Y(n539), .A0(n532), .A1(n540) );
  nor02 U580 ( .Y(n528), .A0(n541), .A1(n542) );
  nor02 U581 ( .Y(n543), .A0(n531), .A1(n532) );
  nor02 U582 ( .Y(n544), .A0(n530), .A1(n532) );
  nor02 U583 ( .Y(n545), .A0(n530), .A1(n531) );
  nor02 U584 ( .Y(n529), .A0(n545), .A1(n546) );
  nor02 U585 ( .Y(n547), .A0(A[1]), .A1(n3) );
  inv01 U586 ( .Y(n534), .A(n547) );
  nor02 U587 ( .Y(n548), .A0(B[1]), .A1(n3) );
  inv01 U588 ( .Y(n536), .A(n548) );
  nor02 U589 ( .Y(n549), .A0(B[1]), .A1(A[1]) );
  inv01 U590 ( .Y(n538), .A(n549) );
  nor02 U591 ( .Y(n550), .A0(n530), .A1(n531) );
  inv01 U592 ( .Y(n540), .A(n550) );
  nor02 U593 ( .Y(n551), .A0(n533), .A1(n535) );
  inv01 U594 ( .Y(n541), .A(n551) );
  nor02 U595 ( .Y(n552), .A0(n537), .A1(n539) );
  inv01 U596 ( .Y(n542), .A(n552) );
  nor02 U597 ( .Y(n553), .A0(n543), .A1(n544) );
  inv01 U598 ( .Y(n546), .A(n553) );
  xor2 U599 ( .Y(n557), .A0(B[0]), .A1(A[0]) );
  fadd1 U1_22 ( .S(n555), .CO(carry_23_), .A(A[22]), .B(B[22]), .CI(carry_22_)
         );
  fadd1 U1_23 ( .S(n554), .A(A[23]), .B(B[23]), .CI(n4) );
endmodule


module mul_24_DW01_add_11_3 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   g_array_0__9_, g_array_0__8_, g_array_0__7_, g_array_0__6_,
         g_array_0__5_, g_array_0__4_, g_array_0__3_, g_array_0__2_,
         g_array_0__1_, g_array_0__0_, g_array_1__9_, g_array_1__8_,
         g_array_1__7_, g_array_1__6_, g_array_1__5_, g_array_1__4_,
         g_array_1__3_, g_array_1__2_, g_array_1__1_, g_array_1__0_,
         g_array_2__9_, g_array_2__8_, g_array_2__7_, g_array_2__6_,
         g_array_2__5_, g_array_2__4_, g_array_2__3_, g_array_2__2_,
         g_array_2__1_, g_array_2__0_, g_array_3__9_, g_array_3__8_,
         g_array_3__7_, g_array_3__6_, g_array_3__5_, g_array_3__4_,
         g_array_3__3_, g_array_3__2_, g_array_3__1_, g_array_3__0_,
         g_array_4__9_, g_array_4__7_, g_array_4__6_, g_array_4__5_,
         g_array_4__4_, g_array_4__3_, g_array_4__2_, g_array_4__1_,
         g_array_4__0_, pog_array_0__9_, pog_array_0__0_, pog_array_1__9_,
         pog_array_1__8_, pog_array_1__7_, pog_array_1__6_, pog_array_1__5_,
         pog_array_1__3_, pog_array_1__2_, pog_array_1__1_, pog_array_2__9_,
         pog_array_2__8_, pog_array_2__7_, pog_array_2__6_, pog_array_2__5_,
         pog_array_2__4_, pog_array_2__3_, pog_array_2__1_, pog_array_3__9_,
         pog_array_3__8_, pog_array_3__7_, pog_array_3__5_, pog_array_3__4_,
         pog_array_3__3_, part_sum_9_, part_sum_8_, part_sum_7_, part_sum_6_,
         part_sum_5_, part_sum_4_, part_sum_3_, part_sum_2_, part_sum_1_, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n93, n95, n97, n99, n101, n103, n105, n107, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140;

  inv02 U1_2_0_7 ( .Y(g_array_1__7_), .A(g_array_0__7_) );
  inv02 U1_2_0_5 ( .Y(g_array_1__5_), .A(g_array_0__5_) );
  inv01 U7 ( .Y(g_array_3__5_), .A(n31) );
  nor02 U8 ( .Y(n32), .A0(pog_array_2__5_), .A1(g_array_2__4_) );
  inv01 U9 ( .Y(n33), .A(g_array_2__5_) );
  nor02 U10 ( .Y(n31), .A0(n32), .A1(n33) );
  inv02 U1_3_1_5 ( .Y(pog_array_2__5_), .A(pog_array_1__5_) );
  inv02 U1_2_1_5 ( .Y(g_array_2__5_), .A(g_array_1__5_) );
  inv01 U11 ( .Y(g_array_3__9_), .A(n34) );
  nor02 U12 ( .Y(n35), .A0(pog_array_2__9_), .A1(g_array_2__8_) );
  inv01 U13 ( .Y(n36), .A(g_array_2__9_) );
  nor02 U14 ( .Y(n34), .A0(n35), .A1(n36) );
  inv02 U1_3_1_9 ( .Y(pog_array_2__9_), .A(pog_array_1__9_) );
  inv02 U1_2_1_9 ( .Y(g_array_2__9_), .A(g_array_1__9_) );
  inv01 U15 ( .Y(g_array_1__2_), .A(n37) );
  nor02 U16 ( .Y(n38), .A0(n115), .A1(g_array_0__1_) );
  inv01 U17 ( .Y(n39), .A(g_array_0__2_) );
  nor02 U18 ( .Y(n37), .A0(n38), .A1(n39) );
  nand02 U19 ( .Y(g_array_1__6_), .A0(n40), .A1(g_array_0__6_) );
  inv01 U20 ( .Y(n41), .A(g_array_0__5_) );
  inv01 U21 ( .Y(n42), .A(n121) );
  nand02 U22 ( .Y(n40), .A0(n41), .A1(n42) );
  nand02 U23 ( .Y(g_array_4__9_), .A0(n43), .A1(n44) );
  inv01 U24 ( .Y(n45), .A(g_array_3__9_) );
  inv01 U25 ( .Y(n46), .A(g_array_3__6_) );
  inv01 U26 ( .Y(n47), .A(pog_array_3__9_) );
  nand02 U27 ( .Y(n43), .A0(n45), .A1(n46) );
  nand02 U28 ( .Y(n44), .A0(n45), .A1(n47) );
  inv02 U1_2_0_9 ( .Y(g_array_1__9_), .A(g_array_0__9_) );
  inv02 U1_3_1_8 ( .Y(pog_array_2__8_), .A(pog_array_1__8_) );
  inv02 U1_3_2_8 ( .Y(pog_array_3__8_), .A(pog_array_2__8_) );
  inv02 U1_3_0_9 ( .Y(pog_array_1__9_), .A(pog_array_0__9_) );
  inv02 U29 ( .Y(n136), .A(pog_array_0__0_) );
  inv01 U30 ( .Y(g_array_3__1_), .A(n48) );
  nor02 U31 ( .Y(n49), .A0(pog_array_2__1_), .A1(g_array_2__0_) );
  inv01 U32 ( .Y(n50), .A(g_array_2__1_) );
  nor02 U33 ( .Y(n48), .A0(n49), .A1(n50) );
  inv01 U1_2_3_1 ( .Y(g_array_4__1_), .A(g_array_3__1_) );
  inv02 U1_3_1_1 ( .Y(pog_array_2__1_), .A(pog_array_1__1_) );
  inv02 U1_2_1_0 ( .Y(g_array_2__0_), .A(g_array_1__0_) );
  inv02 U1_2_1_1 ( .Y(g_array_2__1_), .A(g_array_1__1_) );
  nand02 U34 ( .Y(g_array_1__8_), .A0(n51), .A1(g_array_0__8_) );
  inv01 U35 ( .Y(n52), .A(g_array_0__7_) );
  inv01 U36 ( .Y(n53), .A(n119) );
  nand02 U37 ( .Y(n51), .A0(n52), .A1(n53) );
  inv02 U1_2_1_8 ( .Y(g_array_2__8_), .A(g_array_1__8_) );
  nand02 U38 ( .Y(g_array_4__7_), .A0(n54), .A1(n55) );
  inv01 U39 ( .Y(n56), .A(g_array_3__7_) );
  inv01 U40 ( .Y(n57), .A(g_array_3__6_) );
  inv01 U41 ( .Y(n58), .A(pog_array_3__7_) );
  nand02 U42 ( .Y(n54), .A0(n56), .A1(n57) );
  nand02 U43 ( .Y(n55), .A0(n56), .A1(n58) );
  ao21 U44 ( .Y(n59), .A0(pog_array_3__8_), .A1(g_array_3__6_), .B0(
        g_array_3__8_) );
  inv01 U45 ( .Y(n60), .A(n59) );
  inv02 U1_3_2_7 ( .Y(pog_array_3__7_), .A(pog_array_2__7_) );
  inv02 U1_2_2_7 ( .Y(g_array_3__7_), .A(g_array_2__7_) );
  inv02 U46 ( .Y(SUM[10]), .A(g_array_4__9_) );
  nand02 U47 ( .Y(g_array_4__3_), .A0(n61), .A1(n62) );
  inv01 U48 ( .Y(n63), .A(g_array_3__3_) );
  inv01 U49 ( .Y(n64), .A(g_array_3__2_) );
  inv01 U50 ( .Y(n65), .A(pog_array_3__3_) );
  nand02 U51 ( .Y(n61), .A0(n63), .A1(n64) );
  nand02 U52 ( .Y(n62), .A0(n63), .A1(n65) );
  nand02 U53 ( .Y(g_array_4__4_), .A0(n66), .A1(n67) );
  inv01 U54 ( .Y(n68), .A(g_array_3__4_) );
  inv01 U55 ( .Y(n69), .A(g_array_3__2_) );
  inv01 U56 ( .Y(n70), .A(pog_array_3__4_) );
  nand02 U57 ( .Y(n66), .A0(n68), .A1(n69) );
  nand02 U58 ( .Y(n67), .A0(n68), .A1(n70) );
  nand02 U59 ( .Y(g_array_4__5_), .A0(n71), .A1(n72) );
  inv01 U60 ( .Y(n73), .A(g_array_3__5_) );
  inv01 U61 ( .Y(n74), .A(g_array_3__2_) );
  inv01 U62 ( .Y(n75), .A(pog_array_3__5_) );
  nand02 U63 ( .Y(n71), .A0(n73), .A1(n74) );
  nand02 U64 ( .Y(n72), .A0(n73), .A1(n75) );
  inv02 U1_3_2_3 ( .Y(pog_array_3__3_), .A(pog_array_2__3_) );
  inv02 U1_2_2_3 ( .Y(g_array_3__3_), .A(g_array_2__3_) );
  inv02 U1_3_2_4 ( .Y(pog_array_3__4_), .A(pog_array_2__4_) );
  inv02 U1_2_2_4 ( .Y(g_array_3__4_), .A(g_array_2__4_) );
  inv02 U1_2_0_3 ( .Y(g_array_1__3_), .A(g_array_0__3_) );
  inv01 U1_2_0_1 ( .Y(g_array_1__1_), .A(g_array_0__1_) );
  nand02 U65 ( .Y(g_array_1__4_), .A0(n76), .A1(g_array_0__4_) );
  inv01 U66 ( .Y(n77), .A(g_array_0__3_) );
  inv01 U67 ( .Y(n78), .A(n117) );
  nand02 U68 ( .Y(n76), .A0(n77), .A1(n78) );
  inv02 U1_2_1_4 ( .Y(g_array_2__4_), .A(g_array_1__4_) );
  or02 U69 ( .Y(n79), .A0(A[3]), .A1(B[3]) );
  inv01 U70 ( .Y(n80), .A(n79) );
  inv02 U1_3_0_3 ( .Y(pog_array_1__3_), .A(n80) );
  or02 U71 ( .Y(n81), .A0(A[5]), .A1(B[5]) );
  inv01 U72 ( .Y(n82), .A(n81) );
  inv01 U73 ( .Y(n83), .A(n81) );
  inv02 U1_3_0_5 ( .Y(pog_array_1__5_), .A(n82) );
  or02 U74 ( .Y(n84), .A0(A[7]), .A1(B[7]) );
  inv01 U75 ( .Y(n85), .A(n84) );
  inv01 U76 ( .Y(n86), .A(n84) );
  inv02 U1_3_0_7 ( .Y(pog_array_1__7_), .A(n85) );
  or02 U77 ( .Y(n87), .A0(A[1]), .A1(B[1]) );
  inv01 U78 ( .Y(n88), .A(n87) );
  inv02 U1_3_0_1 ( .Y(pog_array_1__1_), .A(n88) );
  or02 U79 ( .Y(n89), .A0(n80), .A1(n117) );
  inv01 U80 ( .Y(n90), .A(n89) );
  inv02 U1_3_1_4 ( .Y(pog_array_2__4_), .A(n90) );
  xor2 U81 ( .Y(n91), .A0(part_sum_4_), .A1(g_array_4__3_) );
  inv02 U82 ( .Y(SUM[4]), .A(n91) );
  xor2 U83 ( .Y(n93), .A0(part_sum_8_), .A1(g_array_4__7_) );
  inv02 U84 ( .Y(SUM[8]), .A(n93) );
  xor2 U85 ( .Y(n95), .A0(part_sum_6_), .A1(g_array_4__5_) );
  inv02 U86 ( .Y(SUM[6]), .A(n95) );
  xor2 U87 ( .Y(n97), .A0(part_sum_2_), .A1(g_array_4__1_) );
  inv02 U88 ( .Y(SUM[2]), .A(n97) );
  xor2 U89 ( .Y(n99), .A0(part_sum_9_), .A1(n60) );
  inv02 U90 ( .Y(SUM[9]), .A(n99) );
  xor2 U91 ( .Y(n101), .A0(part_sum_5_), .A1(g_array_4__4_) );
  inv02 U92 ( .Y(SUM[5]), .A(n101) );
  xor2 U93 ( .Y(n103), .A0(part_sum_7_), .A1(g_array_4__6_) );
  inv02 U94 ( .Y(SUM[7]), .A(n103) );
  xor2 U95 ( .Y(n105), .A0(part_sum_3_), .A1(g_array_4__2_) );
  inv02 U96 ( .Y(SUM[3]), .A(n105) );
  xor2 U97 ( .Y(n107), .A0(part_sum_1_), .A1(g_array_4__0_) );
  inv02 U98 ( .Y(SUM[1]), .A(n107) );
  nand02 U99 ( .Y(g_array_2__2_), .A0(n109), .A1(n110) );
  inv01 U100 ( .Y(n111), .A(g_array_1__2_) );
  inv01 U101 ( .Y(n112), .A(g_array_1__0_) );
  inv01 U102 ( .Y(n113), .A(pog_array_1__2_) );
  nand02 U103 ( .Y(n109), .A0(n111), .A1(n112) );
  nand02 U104 ( .Y(n110), .A0(n111), .A1(n113) );
  inv02 U1_2_2_2 ( .Y(g_array_3__2_), .A(g_array_2__2_) );
  inv02 U105 ( .Y(g_array_1__0_), .A(g_array_0__0_) );
  or02 U106 ( .Y(n114), .A0(A[2]), .A1(B[2]) );
  inv02 U107 ( .Y(n115), .A(n114) );
  inv01 U108 ( .Y(n137), .A(n115) );
  or02 U109 ( .Y(n116), .A0(A[4]), .A1(B[4]) );
  inv02 U110 ( .Y(n117), .A(n116) );
  inv01 U111 ( .Y(n138), .A(n117) );
  or02 U112 ( .Y(n118), .A0(A[8]), .A1(B[8]) );
  inv02 U113 ( .Y(n119), .A(n118) );
  inv01 U114 ( .Y(n140), .A(n119) );
  or02 U115 ( .Y(n120), .A0(A[6]), .A1(B[6]) );
  inv01 U116 ( .Y(n121), .A(n120) );
  inv01 U117 ( .Y(n122), .A(n120) );
  inv01 U118 ( .Y(n139), .A(n121) );
  inv02 U119 ( .Y(g_array_3__6_), .A(n123) );
  nor02 U120 ( .Y(n124), .A0(pog_array_2__6_), .A1(g_array_2__2_) );
  inv01 U121 ( .Y(n125), .A(g_array_2__6_) );
  nor02 U122 ( .Y(n123), .A0(n124), .A1(n125) );
  inv01 U1_2_3_6 ( .Y(g_array_4__6_), .A(g_array_3__6_) );
  inv04 U123 ( .Y(part_sum_9_), .A(n126) );
  inv04 U124 ( .Y(part_sum_8_), .A(n127) );
  inv04 U125 ( .Y(part_sum_7_), .A(n128) );
  inv04 U126 ( .Y(part_sum_6_), .A(n129) );
  inv04 U127 ( .Y(part_sum_5_), .A(n130) );
  inv04 U128 ( .Y(part_sum_4_), .A(n131) );
  inv04 U129 ( .Y(part_sum_3_), .A(n132) );
  inv04 U130 ( .Y(part_sum_2_), .A(n133) );
  inv04 U131 ( .Y(part_sum_1_), .A(n134) );
  inv04 U132 ( .Y(SUM[0]), .A(n135) );
  nand02 U0_1_0 ( .Y(g_array_0__0_), .A0(A[0]), .A1(B[0]) );
  nor02 U0_2_0 ( .Y(pog_array_0__0_), .A0(A[0]), .A1(B[0]) );
  nand02 U0_3_0 ( .Y(n135), .A0(g_array_0__0_), .A1(n136) );
  nand02 U0_1_1 ( .Y(g_array_0__1_), .A0(A[1]), .A1(B[1]) );
  nand02 U0_3_1 ( .Y(n134), .A0(g_array_0__1_), .A1(pog_array_1__1_) );
  nand02 U0_1_2 ( .Y(g_array_0__2_), .A0(A[2]), .A1(B[2]) );
  nand02 U0_3_2 ( .Y(n133), .A0(g_array_0__2_), .A1(n137) );
  nand02 U0_1_3 ( .Y(g_array_0__3_), .A0(A[3]), .A1(B[3]) );
  nand02 U0_3_3 ( .Y(n132), .A0(g_array_0__3_), .A1(pog_array_1__3_) );
  nand02 U0_1_4 ( .Y(g_array_0__4_), .A0(A[4]), .A1(B[4]) );
  nand02 U0_3_4 ( .Y(n131), .A0(g_array_0__4_), .A1(n138) );
  nand02 U0_1_5 ( .Y(g_array_0__5_), .A0(A[5]), .A1(B[5]) );
  nand02 U0_3_5 ( .Y(n130), .A0(g_array_0__5_), .A1(pog_array_1__5_) );
  nand02 U0_1_6 ( .Y(g_array_0__6_), .A0(A[6]), .A1(B[6]) );
  nand02 U0_3_6 ( .Y(n129), .A0(g_array_0__6_), .A1(n139) );
  nand02 U0_1_7 ( .Y(g_array_0__7_), .A0(A[7]), .A1(B[7]) );
  nand02 U0_3_7 ( .Y(n128), .A0(g_array_0__7_), .A1(pog_array_1__7_) );
  nand02 U0_1_8 ( .Y(g_array_0__8_), .A0(A[8]), .A1(B[8]) );
  nand02 U0_3_8 ( .Y(n127), .A0(g_array_0__8_), .A1(n140) );
  nand02 U0_1_9 ( .Y(g_array_0__9_), .A0(A[9]), .A1(B[9]) );
  nor02 U0_2_9 ( .Y(pog_array_0__9_), .A0(A[9]), .A1(B[9]) );
  nand02 U0_3_9 ( .Y(n126), .A0(g_array_0__9_), .A1(pog_array_1__9_) );
  nor02 U1_5_0_2 ( .Y(pog_array_1__2_), .A0(n88), .A1(n115) );
  nor02 U1_5_0_6 ( .Y(pog_array_1__6_), .A0(n83), .A1(n122) );
  nor02 U1_5_0_8 ( .Y(pog_array_1__8_), .A0(n86), .A1(n119) );
  inv04 U1_2_1_3 ( .Y(g_array_2__3_), .A(g_array_1__3_) );
  inv04 U1_3_1_3 ( .Y(pog_array_2__3_), .A(pog_array_1__3_) );
  aoi21 U1_4_1_6 ( .Y(g_array_2__6_), .A0(pog_array_1__6_), .A1(g_array_1__4_), 
        .B0(g_array_1__6_) );
  nand02 U1_5_1_6 ( .Y(pog_array_2__6_), .A0(pog_array_1__6_), .A1(n90) );
  inv04 U1_2_1_7 ( .Y(g_array_2__7_), .A(g_array_1__7_) );
  inv04 U1_3_1_7 ( .Y(pog_array_2__7_), .A(pog_array_1__7_) );
  inv04 U1_2_2_0 ( .Y(g_array_3__0_), .A(g_array_2__0_) );
  nor02 U1_5_2_5 ( .Y(pog_array_3__5_), .A0(pog_array_2__4_), .A1(
        pog_array_2__5_) );
  inv04 U1_2_2_8 ( .Y(g_array_3__8_), .A(g_array_2__8_) );
  nor02 U1_5_2_9 ( .Y(pog_array_3__9_), .A0(pog_array_2__8_), .A1(
        pog_array_2__9_) );
  inv04 U1_2_3_0 ( .Y(g_array_4__0_), .A(g_array_3__0_) );
  inv04 U1_2_3_2 ( .Y(g_array_4__2_), .A(g_array_3__2_) );
endmodule


module mul_24_DW02_mult_6_6_3 ( A, B, TC, PRODUCT );
  input [5:0] A;
  input [5:0] B;
  output [11:0] PRODUCT;
  input TC;
  wire   U1_level_node_1__4__0_, U1_level_node_1__5__0_,
         U1_level_node_1__5__1_, U1_level_node_1__5__2_,
         U1_level_node_1__6__0_, U1_level_node_1__6__1_,
         U1_level_node_1__6__2_, U1_level_node_1__7__0_,
         U1_level_node_1__7__1_, U1_level_node_1__8__0_,
         U1_level_node_2__3__0_, U1_level_node_2__4__0_,
         U1_level_node_2__4__1_, U1_level_node_2__5__0_,
         U1_level_node_2__5__1_, U1_level_node_2__6__0_,
         U1_level_node_2__6__1_, U1_level_node_2__7__0_,
         U1_level_node_2__7__1_, U1_level_node_2__8__0_,
         U1_level_node_2__8__1_, U1_level_node_2__9__0_,
         U1_level_node_3__2__0_, U1_level_node_3__3__0_,
         U1_level_node_3__3__1_, U1_level_node_3__4__0_,
         U1_level_node_3__4__1_, U1_level_node_3__5__0_,
         U1_level_node_3__5__1_, U1_level_node_3__6__0_,
         U1_level_node_3__6__1_, U1_level_node_3__7__0_,
         U1_level_node_3__7__1_, U1_level_node_3__8__0_,
         U1_level_node_3__8__1_, U1_level_node_3__9__0_,
         U1_level_node_3__9__1_, U1_level_node_3__10__0_,
         U1_B_neg_correction_2_, U1_B_neg_correction_1_, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303;

  or02 U5 ( .Y(n1), .A0(n298), .A1(n301) );
  inv01 U6 ( .Y(n2), .A(n1) );
  nor02 U7 ( .Y(n3), .A0(n296), .A1(n303) );
  inv04 U8 ( .Y(n296), .A(A[2]) );
  or02 U9 ( .Y(n4), .A0(n297), .A1(n300) );
  inv01 U10 ( .Y(n5), .A(n4) );
  or02 U11 ( .Y(n6), .A0(n302), .A1(n303) );
  inv01 U12 ( .Y(n7), .A(n6) );
  or02 U13 ( .Y(n8), .A0(n299), .A1(n300) );
  inv01 U14 ( .Y(n9), .A(n8) );
  or02 U15 ( .Y(n10), .A0(n294), .A1(n301) );
  inv01 U16 ( .Y(n11), .A(n10) );
  or02 U17 ( .Y(n12), .A0(n296), .A1(n301) );
  inv01 U18 ( .Y(n13), .A(n12) );
  or02 U19 ( .Y(n14), .A0(n292), .A1(n301) );
  inv01 U20 ( .Y(n15), .A(n14) );
  or02 U21 ( .Y(n16), .A0(n298), .A1(n299) );
  inv02 U22 ( .Y(n17), .A(n16) );
  or02 U23 ( .Y(n18), .A0(n294), .A1(n299) );
  inv02 U24 ( .Y(n19), .A(n18) );
  or02 U25 ( .Y(n20), .A0(n296), .A1(n299) );
  inv02 U26 ( .Y(n21), .A(n20) );
  nand02 U27 ( .Y(n22), .A0(n47), .A1(n49) );
  inv02 U28 ( .Y(n23), .A(n22) );
  nand02 U29 ( .Y(n24), .A0(n51), .A1(n45) );
  inv02 U30 ( .Y(n25), .A(n24) );
  inv01 U31 ( .Y(n26), .A(n174) );
  inv01 U32 ( .Y(n27), .A(n122) );
  inv01 U33 ( .Y(n28), .A(n176) );
  inv01 U34 ( .Y(n29), .A(n63) );
  or02 U35 ( .Y(n30), .A0(n295), .A1(n302) );
  inv02 U36 ( .Y(n31), .A(n30) );
  or02 U37 ( .Y(n32), .A0(n295), .A1(n300) );
  inv02 U38 ( .Y(n33), .A(n32) );
  or02 U39 ( .Y(n34), .A0(n293), .A1(n300) );
  inv02 U40 ( .Y(n35), .A(n34) );
  or02 U41 ( .Y(n36), .A0(n301), .A1(n302) );
  inv02 U42 ( .Y(n37), .A(n36) );
  or02 U43 ( .Y(n38), .A0(n297), .A1(n302) );
  inv02 U44 ( .Y(n39), .A(n38) );
  or02 U45 ( .Y(n40), .A0(n293), .A1(n302) );
  inv02 U46 ( .Y(n41), .A(n40) );
  buf02 U47 ( .Y(n42), .A(U1_level_node_2__4__1_) );
  buf02 U48 ( .Y(n43), .A(U1_level_node_2__3__0_) );
  buf02 U49 ( .Y(n44), .A(U1_B_neg_correction_1_) );
  buf02 U50 ( .Y(n45), .A(U1_B_neg_correction_1_) );
  or02 U51 ( .Y(n46), .A0(n300), .A1(n303) );
  inv02 U52 ( .Y(n47), .A(n46) );
  or02 U53 ( .Y(n48), .A0(n293), .A1(n298) );
  inv02 U54 ( .Y(n49), .A(n48) );
  or02 U55 ( .Y(n50), .A0(n299), .A1(n302) );
  inv02 U56 ( .Y(n51), .A(n50) );
  or02 U57 ( .Y(n52), .A0(n292), .A1(n303) );
  inv02 U58 ( .Y(n53), .A(n52) );
  or02 U59 ( .Y(n54), .A0(n297), .A1(n298) );
  inv02 U60 ( .Y(n55), .A(n54) );
  or02 U61 ( .Y(n56), .A0(n296), .A1(n297) );
  inv02 U62 ( .Y(n57), .A(n56) );
  or02 U63 ( .Y(n58), .A0(n295), .A1(n298) );
  inv02 U64 ( .Y(n59), .A(n58) );
  inv02 U65 ( .Y(U1_level_node_2__4__0_), .A(n60) );
  inv02 U66 ( .Y(U1_level_node_2__5__1_), .A(n61) );
  inv02 U67 ( .Y(n62), .A(n57) );
  inv02 U68 ( .Y(n63), .A(U1_level_node_1__4__0_) );
  inv02 U69 ( .Y(n64), .A(n59) );
  nor02 U70 ( .Y(n65), .A0(n62), .A1(n66) );
  nor02 U71 ( .Y(n67), .A0(n63), .A1(n68) );
  nor02 U72 ( .Y(n69), .A0(n64), .A1(n70) );
  nor02 U73 ( .Y(n71), .A0(n64), .A1(n72) );
  nor02 U74 ( .Y(n60), .A0(n73), .A1(n74) );
  nor02 U75 ( .Y(n75), .A0(n63), .A1(n64) );
  nor02 U76 ( .Y(n76), .A0(n62), .A1(n64) );
  nor02 U77 ( .Y(n77), .A0(n62), .A1(n63) );
  nor02 U78 ( .Y(n61), .A0(n77), .A1(n78) );
  nor02 U79 ( .Y(n79), .A0(U1_level_node_1__4__0_), .A1(n59) );
  inv01 U80 ( .Y(n66), .A(n79) );
  nor02 U81 ( .Y(n80), .A0(n57), .A1(n59) );
  inv01 U82 ( .Y(n68), .A(n80) );
  nor02 U83 ( .Y(n81), .A0(n57), .A1(n29) );
  inv01 U84 ( .Y(n70), .A(n81) );
  nor02 U85 ( .Y(n82), .A0(n62), .A1(n63) );
  inv01 U86 ( .Y(n72), .A(n82) );
  nor02 U87 ( .Y(n83), .A0(n65), .A1(n67) );
  inv01 U88 ( .Y(n73), .A(n83) );
  nor02 U89 ( .Y(n84), .A0(n69), .A1(n71) );
  inv01 U90 ( .Y(n74), .A(n84) );
  nor02 U91 ( .Y(n85), .A0(n75), .A1(n76) );
  inv01 U92 ( .Y(n78), .A(n85) );
  or02 U93 ( .Y(n86), .A0(n292), .A1(n293) );
  inv02 U94 ( .Y(n87), .A(n86) );
  or02 U95 ( .Y(n88), .A0(n294), .A1(n303) );
  inv02 U96 ( .Y(n89), .A(n88) );
  inv02 U97 ( .Y(U1_level_node_2__8__0_), .A(n90) );
  inv02 U98 ( .Y(U1_level_node_2__9__0_), .A(n91) );
  inv02 U99 ( .Y(n92), .A(n87) );
  inv02 U100 ( .Y(n93), .A(U1_level_node_1__8__0_) );
  inv02 U101 ( .Y(n94), .A(n89) );
  nor02 U102 ( .Y(n95), .A0(n92), .A1(n96) );
  nor02 U103 ( .Y(n97), .A0(n93), .A1(n98) );
  nor02 U104 ( .Y(n99), .A0(n94), .A1(n100) );
  nor02 U105 ( .Y(n101), .A0(n94), .A1(n102) );
  nor02 U106 ( .Y(n90), .A0(n103), .A1(n104) );
  nor02 U107 ( .Y(n105), .A0(n93), .A1(n94) );
  nor02 U108 ( .Y(n106), .A0(n92), .A1(n94) );
  nor02 U109 ( .Y(n107), .A0(n92), .A1(n93) );
  nor02 U110 ( .Y(n91), .A0(n107), .A1(n108) );
  nor02 U111 ( .Y(n109), .A0(U1_level_node_1__8__0_), .A1(n89) );
  inv01 U112 ( .Y(n96), .A(n109) );
  nor02 U113 ( .Y(n110), .A0(n87), .A1(n89) );
  inv01 U114 ( .Y(n98), .A(n110) );
  nor02 U115 ( .Y(n111), .A0(n87), .A1(U1_level_node_1__8__0_) );
  inv01 U116 ( .Y(n100), .A(n111) );
  nor02 U117 ( .Y(n112), .A0(n92), .A1(n93) );
  inv01 U118 ( .Y(n102), .A(n112) );
  nor02 U119 ( .Y(n113), .A0(n95), .A1(n97) );
  inv01 U120 ( .Y(n103), .A(n113) );
  nor02 U121 ( .Y(n114), .A0(n99), .A1(n101) );
  inv01 U122 ( .Y(n104), .A(n114) );
  nor02 U123 ( .Y(n115), .A0(n105), .A1(n106) );
  inv01 U124 ( .Y(n108), .A(n115) );
  or02 U125 ( .Y(n116), .A0(n294), .A1(n297) );
  inv02 U126 ( .Y(n117), .A(n116) );
  or02 U127 ( .Y(n118), .A0(n295), .A1(n296) );
  inv02 U128 ( .Y(n119), .A(n118) );
  inv02 U129 ( .Y(U1_level_node_2__6__0_), .A(n120) );
  inv02 U130 ( .Y(U1_level_node_2__7__1_), .A(n121) );
  inv02 U131 ( .Y(n122), .A(U1_level_node_1__6__1_) );
  inv02 U132 ( .Y(n123), .A(U1_level_node_1__6__0_) );
  inv02 U133 ( .Y(n124), .A(U1_level_node_1__6__2_) );
  nor02 U134 ( .Y(n125), .A0(n122), .A1(n126) );
  nor02 U135 ( .Y(n127), .A0(n123), .A1(n128) );
  nor02 U136 ( .Y(n129), .A0(n124), .A1(n130) );
  nor02 U137 ( .Y(n131), .A0(n124), .A1(n132) );
  nor02 U138 ( .Y(n120), .A0(n133), .A1(n134) );
  nor02 U139 ( .Y(n135), .A0(n123), .A1(n124) );
  nor02 U140 ( .Y(n136), .A0(n122), .A1(n124) );
  nor02 U141 ( .Y(n137), .A0(n122), .A1(n123) );
  nor02 U142 ( .Y(n121), .A0(n137), .A1(n138) );
  nor02 U143 ( .Y(n139), .A0(U1_level_node_1__6__0_), .A1(
        U1_level_node_1__6__2_) );
  inv01 U144 ( .Y(n126), .A(n139) );
  nor02 U145 ( .Y(n140), .A0(n27), .A1(U1_level_node_1__6__2_) );
  inv01 U146 ( .Y(n128), .A(n140) );
  nor02 U147 ( .Y(n141), .A0(U1_level_node_1__6__1_), .A1(
        U1_level_node_1__6__0_) );
  inv01 U148 ( .Y(n130), .A(n141) );
  nor02 U149 ( .Y(n142), .A0(n122), .A1(n123) );
  inv01 U150 ( .Y(n132), .A(n142) );
  nor02 U151 ( .Y(n143), .A0(n125), .A1(n127) );
  inv01 U152 ( .Y(n133), .A(n143) );
  nor02 U153 ( .Y(n144), .A0(n129), .A1(n131) );
  inv01 U154 ( .Y(n134), .A(n144) );
  nor02 U155 ( .Y(n145), .A0(n135), .A1(n136) );
  inv01 U156 ( .Y(n138), .A(n145) );
  inv02 U157 ( .Y(U1_level_node_1__5__0_), .A(n146) );
  inv02 U158 ( .Y(U1_level_node_1__6__2_), .A(n147) );
  inv02 U159 ( .Y(n148), .A(n117) );
  inv02 U160 ( .Y(n149), .A(n288) );
  inv02 U161 ( .Y(n150), .A(n119) );
  nor02 U162 ( .Y(n151), .A0(n148), .A1(n152) );
  nor02 U163 ( .Y(n153), .A0(n149), .A1(n154) );
  nor02 U164 ( .Y(n155), .A0(n150), .A1(n156) );
  nor02 U165 ( .Y(n157), .A0(n150), .A1(n158) );
  nor02 U166 ( .Y(n146), .A0(n159), .A1(n160) );
  nor02 U167 ( .Y(n161), .A0(n149), .A1(n150) );
  nor02 U168 ( .Y(n162), .A0(n148), .A1(n150) );
  nor02 U169 ( .Y(n163), .A0(n148), .A1(n149) );
  nor02 U170 ( .Y(n147), .A0(n163), .A1(n164) );
  nor02 U171 ( .Y(n165), .A0(n288), .A1(n119) );
  inv01 U172 ( .Y(n152), .A(n165) );
  nor02 U173 ( .Y(n166), .A0(n117), .A1(n119) );
  inv01 U174 ( .Y(n154), .A(n166) );
  nor02 U175 ( .Y(n167), .A0(n117), .A1(n288) );
  inv01 U176 ( .Y(n156), .A(n167) );
  nor02 U177 ( .Y(n168), .A0(n148), .A1(n149) );
  inv01 U178 ( .Y(n158), .A(n168) );
  nor02 U179 ( .Y(n169), .A0(n151), .A1(n153) );
  inv01 U180 ( .Y(n159), .A(n169) );
  nor02 U181 ( .Y(n170), .A0(n155), .A1(n157) );
  inv01 U182 ( .Y(n160), .A(n170) );
  nor02 U183 ( .Y(n171), .A0(n161), .A1(n162) );
  inv01 U184 ( .Y(n164), .A(n171) );
  inv02 U185 ( .Y(U1_level_node_2__5__0_), .A(n172) );
  inv02 U186 ( .Y(U1_level_node_2__6__1_), .A(n173) );
  inv02 U187 ( .Y(n174), .A(U1_level_node_1__5__1_) );
  inv02 U188 ( .Y(n175), .A(U1_level_node_1__5__0_) );
  inv02 U189 ( .Y(n176), .A(U1_level_node_1__5__2_) );
  nor02 U190 ( .Y(n177), .A0(n174), .A1(n178) );
  nor02 U191 ( .Y(n179), .A0(n175), .A1(n180) );
  nor02 U192 ( .Y(n181), .A0(n176), .A1(n182) );
  nor02 U193 ( .Y(n183), .A0(n176), .A1(n184) );
  nor02 U194 ( .Y(n172), .A0(n185), .A1(n186) );
  nor02 U195 ( .Y(n187), .A0(n175), .A1(n176) );
  nor02 U196 ( .Y(n188), .A0(n174), .A1(n176) );
  nor02 U197 ( .Y(n189), .A0(n174), .A1(n175) );
  nor02 U198 ( .Y(n173), .A0(n189), .A1(n190) );
  nor02 U199 ( .Y(n191), .A0(U1_level_node_1__5__0_), .A1(
        U1_level_node_1__5__2_) );
  inv01 U200 ( .Y(n178), .A(n191) );
  nor02 U201 ( .Y(n192), .A0(n26), .A1(n28) );
  inv01 U202 ( .Y(n180), .A(n192) );
  nor02 U203 ( .Y(n193), .A0(U1_level_node_1__5__1_), .A1(
        U1_level_node_1__5__0_) );
  inv01 U204 ( .Y(n182), .A(n193) );
  nor02 U205 ( .Y(n194), .A0(n174), .A1(n175) );
  inv01 U206 ( .Y(n184), .A(n194) );
  nor02 U207 ( .Y(n195), .A0(n177), .A1(n179) );
  inv01 U208 ( .Y(n185), .A(n195) );
  nor02 U209 ( .Y(n196), .A0(n181), .A1(n183) );
  inv01 U210 ( .Y(n186), .A(n196) );
  nor02 U211 ( .Y(n197), .A0(n187), .A1(n188) );
  inv01 U212 ( .Y(n190), .A(n197) );
  nor02 U213 ( .Y(n198), .A0(n296), .A1(n303) );
  or02 U214 ( .Y(n199), .A0(n293), .A1(n296) );
  inv02 U215 ( .Y(n200), .A(n199) );
  or02 U216 ( .Y(n201), .A0(n293), .A1(n294) );
  inv02 U217 ( .Y(n202), .A(n201) );
  or02 U218 ( .Y(n203), .A0(n294), .A1(n295) );
  inv02 U219 ( .Y(n204), .A(n203) );
  inv04 U220 ( .Y(n303), .A(B[5]) );
  inv02 U221 ( .Y(U1_level_node_1__7__0_), .A(n205) );
  inv02 U222 ( .Y(U1_level_node_1__8__0_), .A(n206) );
  inv02 U223 ( .Y(n207), .A(n202) );
  inv02 U224 ( .Y(n208), .A(n284) );
  inv02 U225 ( .Y(n209), .A(U1_B_neg_correction_2_) );
  nor02 U226 ( .Y(n210), .A0(n207), .A1(n211) );
  nor02 U227 ( .Y(n212), .A0(n208), .A1(n213) );
  nor02 U228 ( .Y(n214), .A0(n209), .A1(n215) );
  nor02 U229 ( .Y(n216), .A0(n209), .A1(n217) );
  nor02 U230 ( .Y(n205), .A0(n218), .A1(n219) );
  nor02 U231 ( .Y(n220), .A0(n208), .A1(n209) );
  nor02 U232 ( .Y(n221), .A0(n207), .A1(n209) );
  nor02 U233 ( .Y(n222), .A0(n207), .A1(n208) );
  nor02 U234 ( .Y(n206), .A0(n222), .A1(n223) );
  nor02 U235 ( .Y(n224), .A0(n284), .A1(n198) );
  inv01 U236 ( .Y(n211), .A(n224) );
  nor02 U237 ( .Y(n225), .A0(n202), .A1(n3) );
  inv01 U238 ( .Y(n213), .A(n225) );
  nor02 U239 ( .Y(n226), .A0(n202), .A1(n284) );
  inv01 U240 ( .Y(n215), .A(n226) );
  nor02 U241 ( .Y(n227), .A0(n207), .A1(n208) );
  inv01 U242 ( .Y(n217), .A(n227) );
  nor02 U243 ( .Y(n228), .A0(n210), .A1(n212) );
  inv01 U244 ( .Y(n218), .A(n228) );
  nor02 U245 ( .Y(n229), .A0(n214), .A1(n216) );
  inv01 U246 ( .Y(n219), .A(n229) );
  nor02 U247 ( .Y(n230), .A0(n220), .A1(n221) );
  inv01 U248 ( .Y(n223), .A(n230) );
  inv02 U249 ( .Y(U1_level_node_1__6__0_), .A(n231) );
  inv02 U250 ( .Y(U1_level_node_1__7__1_), .A(n232) );
  inv02 U251 ( .Y(n233), .A(n204) );
  inv02 U252 ( .Y(n234), .A(n286) );
  inv02 U253 ( .Y(n235), .A(n200) );
  nor02 U254 ( .Y(n236), .A0(n233), .A1(n237) );
  nor02 U255 ( .Y(n238), .A0(n234), .A1(n239) );
  nor02 U256 ( .Y(n240), .A0(n235), .A1(n241) );
  nor02 U257 ( .Y(n242), .A0(n235), .A1(n243) );
  nor02 U258 ( .Y(n231), .A0(n244), .A1(n245) );
  nor02 U259 ( .Y(n246), .A0(n234), .A1(n235) );
  nor02 U260 ( .Y(n247), .A0(n233), .A1(n235) );
  nor02 U261 ( .Y(n248), .A0(n233), .A1(n234) );
  nor02 U262 ( .Y(n232), .A0(n248), .A1(n249) );
  nor02 U263 ( .Y(n250), .A0(n286), .A1(n200) );
  inv01 U264 ( .Y(n237), .A(n250) );
  nor02 U265 ( .Y(n251), .A0(n204), .A1(n200) );
  inv01 U266 ( .Y(n239), .A(n251) );
  nor02 U267 ( .Y(n252), .A0(n204), .A1(n286) );
  inv01 U268 ( .Y(n241), .A(n252) );
  nor02 U269 ( .Y(n253), .A0(n233), .A1(n234) );
  inv01 U270 ( .Y(n243), .A(n253) );
  nor02 U271 ( .Y(n254), .A0(n236), .A1(n238) );
  inv01 U272 ( .Y(n244), .A(n254) );
  nor02 U273 ( .Y(n255), .A0(n240), .A1(n242) );
  inv01 U274 ( .Y(n245), .A(n255) );
  nor02 U275 ( .Y(n256), .A0(n246), .A1(n247) );
  inv01 U276 ( .Y(n249), .A(n256) );
  inv02 U277 ( .Y(U1_level_node_2__7__0_), .A(n257) );
  inv02 U278 ( .Y(U1_level_node_2__8__1_), .A(n258) );
  inv02 U279 ( .Y(n259), .A(U1_level_node_1__7__1_) );
  inv02 U280 ( .Y(n260), .A(U1_level_node_1__7__0_) );
  inv02 U281 ( .Y(n261), .A(n25) );
  nor02 U282 ( .Y(n262), .A0(n259), .A1(n263) );
  nor02 U283 ( .Y(n264), .A0(n260), .A1(n265) );
  nor02 U284 ( .Y(n266), .A0(n261), .A1(n267) );
  nor02 U285 ( .Y(n268), .A0(n261), .A1(n269) );
  nor02 U286 ( .Y(n257), .A0(n270), .A1(n271) );
  nor02 U287 ( .Y(n272), .A0(n260), .A1(n261) );
  nor02 U288 ( .Y(n273), .A0(n259), .A1(n261) );
  nor02 U289 ( .Y(n274), .A0(n259), .A1(n260) );
  nor02 U290 ( .Y(n258), .A0(n274), .A1(n275) );
  nor02 U291 ( .Y(n276), .A0(U1_level_node_1__7__0_), .A1(n25) );
  inv01 U292 ( .Y(n263), .A(n276) );
  nor02 U293 ( .Y(n277), .A0(U1_level_node_1__7__1_), .A1(n25) );
  inv01 U294 ( .Y(n265), .A(n277) );
  nor02 U295 ( .Y(n278), .A0(U1_level_node_1__7__1_), .A1(
        U1_level_node_1__7__0_) );
  inv01 U296 ( .Y(n267), .A(n278) );
  nor02 U297 ( .Y(n279), .A0(n259), .A1(n260) );
  inv01 U298 ( .Y(n269), .A(n279) );
  nor02 U299 ( .Y(n280), .A0(n262), .A1(n264) );
  inv01 U300 ( .Y(n270), .A(n280) );
  nor02 U301 ( .Y(n281), .A0(n266), .A1(n268) );
  inv01 U302 ( .Y(n271), .A(n281) );
  nor02 U303 ( .Y(n282), .A0(n272), .A1(n273) );
  inv01 U304 ( .Y(n275), .A(n282) );
  or02 U305 ( .Y(n283), .A0(n292), .A1(n295) );
  inv02 U306 ( .Y(n284), .A(n283) );
  or02 U307 ( .Y(n285), .A0(n292), .A1(n297) );
  inv02 U308 ( .Y(n286), .A(n285) );
  or02 U309 ( .Y(n287), .A0(n292), .A1(n299) );
  inv02 U310 ( .Y(n288), .A(n287) );
  or02 U311 ( .Y(n289), .A0(n300), .A1(n301) );
  inv02 U312 ( .Y(PRODUCT[0]), .A(n289) );
  inv02 U313 ( .Y(n292), .A(A[4]) );
  inv02 U314 ( .Y(n298), .A(A[1]) );
  inv02 U315 ( .Y(n293), .A(B[4]) );
  inv02 U316 ( .Y(n299), .A(B[1]) );
  inv02 U317 ( .Y(n302), .A(A[5]) );
  inv02 U318 ( .Y(n297), .A(B[2]) );
  inv02 U319 ( .Y(n301), .A(B[0]) );
  inv02 U320 ( .Y(n295), .A(B[3]) );
  inv02 U321 ( .Y(n300), .A(A[0]) );
  inv02 U322 ( .Y(n294), .A(A[3]) );
  xor2 U323 ( .Y(U1_level_node_1__5__1_), .A0(n49), .A1(n47) );
  xor2 U324 ( .Y(U1_level_node_1__6__1_), .A0(n44), .A1(n51) );
  mul_24_DW01_add_11_3 U1_U9720 ( .A({1'b0, U1_level_node_3__10__0_, 
        U1_level_node_3__9__0_, U1_level_node_3__8__0_, U1_level_node_3__7__0_, 
        U1_level_node_3__6__0_, U1_level_node_3__5__0_, U1_level_node_3__4__0_, 
        U1_level_node_3__3__0_, U1_level_node_3__2__0_, n2}), .B({1'b0, n7, 
        U1_level_node_3__9__1_, U1_level_node_3__8__1_, U1_level_node_3__7__1_, 
        U1_level_node_3__6__1_, U1_level_node_3__5__1_, U1_level_node_3__4__1_, 
        U1_level_node_3__3__1_, n5, n9}), .CI(1'b0), .SUM(PRODUCT[11:1]) );
  nor02 U325 ( .Y(U1_B_neg_correction_2_), .A0(n296), .A1(n303) );
  nor02 U326 ( .Y(U1_B_neg_correction_1_), .A0(n298), .A1(n303) );
  hadd1 U1_U3220_1_4 ( .S(U1_level_node_1__4__0_), .CO(U1_level_node_1__5__2_), 
        .A(n15), .B(n19) );
  hadd1 U1_U3220_2_3 ( .S(U1_level_node_2__3__0_), .CO(U1_level_node_2__4__1_), 
        .A(n11), .B(n21) );
  fadd1 U1_U3140_3_9_0 ( .S(U1_level_node_3__9__0_), .CO(
        U1_level_node_3__10__0_), .A(U1_level_node_2__9__0_), .B(n53), .CI(n41) );
  fadd1 U1_U3140_3_8_0 ( .S(U1_level_node_3__8__0_), .CO(
        U1_level_node_3__9__1_), .A(U1_level_node_2__8__0_), .B(
        U1_level_node_2__8__1_), .CI(n31) );
  fadd1 U1_U3140_3_7_0 ( .S(U1_level_node_3__7__0_), .CO(
        U1_level_node_3__8__1_), .A(U1_level_node_2__7__0_), .B(
        U1_level_node_2__7__1_), .CI(n39) );
  fadd1 U1_U3140_3_6_0 ( .S(U1_level_node_3__6__0_), .CO(
        U1_level_node_3__7__1_), .A(U1_level_node_2__6__0_), .B(
        U1_level_node_2__6__1_), .CI(n23) );
  fadd1 U1_U3140_3_5_0 ( .S(U1_level_node_3__5__0_), .CO(
        U1_level_node_3__6__1_), .A(U1_level_node_2__5__0_), .B(
        U1_level_node_2__5__1_), .CI(n37) );
  fadd1 U1_U3140_3_4_0 ( .S(U1_level_node_3__4__0_), .CO(
        U1_level_node_3__5__1_), .A(U1_level_node_2__4__0_), .B(n42), .CI(n35)
         );
  fadd1 U1_U3140_3_3_0 ( .S(U1_level_node_3__3__0_), .CO(
        U1_level_node_3__4__1_), .A(n43), .B(n55), .CI(n33) );
  hadd1 U1_U3220_3_2 ( .S(U1_level_node_3__2__0_), .CO(U1_level_node_3__3__1_), 
        .A(n13), .B(n17) );
endmodule


module mul_24_DW01_add_11_2 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   g_array_0__9_, g_array_0__8_, g_array_0__7_, g_array_0__6_,
         g_array_0__5_, g_array_0__4_, g_array_0__3_, g_array_0__2_,
         g_array_0__1_, g_array_0__0_, g_array_1__9_, g_array_1__8_,
         g_array_1__7_, g_array_1__6_, g_array_1__5_, g_array_1__4_,
         g_array_1__3_, g_array_1__2_, g_array_1__1_, g_array_1__0_,
         g_array_2__9_, g_array_2__8_, g_array_2__7_, g_array_2__6_,
         g_array_2__5_, g_array_2__4_, g_array_2__3_, g_array_2__2_,
         g_array_2__1_, g_array_2__0_, g_array_3__9_, g_array_3__8_,
         g_array_3__7_, g_array_3__6_, g_array_3__5_, g_array_3__4_,
         g_array_3__3_, g_array_3__2_, g_array_3__1_, g_array_3__0_,
         g_array_4__9_, g_array_4__6_, g_array_4__5_, g_array_4__3_,
         g_array_4__2_, g_array_4__1_, g_array_4__0_, pog_array_0__9_,
         pog_array_0__0_, pog_array_1__9_, pog_array_1__8_, pog_array_1__7_,
         pog_array_1__6_, pog_array_1__5_, pog_array_1__3_, pog_array_1__2_,
         pog_array_1__1_, pog_array_2__9_, pog_array_2__8_, pog_array_2__7_,
         pog_array_2__6_, pog_array_2__5_, pog_array_2__4_, pog_array_2__3_,
         pog_array_2__1_, pog_array_3__9_, pog_array_3__8_, pog_array_3__7_,
         pog_array_3__5_, pog_array_3__4_, pog_array_3__3_, part_sum_9_,
         part_sum_8_, part_sum_7_, part_sum_6_, part_sum_5_, part_sum_4_,
         part_sum_3_, part_sum_2_, part_sum_1_, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n87, n89, n91, n93, n95, n97, n99,
         n101, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134;

  inv02 U1_2_0_7 ( .Y(g_array_1__7_), .A(g_array_0__7_) );
  inv02 U1_2_0_5 ( .Y(g_array_1__5_), .A(g_array_0__5_) );
  inv02 U1_2_0_3 ( .Y(g_array_1__3_), .A(g_array_0__3_) );
  inv02 U7 ( .Y(part_sum_3_), .A(n126) );
  inv02 U8 ( .Y(part_sum_7_), .A(n122) );
  inv02 U9 ( .Y(part_sum_5_), .A(n124) );
  inv01 U10 ( .Y(g_array_3__5_), .A(n31) );
  nor02 U11 ( .Y(n32), .A0(pog_array_2__5_), .A1(g_array_2__4_) );
  inv01 U12 ( .Y(n33), .A(g_array_2__5_) );
  nor02 U13 ( .Y(n31), .A0(n32), .A1(n33) );
  inv02 U1_3_1_5 ( .Y(pog_array_2__5_), .A(pog_array_1__5_) );
  inv02 U1_2_1_5 ( .Y(g_array_2__5_), .A(g_array_1__5_) );
  inv01 U14 ( .Y(g_array_3__9_), .A(n34) );
  nor02 U15 ( .Y(n35), .A0(pog_array_2__9_), .A1(g_array_2__8_) );
  inv01 U16 ( .Y(n36), .A(g_array_2__9_) );
  nor02 U17 ( .Y(n34), .A0(n35), .A1(n36) );
  inv02 U1_3_1_9 ( .Y(pog_array_2__9_), .A(pog_array_1__9_) );
  inv02 U1_2_1_9 ( .Y(g_array_2__9_), .A(g_array_1__9_) );
  inv01 U18 ( .Y(g_array_1__2_), .A(n37) );
  nor02 U19 ( .Y(n38), .A0(n109), .A1(g_array_0__1_) );
  inv01 U20 ( .Y(n39), .A(g_array_0__2_) );
  nor02 U21 ( .Y(n37), .A0(n38), .A1(n39) );
  nand02 U22 ( .Y(g_array_1__6_), .A0(n40), .A1(g_array_0__6_) );
  inv01 U23 ( .Y(n41), .A(g_array_0__5_) );
  inv01 U24 ( .Y(n42), .A(n115) );
  nand02 U25 ( .Y(n40), .A0(n41), .A1(n42) );
  nand02 U26 ( .Y(g_array_4__9_), .A0(n43), .A1(n44) );
  inv01 U27 ( .Y(n45), .A(g_array_3__9_) );
  inv01 U28 ( .Y(n46), .A(g_array_3__6_) );
  inv01 U29 ( .Y(n47), .A(pog_array_3__9_) );
  nand02 U30 ( .Y(n43), .A0(n45), .A1(n46) );
  nand02 U31 ( .Y(n44), .A0(n45), .A1(n47) );
  inv02 U1_2_0_9 ( .Y(g_array_1__9_), .A(g_array_0__9_) );
  inv02 U1_3_1_8 ( .Y(pog_array_2__8_), .A(pog_array_1__8_) );
  inv02 U1_3_2_8 ( .Y(pog_array_3__8_), .A(pog_array_2__8_) );
  inv02 U1_3_0_9 ( .Y(pog_array_1__9_), .A(pog_array_0__9_) );
  inv02 U32 ( .Y(n130), .A(pog_array_0__0_) );
  inv01 U33 ( .Y(g_array_3__1_), .A(n48) );
  nor02 U34 ( .Y(n49), .A0(pog_array_2__1_), .A1(g_array_2__0_) );
  inv01 U35 ( .Y(n50), .A(g_array_2__1_) );
  nor02 U36 ( .Y(n48), .A0(n49), .A1(n50) );
  inv01 U1_2_3_1 ( .Y(g_array_4__1_), .A(g_array_3__1_) );
  inv02 U1_3_1_1 ( .Y(pog_array_2__1_), .A(pog_array_1__1_) );
  inv02 U1_2_1_0 ( .Y(g_array_2__0_), .A(g_array_1__0_) );
  inv02 U1_2_1_1 ( .Y(g_array_2__1_), .A(g_array_1__1_) );
  nand02 U37 ( .Y(g_array_1__8_), .A0(n51), .A1(g_array_0__8_) );
  inv01 U38 ( .Y(n52), .A(g_array_0__7_) );
  inv01 U39 ( .Y(n53), .A(n113) );
  nand02 U40 ( .Y(n51), .A0(n52), .A1(n53) );
  inv02 U1_2_1_8 ( .Y(g_array_2__8_), .A(g_array_1__8_) );
  ao21 U41 ( .Y(n54), .A0(pog_array_3__8_), .A1(g_array_3__6_), .B0(
        g_array_3__8_) );
  inv01 U42 ( .Y(n55), .A(n54) );
  ao21 U43 ( .Y(n56), .A0(pog_array_3__7_), .A1(g_array_3__6_), .B0(
        g_array_3__7_) );
  inv01 U44 ( .Y(n57), .A(n56) );
  inv02 U45 ( .Y(SUM[10]), .A(g_array_4__9_) );
  ao21 U46 ( .Y(n58), .A0(pog_array_3__4_), .A1(g_array_3__2_), .B0(
        g_array_3__4_) );
  inv01 U47 ( .Y(n59), .A(n58) );
  nand02 U48 ( .Y(g_array_4__3_), .A0(n60), .A1(n61) );
  inv01 U49 ( .Y(n62), .A(g_array_3__3_) );
  inv01 U50 ( .Y(n63), .A(g_array_3__2_) );
  inv01 U51 ( .Y(n64), .A(pog_array_3__3_) );
  nand02 U52 ( .Y(n60), .A0(n62), .A1(n63) );
  nand02 U53 ( .Y(n61), .A0(n62), .A1(n64) );
  nand02 U54 ( .Y(g_array_4__5_), .A0(n65), .A1(n66) );
  inv01 U55 ( .Y(n67), .A(g_array_3__5_) );
  inv01 U56 ( .Y(n68), .A(g_array_3__2_) );
  inv01 U57 ( .Y(n69), .A(pog_array_3__5_) );
  nand02 U58 ( .Y(n65), .A0(n67), .A1(n68) );
  nand02 U59 ( .Y(n66), .A0(n67), .A1(n69) );
  inv02 U1_3_2_3 ( .Y(pog_array_3__3_), .A(pog_array_2__3_) );
  inv02 U1_2_2_3 ( .Y(g_array_3__3_), .A(g_array_2__3_) );
  inv01 U1_2_0_1 ( .Y(g_array_1__1_), .A(g_array_0__1_) );
  nand02 U60 ( .Y(g_array_1__4_), .A0(n70), .A1(g_array_0__4_) );
  inv01 U61 ( .Y(n71), .A(g_array_0__3_) );
  inv01 U62 ( .Y(n72), .A(n111) );
  nand02 U63 ( .Y(n70), .A0(n71), .A1(n72) );
  inv02 U1_2_1_4 ( .Y(g_array_2__4_), .A(g_array_1__4_) );
  or02 U64 ( .Y(n73), .A0(A[3]), .A1(B[3]) );
  inv01 U65 ( .Y(n74), .A(n73) );
  inv02 U1_3_0_3 ( .Y(pog_array_1__3_), .A(n74) );
  or02 U66 ( .Y(n75), .A0(A[5]), .A1(B[5]) );
  inv01 U67 ( .Y(n76), .A(n75) );
  inv01 U68 ( .Y(n77), .A(n75) );
  inv02 U1_3_0_5 ( .Y(pog_array_1__5_), .A(n76) );
  or02 U69 ( .Y(n78), .A0(A[7]), .A1(B[7]) );
  inv01 U70 ( .Y(n79), .A(n78) );
  inv01 U71 ( .Y(n80), .A(n78) );
  inv02 U1_3_0_7 ( .Y(pog_array_1__7_), .A(n79) );
  or02 U72 ( .Y(n81), .A0(A[1]), .A1(B[1]) );
  inv01 U73 ( .Y(n82), .A(n81) );
  inv02 U1_3_0_1 ( .Y(pog_array_1__1_), .A(n82) );
  or02 U74 ( .Y(n83), .A0(n74), .A1(n111) );
  inv01 U75 ( .Y(n84), .A(n83) );
  inv02 U1_3_1_4 ( .Y(pog_array_2__4_), .A(n84) );
  xor2 U76 ( .Y(n85), .A0(part_sum_8_), .A1(n57) );
  inv02 U77 ( .Y(SUM[8]), .A(n85) );
  xor2 U78 ( .Y(n87), .A0(part_sum_4_), .A1(g_array_4__3_) );
  inv02 U79 ( .Y(SUM[4]), .A(n87) );
  xor2 U80 ( .Y(n89), .A0(part_sum_2_), .A1(g_array_4__1_) );
  inv02 U81 ( .Y(SUM[2]), .A(n89) );
  xor2 U82 ( .Y(n91), .A0(part_sum_6_), .A1(g_array_4__5_) );
  inv02 U83 ( .Y(SUM[6]), .A(n91) );
  xor2 U84 ( .Y(n93), .A0(part_sum_9_), .A1(n55) );
  inv02 U85 ( .Y(SUM[9]), .A(n93) );
  xor2 U86 ( .Y(n95), .A0(part_sum_5_), .A1(n59) );
  inv02 U87 ( .Y(SUM[5]), .A(n95) );
  xor2 U88 ( .Y(n97), .A0(part_sum_3_), .A1(g_array_4__2_) );
  inv02 U89 ( .Y(SUM[3]), .A(n97) );
  xor2 U90 ( .Y(n99), .A0(part_sum_7_), .A1(g_array_4__6_) );
  inv02 U91 ( .Y(SUM[7]), .A(n99) );
  xor2 U92 ( .Y(n101), .A0(part_sum_1_), .A1(g_array_4__0_) );
  inv02 U93 ( .Y(SUM[1]), .A(n101) );
  nand02 U94 ( .Y(g_array_2__2_), .A0(n103), .A1(n104) );
  inv01 U95 ( .Y(n105), .A(g_array_1__2_) );
  inv01 U96 ( .Y(n106), .A(g_array_1__0_) );
  inv01 U97 ( .Y(n107), .A(pog_array_1__2_) );
  nand02 U98 ( .Y(n103), .A0(n105), .A1(n106) );
  nand02 U99 ( .Y(n104), .A0(n105), .A1(n107) );
  inv02 U1_2_2_2 ( .Y(g_array_3__2_), .A(g_array_2__2_) );
  inv02 U100 ( .Y(g_array_1__0_), .A(g_array_0__0_) );
  or02 U101 ( .Y(n108), .A0(A[2]), .A1(B[2]) );
  inv02 U102 ( .Y(n109), .A(n108) );
  inv01 U103 ( .Y(n131), .A(n109) );
  or02 U104 ( .Y(n110), .A0(A[4]), .A1(B[4]) );
  inv02 U105 ( .Y(n111), .A(n110) );
  inv01 U106 ( .Y(n132), .A(n111) );
  or02 U107 ( .Y(n112), .A0(A[8]), .A1(B[8]) );
  inv02 U108 ( .Y(n113), .A(n112) );
  inv01 U109 ( .Y(n134), .A(n113) );
  or02 U110 ( .Y(n114), .A0(A[6]), .A1(B[6]) );
  inv01 U111 ( .Y(n115), .A(n114) );
  inv01 U112 ( .Y(n116), .A(n114) );
  inv01 U113 ( .Y(n133), .A(n115) );
  inv02 U114 ( .Y(g_array_3__6_), .A(n117) );
  nor02 U115 ( .Y(n118), .A0(pog_array_2__6_), .A1(g_array_2__2_) );
  inv01 U116 ( .Y(n119), .A(g_array_2__6_) );
  nor02 U117 ( .Y(n117), .A0(n118), .A1(n119) );
  inv01 U1_2_3_6 ( .Y(g_array_4__6_), .A(g_array_3__6_) );
  inv04 U118 ( .Y(part_sum_9_), .A(n120) );
  inv04 U119 ( .Y(part_sum_8_), .A(n121) );
  inv04 U120 ( .Y(part_sum_6_), .A(n123) );
  inv04 U121 ( .Y(part_sum_4_), .A(n125) );
  inv04 U122 ( .Y(part_sum_2_), .A(n127) );
  inv04 U123 ( .Y(part_sum_1_), .A(n128) );
  inv04 U124 ( .Y(SUM[0]), .A(n129) );
  nand02 U0_1_0 ( .Y(g_array_0__0_), .A0(A[0]), .A1(B[0]) );
  nor02 U0_2_0 ( .Y(pog_array_0__0_), .A0(A[0]), .A1(B[0]) );
  nand02 U0_3_0 ( .Y(n129), .A0(g_array_0__0_), .A1(n130) );
  nand02 U0_1_1 ( .Y(g_array_0__1_), .A0(A[1]), .A1(B[1]) );
  nand02 U0_3_1 ( .Y(n128), .A0(g_array_0__1_), .A1(pog_array_1__1_) );
  nand02 U0_1_2 ( .Y(g_array_0__2_), .A0(A[2]), .A1(B[2]) );
  nand02 U0_3_2 ( .Y(n127), .A0(g_array_0__2_), .A1(n131) );
  nand02 U0_1_3 ( .Y(g_array_0__3_), .A0(A[3]), .A1(B[3]) );
  nand02 U0_3_3 ( .Y(n126), .A0(g_array_0__3_), .A1(pog_array_1__3_) );
  nand02 U0_1_4 ( .Y(g_array_0__4_), .A0(A[4]), .A1(B[4]) );
  nand02 U0_3_4 ( .Y(n125), .A0(g_array_0__4_), .A1(n132) );
  nand02 U0_1_5 ( .Y(g_array_0__5_), .A0(A[5]), .A1(B[5]) );
  nand02 U0_3_5 ( .Y(n124), .A0(g_array_0__5_), .A1(pog_array_1__5_) );
  nand02 U0_1_6 ( .Y(g_array_0__6_), .A0(A[6]), .A1(B[6]) );
  nand02 U0_3_6 ( .Y(n123), .A0(g_array_0__6_), .A1(n133) );
  nand02 U0_1_7 ( .Y(g_array_0__7_), .A0(A[7]), .A1(B[7]) );
  nand02 U0_3_7 ( .Y(n122), .A0(g_array_0__7_), .A1(pog_array_1__7_) );
  nand02 U0_1_8 ( .Y(g_array_0__8_), .A0(A[8]), .A1(B[8]) );
  nand02 U0_3_8 ( .Y(n121), .A0(g_array_0__8_), .A1(n134) );
  nand02 U0_1_9 ( .Y(g_array_0__9_), .A0(A[9]), .A1(B[9]) );
  nor02 U0_2_9 ( .Y(pog_array_0__9_), .A0(A[9]), .A1(B[9]) );
  nand02 U0_3_9 ( .Y(n120), .A0(g_array_0__9_), .A1(pog_array_1__9_) );
  nor02 U1_5_0_2 ( .Y(pog_array_1__2_), .A0(n82), .A1(n109) );
  nor02 U1_5_0_6 ( .Y(pog_array_1__6_), .A0(n77), .A1(n116) );
  nor02 U1_5_0_8 ( .Y(pog_array_1__8_), .A0(n80), .A1(n113) );
  inv04 U1_2_1_3 ( .Y(g_array_2__3_), .A(g_array_1__3_) );
  inv04 U1_3_1_3 ( .Y(pog_array_2__3_), .A(pog_array_1__3_) );
  aoi21 U1_4_1_6 ( .Y(g_array_2__6_), .A0(pog_array_1__6_), .A1(g_array_1__4_), 
        .B0(g_array_1__6_) );
  nand02 U1_5_1_6 ( .Y(pog_array_2__6_), .A0(pog_array_1__6_), .A1(n84) );
  inv04 U1_2_1_7 ( .Y(g_array_2__7_), .A(g_array_1__7_) );
  inv04 U1_3_1_7 ( .Y(pog_array_2__7_), .A(pog_array_1__7_) );
  inv04 U1_2_2_0 ( .Y(g_array_3__0_), .A(g_array_2__0_) );
  inv04 U1_2_2_4 ( .Y(g_array_3__4_), .A(g_array_2__4_) );
  inv04 U1_3_2_4 ( .Y(pog_array_3__4_), .A(pog_array_2__4_) );
  nor02 U1_5_2_5 ( .Y(pog_array_3__5_), .A0(pog_array_2__4_), .A1(
        pog_array_2__5_) );
  inv04 U1_2_2_7 ( .Y(g_array_3__7_), .A(g_array_2__7_) );
  inv04 U1_3_2_7 ( .Y(pog_array_3__7_), .A(pog_array_2__7_) );
  inv04 U1_2_2_8 ( .Y(g_array_3__8_), .A(g_array_2__8_) );
  nor02 U1_5_2_9 ( .Y(pog_array_3__9_), .A0(pog_array_2__8_), .A1(
        pog_array_2__9_) );
  inv04 U1_2_3_0 ( .Y(g_array_4__0_), .A(g_array_3__0_) );
  inv04 U1_2_3_2 ( .Y(g_array_4__2_), .A(g_array_3__2_) );
endmodule


module mul_24_DW02_mult_6_6_2 ( A, B, TC, PRODUCT );
  input [5:0] A;
  input [5:0] B;
  output [11:0] PRODUCT;
  input TC;
  wire   U1_level_node_0__5__3_, U1_level_node_1__4__0_,
         U1_level_node_1__5__0_, U1_level_node_1__5__1_,
         U1_level_node_1__5__2_, U1_level_node_1__6__0_,
         U1_level_node_1__6__1_, U1_level_node_1__6__2_,
         U1_level_node_1__7__0_, U1_level_node_1__7__1_,
         U1_level_node_1__8__0_, U1_level_node_2__3__0_,
         U1_level_node_2__4__0_, U1_level_node_2__4__1_,
         U1_level_node_2__5__0_, U1_level_node_2__5__1_,
         U1_level_node_2__6__0_, U1_level_node_2__6__1_,
         U1_level_node_2__7__0_, U1_level_node_2__7__1_,
         U1_level_node_2__8__0_, U1_level_node_2__8__1_,
         U1_level_node_2__9__0_, U1_level_node_3__2__0_,
         U1_level_node_3__3__0_, U1_level_node_3__3__1_,
         U1_level_node_3__4__0_, U1_level_node_3__4__1_,
         U1_level_node_3__5__0_, U1_level_node_3__5__1_,
         U1_level_node_3__6__0_, U1_level_node_3__6__1_,
         U1_level_node_3__7__0_, U1_level_node_3__7__1_,
         U1_level_node_3__8__0_, U1_level_node_3__8__1_,
         U1_level_node_3__9__0_, U1_level_node_3__9__1_,
         U1_level_node_3__10__0_, U1_B_neg_correction_1_, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303;

  or02 U5 ( .Y(n1), .A0(n298), .A1(n301) );
  inv01 U6 ( .Y(n2), .A(n1) );
  or02 U7 ( .Y(n3), .A0(n297), .A1(n300) );
  inv01 U8 ( .Y(n4), .A(n3) );
  or02 U9 ( .Y(n5), .A0(n299), .A1(n300) );
  inv01 U10 ( .Y(n6), .A(n5) );
  or02 U11 ( .Y(n7), .A0(n302), .A1(n303) );
  inv01 U12 ( .Y(n8), .A(n7) );
  or02 U13 ( .Y(n9), .A0(n294), .A1(n301) );
  inv01 U14 ( .Y(n10), .A(n9) );
  or02 U15 ( .Y(n11), .A0(n292), .A1(n301) );
  inv01 U16 ( .Y(n12), .A(n11) );
  or02 U17 ( .Y(n13), .A0(n296), .A1(n301) );
  inv01 U18 ( .Y(n14), .A(n13) );
  or02 U19 ( .Y(n15), .A0(n296), .A1(n299) );
  inv02 U20 ( .Y(n16), .A(n15) );
  or02 U21 ( .Y(n17), .A0(n298), .A1(n299) );
  inv02 U22 ( .Y(n18), .A(n17) );
  or02 U23 ( .Y(n19), .A0(n294), .A1(n299) );
  inv02 U24 ( .Y(n20), .A(n19) );
  nand02 U25 ( .Y(n21), .A0(n50), .A1(n44) );
  inv02 U26 ( .Y(n22), .A(n21) );
  nand02 U27 ( .Y(n23), .A0(n48), .A1(n46) );
  inv02 U28 ( .Y(n24), .A(n23) );
  inv01 U29 ( .Y(n25), .A(n173) );
  inv01 U30 ( .Y(n26), .A(n117) );
  inv01 U31 ( .Y(n27), .A(n175) );
  inv01 U32 ( .Y(n28), .A(n92) );
  or02 U33 ( .Y(n29), .A0(n293), .A1(n302) );
  inv02 U34 ( .Y(n30), .A(n29) );
  or02 U35 ( .Y(n31), .A0(n295), .A1(n300) );
  inv02 U36 ( .Y(n32), .A(n31) );
  or02 U37 ( .Y(n33), .A0(n293), .A1(n300) );
  inv02 U38 ( .Y(n34), .A(n33) );
  or02 U39 ( .Y(n35), .A0(n295), .A1(n302) );
  inv02 U40 ( .Y(n36), .A(n35) );
  or02 U41 ( .Y(n37), .A0(n297), .A1(n302) );
  inv02 U42 ( .Y(n38), .A(n37) );
  or02 U43 ( .Y(n39), .A0(n301), .A1(n302) );
  inv02 U44 ( .Y(n40), .A(n39) );
  buf02 U45 ( .Y(n41), .A(U1_level_node_2__4__1_) );
  buf02 U46 ( .Y(n42), .A(U1_level_node_2__3__0_) );
  buf02 U47 ( .Y(n43), .A(U1_level_node_0__5__3_) );
  buf02 U48 ( .Y(n44), .A(U1_level_node_0__5__3_) );
  buf02 U49 ( .Y(n45), .A(U1_B_neg_correction_1_) );
  buf02 U50 ( .Y(n46), .A(U1_B_neg_correction_1_) );
  or02 U51 ( .Y(n47), .A0(n299), .A1(n302) );
  inv02 U52 ( .Y(n48), .A(n47) );
  or02 U53 ( .Y(n49), .A0(n300), .A1(n303) );
  inv02 U54 ( .Y(n50), .A(n49) );
  or02 U55 ( .Y(n51), .A0(n297), .A1(n298) );
  inv02 U56 ( .Y(n52), .A(n51) );
  or02 U57 ( .Y(n53), .A0(n294), .A1(n303) );
  inv02 U58 ( .Y(n54), .A(n53) );
  or02 U59 ( .Y(n55), .A0(n292), .A1(n293) );
  inv02 U60 ( .Y(n56), .A(n55) );
  inv02 U61 ( .Y(U1_level_node_2__8__0_), .A(n57) );
  inv02 U62 ( .Y(U1_level_node_2__9__0_), .A(n58) );
  inv02 U63 ( .Y(n59), .A(n56) );
  inv02 U64 ( .Y(n60), .A(U1_level_node_1__8__0_) );
  inv02 U65 ( .Y(n61), .A(n54) );
  nor02 U66 ( .Y(n62), .A0(n59), .A1(n63) );
  nor02 U67 ( .Y(n64), .A0(n60), .A1(n65) );
  nor02 U68 ( .Y(n66), .A0(n61), .A1(n67) );
  nor02 U69 ( .Y(n68), .A0(n61), .A1(n69) );
  nor02 U70 ( .Y(n57), .A0(n70), .A1(n71) );
  nor02 U71 ( .Y(n72), .A0(n60), .A1(n61) );
  nor02 U72 ( .Y(n73), .A0(n59), .A1(n61) );
  nor02 U73 ( .Y(n74), .A0(n59), .A1(n60) );
  nor02 U74 ( .Y(n58), .A0(n74), .A1(n75) );
  nor02 U75 ( .Y(n76), .A0(U1_level_node_1__8__0_), .A1(n54) );
  inv01 U76 ( .Y(n63), .A(n76) );
  nor02 U77 ( .Y(n77), .A0(n56), .A1(n54) );
  inv01 U78 ( .Y(n65), .A(n77) );
  nor02 U79 ( .Y(n78), .A0(n56), .A1(U1_level_node_1__8__0_) );
  inv01 U80 ( .Y(n67), .A(n78) );
  nor02 U81 ( .Y(n79), .A0(n59), .A1(n60) );
  inv01 U82 ( .Y(n69), .A(n79) );
  nor02 U83 ( .Y(n80), .A0(n62), .A1(n64) );
  inv01 U84 ( .Y(n70), .A(n80) );
  nor02 U85 ( .Y(n81), .A0(n66), .A1(n68) );
  inv01 U86 ( .Y(n71), .A(n81) );
  nor02 U87 ( .Y(n82), .A0(n72), .A1(n73) );
  inv01 U88 ( .Y(n75), .A(n82) );
  or02 U89 ( .Y(n83), .A0(n292), .A1(n303) );
  inv02 U90 ( .Y(n84), .A(n83) );
  or02 U91 ( .Y(n85), .A0(n296), .A1(n297) );
  inv02 U92 ( .Y(n86), .A(n85) );
  or02 U93 ( .Y(n87), .A0(n295), .A1(n298) );
  inv02 U94 ( .Y(n88), .A(n87) );
  inv02 U95 ( .Y(U1_level_node_2__4__0_), .A(n89) );
  inv02 U96 ( .Y(U1_level_node_2__5__1_), .A(n90) );
  inv02 U97 ( .Y(n91), .A(n86) );
  inv02 U98 ( .Y(n92), .A(U1_level_node_1__4__0_) );
  inv02 U99 ( .Y(n93), .A(n88) );
  nor02 U100 ( .Y(n94), .A0(n91), .A1(n95) );
  nor02 U101 ( .Y(n96), .A0(n92), .A1(n97) );
  nor02 U102 ( .Y(n98), .A0(n93), .A1(n99) );
  nor02 U103 ( .Y(n100), .A0(n93), .A1(n101) );
  nor02 U104 ( .Y(n89), .A0(n102), .A1(n103) );
  nor02 U105 ( .Y(n104), .A0(n92), .A1(n93) );
  nor02 U106 ( .Y(n105), .A0(n91), .A1(n93) );
  nor02 U107 ( .Y(n106), .A0(n91), .A1(n92) );
  nor02 U108 ( .Y(n90), .A0(n106), .A1(n107) );
  nor02 U109 ( .Y(n108), .A0(U1_level_node_1__4__0_), .A1(n88) );
  inv01 U110 ( .Y(n95), .A(n108) );
  nor02 U111 ( .Y(n109), .A0(n86), .A1(n88) );
  inv01 U112 ( .Y(n97), .A(n109) );
  nor02 U113 ( .Y(n110), .A0(n86), .A1(n28) );
  inv01 U114 ( .Y(n99), .A(n110) );
  nor02 U115 ( .Y(n111), .A0(n91), .A1(n92) );
  inv01 U116 ( .Y(n101), .A(n111) );
  nor02 U117 ( .Y(n112), .A0(n94), .A1(n96) );
  inv01 U118 ( .Y(n102), .A(n112) );
  nor02 U119 ( .Y(n113), .A0(n98), .A1(n100) );
  inv01 U120 ( .Y(n103), .A(n113) );
  nor02 U121 ( .Y(n114), .A0(n104), .A1(n105) );
  inv01 U122 ( .Y(n107), .A(n114) );
  inv02 U123 ( .Y(U1_level_node_2__6__0_), .A(n115) );
  inv02 U124 ( .Y(U1_level_node_2__7__1_), .A(n116) );
  inv02 U125 ( .Y(n117), .A(U1_level_node_1__6__1_) );
  inv02 U126 ( .Y(n118), .A(U1_level_node_1__6__0_) );
  inv02 U127 ( .Y(n119), .A(U1_level_node_1__6__2_) );
  nor02 U128 ( .Y(n120), .A0(n117), .A1(n121) );
  nor02 U129 ( .Y(n122), .A0(n118), .A1(n123) );
  nor02 U130 ( .Y(n124), .A0(n119), .A1(n125) );
  nor02 U131 ( .Y(n126), .A0(n119), .A1(n127) );
  nor02 U132 ( .Y(n115), .A0(n128), .A1(n129) );
  nor02 U133 ( .Y(n130), .A0(n118), .A1(n119) );
  nor02 U134 ( .Y(n131), .A0(n117), .A1(n119) );
  nor02 U135 ( .Y(n132), .A0(n117), .A1(n118) );
  nor02 U136 ( .Y(n116), .A0(n132), .A1(n133) );
  nor02 U137 ( .Y(n134), .A0(U1_level_node_1__6__0_), .A1(
        U1_level_node_1__6__2_) );
  inv01 U138 ( .Y(n121), .A(n134) );
  nor02 U139 ( .Y(n135), .A0(n26), .A1(U1_level_node_1__6__2_) );
  inv01 U140 ( .Y(n123), .A(n135) );
  nor02 U141 ( .Y(n136), .A0(U1_level_node_1__6__1_), .A1(
        U1_level_node_1__6__0_) );
  inv01 U142 ( .Y(n125), .A(n136) );
  nor02 U143 ( .Y(n137), .A0(n117), .A1(n118) );
  inv01 U144 ( .Y(n127), .A(n137) );
  nor02 U145 ( .Y(n138), .A0(n120), .A1(n122) );
  inv01 U146 ( .Y(n128), .A(n138) );
  nor02 U147 ( .Y(n139), .A0(n124), .A1(n126) );
  inv01 U148 ( .Y(n129), .A(n139) );
  nor02 U149 ( .Y(n140), .A0(n130), .A1(n131) );
  inv01 U150 ( .Y(n133), .A(n140) );
  or02 U151 ( .Y(n141), .A0(n295), .A1(n296) );
  inv02 U152 ( .Y(n142), .A(n141) );
  or02 U153 ( .Y(n143), .A0(n294), .A1(n297) );
  inv02 U154 ( .Y(n144), .A(n143) );
  inv02 U155 ( .Y(U1_level_node_1__5__0_), .A(n145) );
  inv02 U156 ( .Y(U1_level_node_1__6__2_), .A(n146) );
  inv02 U157 ( .Y(n147), .A(n144) );
  inv02 U158 ( .Y(n148), .A(n286) );
  inv02 U159 ( .Y(n149), .A(n142) );
  nor02 U160 ( .Y(n150), .A0(n147), .A1(n151) );
  nor02 U161 ( .Y(n152), .A0(n148), .A1(n153) );
  nor02 U162 ( .Y(n154), .A0(n149), .A1(n155) );
  nor02 U163 ( .Y(n156), .A0(n149), .A1(n157) );
  nor02 U164 ( .Y(n145), .A0(n158), .A1(n159) );
  nor02 U165 ( .Y(n160), .A0(n148), .A1(n149) );
  nor02 U166 ( .Y(n161), .A0(n147), .A1(n149) );
  nor02 U167 ( .Y(n162), .A0(n147), .A1(n148) );
  nor02 U168 ( .Y(n146), .A0(n162), .A1(n163) );
  nor02 U169 ( .Y(n164), .A0(n286), .A1(n142) );
  inv01 U170 ( .Y(n151), .A(n164) );
  nor02 U171 ( .Y(n165), .A0(n144), .A1(n142) );
  inv01 U172 ( .Y(n153), .A(n165) );
  nor02 U173 ( .Y(n166), .A0(n144), .A1(n286) );
  inv01 U174 ( .Y(n155), .A(n166) );
  nor02 U175 ( .Y(n167), .A0(n147), .A1(n148) );
  inv01 U176 ( .Y(n157), .A(n167) );
  nor02 U177 ( .Y(n168), .A0(n150), .A1(n152) );
  inv01 U178 ( .Y(n158), .A(n168) );
  nor02 U179 ( .Y(n169), .A0(n154), .A1(n156) );
  inv01 U180 ( .Y(n159), .A(n169) );
  nor02 U181 ( .Y(n170), .A0(n160), .A1(n161) );
  inv01 U182 ( .Y(n163), .A(n170) );
  inv02 U183 ( .Y(U1_level_node_2__5__0_), .A(n171) );
  inv02 U184 ( .Y(U1_level_node_2__6__1_), .A(n172) );
  inv02 U185 ( .Y(n173), .A(U1_level_node_1__5__1_) );
  inv02 U186 ( .Y(n174), .A(U1_level_node_1__5__0_) );
  inv02 U187 ( .Y(n175), .A(U1_level_node_1__5__2_) );
  nor02 U188 ( .Y(n176), .A0(n173), .A1(n177) );
  nor02 U189 ( .Y(n178), .A0(n174), .A1(n179) );
  nor02 U190 ( .Y(n180), .A0(n175), .A1(n181) );
  nor02 U191 ( .Y(n182), .A0(n175), .A1(n183) );
  nor02 U192 ( .Y(n171), .A0(n184), .A1(n185) );
  nor02 U193 ( .Y(n186), .A0(n174), .A1(n175) );
  nor02 U194 ( .Y(n187), .A0(n173), .A1(n175) );
  nor02 U195 ( .Y(n188), .A0(n173), .A1(n174) );
  nor02 U196 ( .Y(n172), .A0(n188), .A1(n189) );
  nor02 U197 ( .Y(n190), .A0(U1_level_node_1__5__0_), .A1(
        U1_level_node_1__5__2_) );
  inv01 U198 ( .Y(n177), .A(n190) );
  nor02 U199 ( .Y(n191), .A0(n25), .A1(n27) );
  inv01 U200 ( .Y(n179), .A(n191) );
  nor02 U201 ( .Y(n192), .A0(U1_level_node_1__5__1_), .A1(
        U1_level_node_1__5__0_) );
  inv01 U202 ( .Y(n181), .A(n192) );
  nor02 U203 ( .Y(n193), .A0(n173), .A1(n174) );
  inv01 U204 ( .Y(n183), .A(n193) );
  nor02 U205 ( .Y(n194), .A0(n176), .A1(n178) );
  inv01 U206 ( .Y(n184), .A(n194) );
  nor02 U207 ( .Y(n195), .A0(n180), .A1(n182) );
  inv01 U208 ( .Y(n185), .A(n195) );
  nor02 U209 ( .Y(n196), .A0(n186), .A1(n187) );
  inv01 U210 ( .Y(n189), .A(n196) );
  or02 U211 ( .Y(n197), .A0(n293), .A1(n296) );
  inv02 U212 ( .Y(n198), .A(n197) );
  or02 U213 ( .Y(n199), .A0(n296), .A1(n303) );
  inv02 U214 ( .Y(n200), .A(n199) );
  or02 U215 ( .Y(n201), .A0(n293), .A1(n294) );
  inv02 U216 ( .Y(n202), .A(n201) );
  or02 U217 ( .Y(n203), .A0(n294), .A1(n295) );
  inv02 U218 ( .Y(n204), .A(n203) );
  inv02 U219 ( .Y(U1_level_node_1__7__0_), .A(n205) );
  inv02 U220 ( .Y(U1_level_node_1__8__0_), .A(n206) );
  inv02 U221 ( .Y(n207), .A(n202) );
  inv02 U222 ( .Y(n208), .A(n284) );
  inv02 U223 ( .Y(n209), .A(n200) );
  nor02 U224 ( .Y(n210), .A0(n207), .A1(n211) );
  nor02 U225 ( .Y(n212), .A0(n208), .A1(n213) );
  nor02 U226 ( .Y(n214), .A0(n209), .A1(n215) );
  nor02 U227 ( .Y(n216), .A0(n209), .A1(n217) );
  nor02 U228 ( .Y(n205), .A0(n218), .A1(n219) );
  nor02 U229 ( .Y(n220), .A0(n208), .A1(n209) );
  nor02 U230 ( .Y(n221), .A0(n207), .A1(n209) );
  nor02 U231 ( .Y(n222), .A0(n207), .A1(n208) );
  nor02 U232 ( .Y(n206), .A0(n222), .A1(n223) );
  nor02 U233 ( .Y(n224), .A0(n284), .A1(n200) );
  inv01 U234 ( .Y(n211), .A(n224) );
  nor02 U235 ( .Y(n225), .A0(n202), .A1(n200) );
  inv01 U236 ( .Y(n213), .A(n225) );
  nor02 U237 ( .Y(n226), .A0(n202), .A1(n284) );
  inv01 U238 ( .Y(n215), .A(n226) );
  nor02 U239 ( .Y(n227), .A0(n207), .A1(n208) );
  inv01 U240 ( .Y(n217), .A(n227) );
  nor02 U241 ( .Y(n228), .A0(n210), .A1(n212) );
  inv01 U242 ( .Y(n218), .A(n228) );
  nor02 U243 ( .Y(n229), .A0(n214), .A1(n216) );
  inv01 U244 ( .Y(n219), .A(n229) );
  nor02 U245 ( .Y(n230), .A0(n220), .A1(n221) );
  inv01 U246 ( .Y(n223), .A(n230) );
  inv02 U247 ( .Y(U1_level_node_1__6__0_), .A(n231) );
  inv02 U248 ( .Y(U1_level_node_1__7__1_), .A(n232) );
  inv02 U249 ( .Y(n233), .A(n204) );
  inv02 U250 ( .Y(n234), .A(n288) );
  inv02 U251 ( .Y(n235), .A(n198) );
  nor02 U252 ( .Y(n236), .A0(n233), .A1(n237) );
  nor02 U253 ( .Y(n238), .A0(n234), .A1(n239) );
  nor02 U254 ( .Y(n240), .A0(n235), .A1(n241) );
  nor02 U255 ( .Y(n242), .A0(n235), .A1(n243) );
  nor02 U256 ( .Y(n231), .A0(n244), .A1(n245) );
  nor02 U257 ( .Y(n246), .A0(n234), .A1(n235) );
  nor02 U258 ( .Y(n247), .A0(n233), .A1(n235) );
  nor02 U259 ( .Y(n248), .A0(n233), .A1(n234) );
  nor02 U260 ( .Y(n232), .A0(n248), .A1(n249) );
  nor02 U261 ( .Y(n250), .A0(n288), .A1(n198) );
  inv01 U262 ( .Y(n237), .A(n250) );
  nor02 U263 ( .Y(n251), .A0(n204), .A1(n198) );
  inv01 U264 ( .Y(n239), .A(n251) );
  nor02 U265 ( .Y(n252), .A0(n204), .A1(n288) );
  inv01 U266 ( .Y(n241), .A(n252) );
  nor02 U267 ( .Y(n253), .A0(n233), .A1(n234) );
  inv01 U268 ( .Y(n243), .A(n253) );
  nor02 U269 ( .Y(n254), .A0(n236), .A1(n238) );
  inv01 U270 ( .Y(n244), .A(n254) );
  nor02 U271 ( .Y(n255), .A0(n240), .A1(n242) );
  inv01 U272 ( .Y(n245), .A(n255) );
  nor02 U273 ( .Y(n256), .A0(n246), .A1(n247) );
  inv01 U274 ( .Y(n249), .A(n256) );
  inv02 U275 ( .Y(U1_level_node_2__7__0_), .A(n257) );
  inv02 U276 ( .Y(U1_level_node_2__8__1_), .A(n258) );
  inv02 U277 ( .Y(n259), .A(U1_level_node_1__7__1_) );
  inv02 U278 ( .Y(n260), .A(U1_level_node_1__7__0_) );
  inv02 U279 ( .Y(n261), .A(n24) );
  nor02 U280 ( .Y(n262), .A0(n259), .A1(n263) );
  nor02 U281 ( .Y(n264), .A0(n260), .A1(n265) );
  nor02 U282 ( .Y(n266), .A0(n261), .A1(n267) );
  nor02 U283 ( .Y(n268), .A0(n261), .A1(n269) );
  nor02 U284 ( .Y(n257), .A0(n270), .A1(n271) );
  nor02 U285 ( .Y(n272), .A0(n260), .A1(n261) );
  nor02 U286 ( .Y(n273), .A0(n259), .A1(n261) );
  nor02 U287 ( .Y(n274), .A0(n259), .A1(n260) );
  nor02 U288 ( .Y(n258), .A0(n274), .A1(n275) );
  nor02 U289 ( .Y(n276), .A0(U1_level_node_1__7__0_), .A1(n24) );
  inv01 U290 ( .Y(n263), .A(n276) );
  nor02 U291 ( .Y(n277), .A0(U1_level_node_1__7__1_), .A1(n24) );
  inv01 U292 ( .Y(n265), .A(n277) );
  nor02 U293 ( .Y(n278), .A0(U1_level_node_1__7__1_), .A1(
        U1_level_node_1__7__0_) );
  inv01 U294 ( .Y(n267), .A(n278) );
  nor02 U295 ( .Y(n279), .A0(n259), .A1(n260) );
  inv01 U296 ( .Y(n269), .A(n279) );
  nor02 U297 ( .Y(n280), .A0(n262), .A1(n264) );
  inv01 U298 ( .Y(n270), .A(n280) );
  nor02 U299 ( .Y(n281), .A0(n266), .A1(n268) );
  inv01 U300 ( .Y(n271), .A(n281) );
  nor02 U301 ( .Y(n282), .A0(n272), .A1(n273) );
  inv01 U302 ( .Y(n275), .A(n282) );
  or02 U303 ( .Y(n283), .A0(n292), .A1(n295) );
  inv02 U304 ( .Y(n284), .A(n283) );
  or02 U305 ( .Y(n285), .A0(n292), .A1(n299) );
  inv02 U306 ( .Y(n286), .A(n285) );
  or02 U307 ( .Y(n287), .A0(n292), .A1(n297) );
  inv02 U308 ( .Y(n288), .A(n287) );
  or02 U309 ( .Y(n289), .A0(n300), .A1(n301) );
  inv02 U310 ( .Y(PRODUCT[0]), .A(n289) );
  inv02 U311 ( .Y(n292), .A(A[4]) );
  inv02 U312 ( .Y(n296), .A(A[2]) );
  inv02 U313 ( .Y(n299), .A(B[1]) );
  inv02 U314 ( .Y(n295), .A(B[3]) );
  inv02 U315 ( .Y(n298), .A(A[1]) );
  inv02 U316 ( .Y(n297), .A(B[2]) );
  inv02 U317 ( .Y(n301), .A(B[0]) );
  inv02 U318 ( .Y(n303), .A(B[5]) );
  inv02 U319 ( .Y(n302), .A(A[5]) );
  inv02 U320 ( .Y(n293), .A(B[4]) );
  inv02 U321 ( .Y(n300), .A(A[0]) );
  inv02 U322 ( .Y(n294), .A(A[3]) );
  xor2 U323 ( .Y(U1_level_node_1__5__1_), .A0(n43), .A1(n50) );
  xor2 U324 ( .Y(U1_level_node_1__6__1_), .A0(n45), .A1(n48) );
  mul_24_DW01_add_11_2 U1_U9720 ( .A({1'b0, U1_level_node_3__10__0_, 
        U1_level_node_3__9__0_, U1_level_node_3__8__0_, U1_level_node_3__7__0_, 
        U1_level_node_3__6__0_, U1_level_node_3__5__0_, U1_level_node_3__4__0_, 
        U1_level_node_3__3__0_, U1_level_node_3__2__0_, n2}), .B({1'b0, n8, 
        U1_level_node_3__9__1_, U1_level_node_3__8__1_, U1_level_node_3__7__1_, 
        U1_level_node_3__6__1_, U1_level_node_3__5__1_, U1_level_node_3__4__1_, 
        U1_level_node_3__3__1_, n4, n6}), .CI(1'b0), .SUM(PRODUCT[11:1]) );
  nor02 U325 ( .Y(U1_level_node_0__5__3_), .A0(n293), .A1(n298) );
  nor02 U326 ( .Y(U1_B_neg_correction_1_), .A0(n298), .A1(n303) );
  hadd1 U1_U3220_1_4 ( .S(U1_level_node_1__4__0_), .CO(U1_level_node_1__5__2_), 
        .A(n12), .B(n20) );
  hadd1 U1_U3220_2_3 ( .S(U1_level_node_2__3__0_), .CO(U1_level_node_2__4__1_), 
        .A(n10), .B(n16) );
  fadd1 U1_U3140_3_9_0 ( .S(U1_level_node_3__9__0_), .CO(
        U1_level_node_3__10__0_), .A(U1_level_node_2__9__0_), .B(n84), .CI(n30) );
  fadd1 U1_U3140_3_8_0 ( .S(U1_level_node_3__8__0_), .CO(
        U1_level_node_3__9__1_), .A(U1_level_node_2__8__0_), .B(
        U1_level_node_2__8__1_), .CI(n36) );
  fadd1 U1_U3140_3_7_0 ( .S(U1_level_node_3__7__0_), .CO(
        U1_level_node_3__8__1_), .A(U1_level_node_2__7__0_), .B(
        U1_level_node_2__7__1_), .CI(n38) );
  fadd1 U1_U3140_3_6_0 ( .S(U1_level_node_3__6__0_), .CO(
        U1_level_node_3__7__1_), .A(U1_level_node_2__6__0_), .B(
        U1_level_node_2__6__1_), .CI(n22) );
  fadd1 U1_U3140_3_5_0 ( .S(U1_level_node_3__5__0_), .CO(
        U1_level_node_3__6__1_), .A(U1_level_node_2__5__0_), .B(
        U1_level_node_2__5__1_), .CI(n40) );
  fadd1 U1_U3140_3_4_0 ( .S(U1_level_node_3__4__0_), .CO(
        U1_level_node_3__5__1_), .A(U1_level_node_2__4__0_), .B(n41), .CI(n34)
         );
  fadd1 U1_U3140_3_3_0 ( .S(U1_level_node_3__3__0_), .CO(
        U1_level_node_3__4__1_), .A(n42), .B(n52), .CI(n32) );
  hadd1 U1_U3220_3_2 ( .S(U1_level_node_3__2__0_), .CO(U1_level_node_3__3__1_), 
        .A(n14), .B(n18) );
endmodule


module mul_24_DW01_add_11_1 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   g_array_0__9_, g_array_0__8_, g_array_0__7_, g_array_0__6_,
         g_array_0__5_, g_array_0__4_, g_array_0__3_, g_array_0__2_,
         g_array_0__1_, g_array_0__0_, g_array_1__9_, g_array_1__8_,
         g_array_1__7_, g_array_1__6_, g_array_1__5_, g_array_1__4_,
         g_array_1__3_, g_array_1__2_, g_array_1__1_, g_array_1__0_,
         g_array_2__9_, g_array_2__8_, g_array_2__7_, g_array_2__6_,
         g_array_2__5_, g_array_2__4_, g_array_2__3_, g_array_2__2_,
         g_array_2__1_, g_array_2__0_, g_array_3__9_, g_array_3__8_,
         g_array_3__7_, g_array_3__6_, g_array_3__5_, g_array_3__4_,
         g_array_3__3_, g_array_3__2_, g_array_3__1_, g_array_3__0_,
         g_array_4__9_, g_array_4__6_, g_array_4__5_, g_array_4__2_,
         g_array_4__1_, g_array_4__0_, pog_array_0__9_, pog_array_0__0_,
         pog_array_1__9_, pog_array_1__8_, pog_array_1__7_, pog_array_1__6_,
         pog_array_1__5_, pog_array_1__3_, pog_array_1__2_, pog_array_1__1_,
         pog_array_2__9_, pog_array_2__8_, pog_array_2__7_, pog_array_2__6_,
         pog_array_2__5_, pog_array_2__4_, pog_array_2__3_, pog_array_2__1_,
         pog_array_3__9_, pog_array_3__8_, pog_array_3__7_, pog_array_3__5_,
         pog_array_3__4_, pog_array_3__3_, part_sum_9_, part_sum_8_,
         part_sum_7_, part_sum_6_, part_sum_5_, part_sum_4_, part_sum_3_,
         part_sum_2_, part_sum_1_, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n84, n86, n88, n90, n92, n94, n96, n98, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131;

  inv02 U1_2_0_7 ( .Y(g_array_1__7_), .A(g_array_0__7_) );
  inv02 U1_2_0_5 ( .Y(g_array_1__5_), .A(g_array_0__5_) );
  inv02 U7 ( .Y(part_sum_5_), .A(n121) );
  inv02 U8 ( .Y(part_sum_7_), .A(n119) );
  inv01 U9 ( .Y(g_array_3__5_), .A(n31) );
  nor02 U10 ( .Y(n32), .A0(pog_array_2__5_), .A1(g_array_2__4_) );
  inv01 U11 ( .Y(n33), .A(g_array_2__5_) );
  nor02 U12 ( .Y(n31), .A0(n32), .A1(n33) );
  inv02 U1_3_1_5 ( .Y(pog_array_2__5_), .A(pog_array_1__5_) );
  inv02 U1_2_1_5 ( .Y(g_array_2__5_), .A(g_array_1__5_) );
  inv01 U13 ( .Y(g_array_3__9_), .A(n34) );
  nor02 U14 ( .Y(n35), .A0(pog_array_2__9_), .A1(g_array_2__8_) );
  inv01 U15 ( .Y(n36), .A(g_array_2__9_) );
  nor02 U16 ( .Y(n34), .A0(n35), .A1(n36) );
  inv02 U1_3_1_9 ( .Y(pog_array_2__9_), .A(pog_array_1__9_) );
  inv02 U1_2_1_9 ( .Y(g_array_2__9_), .A(g_array_1__9_) );
  inv01 U17 ( .Y(g_array_1__2_), .A(n37) );
  nor02 U18 ( .Y(n38), .A0(n106), .A1(g_array_0__1_) );
  inv01 U19 ( .Y(n39), .A(g_array_0__2_) );
  nor02 U20 ( .Y(n37), .A0(n38), .A1(n39) );
  nand02 U21 ( .Y(g_array_1__6_), .A0(n40), .A1(g_array_0__6_) );
  inv01 U22 ( .Y(n41), .A(g_array_0__5_) );
  inv01 U23 ( .Y(n42), .A(n112) );
  nand02 U24 ( .Y(n40), .A0(n41), .A1(n42) );
  nand02 U25 ( .Y(g_array_4__9_), .A0(n43), .A1(n44) );
  inv01 U26 ( .Y(n45), .A(g_array_3__9_) );
  inv01 U27 ( .Y(n46), .A(g_array_3__6_) );
  inv01 U28 ( .Y(n47), .A(pog_array_3__9_) );
  nand02 U29 ( .Y(n43), .A0(n45), .A1(n46) );
  nand02 U30 ( .Y(n44), .A0(n45), .A1(n47) );
  inv02 U1_2_0_9 ( .Y(g_array_1__9_), .A(g_array_0__9_) );
  inv02 U1_3_1_8 ( .Y(pog_array_2__8_), .A(pog_array_1__8_) );
  inv02 U1_3_0_9 ( .Y(pog_array_1__9_), .A(pog_array_0__9_) );
  inv02 U31 ( .Y(n127), .A(pog_array_0__0_) );
  inv01 U32 ( .Y(g_array_3__1_), .A(n48) );
  nor02 U33 ( .Y(n49), .A0(pog_array_2__1_), .A1(g_array_2__0_) );
  inv01 U34 ( .Y(n50), .A(g_array_2__1_) );
  nor02 U35 ( .Y(n48), .A0(n49), .A1(n50) );
  inv01 U1_2_3_1 ( .Y(g_array_4__1_), .A(g_array_3__1_) );
  inv02 U1_3_1_1 ( .Y(pog_array_2__1_), .A(pog_array_1__1_) );
  inv02 U1_2_1_0 ( .Y(g_array_2__0_), .A(g_array_1__0_) );
  inv02 U1_2_1_1 ( .Y(g_array_2__1_), .A(g_array_1__1_) );
  nand02 U36 ( .Y(g_array_1__8_), .A0(n51), .A1(g_array_0__8_) );
  inv01 U37 ( .Y(n52), .A(g_array_0__7_) );
  inv01 U38 ( .Y(n53), .A(n110) );
  nand02 U39 ( .Y(n51), .A0(n52), .A1(n53) );
  inv02 U1_2_1_8 ( .Y(g_array_2__8_), .A(g_array_1__8_) );
  ao21 U40 ( .Y(n54), .A0(pog_array_3__7_), .A1(g_array_3__6_), .B0(
        g_array_3__7_) );
  inv01 U41 ( .Y(n55), .A(n54) );
  ao21 U42 ( .Y(n56), .A0(pog_array_3__8_), .A1(g_array_3__6_), .B0(
        g_array_3__8_) );
  inv01 U43 ( .Y(n57), .A(n56) );
  inv02 U44 ( .Y(SUM[10]), .A(g_array_4__9_) );
  nand02 U45 ( .Y(g_array_4__5_), .A0(n58), .A1(n59) );
  inv01 U46 ( .Y(n60), .A(g_array_3__5_) );
  inv01 U47 ( .Y(n61), .A(g_array_3__2_) );
  inv01 U48 ( .Y(n62), .A(pog_array_3__5_) );
  nand02 U49 ( .Y(n58), .A0(n60), .A1(n61) );
  nand02 U50 ( .Y(n59), .A0(n60), .A1(n62) );
  ao21 U51 ( .Y(n63), .A0(pog_array_3__3_), .A1(g_array_3__2_), .B0(
        g_array_3__3_) );
  inv01 U52 ( .Y(n64), .A(n63) );
  ao21 U53 ( .Y(n65), .A0(pog_array_3__4_), .A1(g_array_3__2_), .B0(
        g_array_3__4_) );
  inv01 U54 ( .Y(n66), .A(n65) );
  inv02 U1_2_0_3 ( .Y(g_array_1__3_), .A(g_array_0__3_) );
  inv01 U1_2_0_1 ( .Y(g_array_1__1_), .A(g_array_0__1_) );
  nand02 U55 ( .Y(g_array_1__4_), .A0(n67), .A1(g_array_0__4_) );
  inv01 U56 ( .Y(n68), .A(g_array_0__3_) );
  inv01 U57 ( .Y(n69), .A(n108) );
  nand02 U58 ( .Y(n67), .A0(n68), .A1(n69) );
  inv02 U1_2_1_4 ( .Y(g_array_2__4_), .A(g_array_1__4_) );
  or02 U59 ( .Y(n70), .A0(A[3]), .A1(B[3]) );
  inv01 U60 ( .Y(n71), .A(n70) );
  inv02 U1_3_0_3 ( .Y(pog_array_1__3_), .A(n71) );
  or02 U61 ( .Y(n72), .A0(A[5]), .A1(B[5]) );
  inv01 U62 ( .Y(n73), .A(n72) );
  inv01 U63 ( .Y(n74), .A(n72) );
  inv02 U1_3_0_5 ( .Y(pog_array_1__5_), .A(n73) );
  or02 U64 ( .Y(n75), .A0(A[7]), .A1(B[7]) );
  inv01 U65 ( .Y(n76), .A(n75) );
  inv01 U66 ( .Y(n77), .A(n75) );
  inv02 U1_3_0_7 ( .Y(pog_array_1__7_), .A(n76) );
  or02 U67 ( .Y(n78), .A0(A[1]), .A1(B[1]) );
  inv01 U68 ( .Y(n79), .A(n78) );
  inv02 U1_3_0_1 ( .Y(pog_array_1__1_), .A(n79) );
  or02 U69 ( .Y(n80), .A0(n71), .A1(n108) );
  inv01 U70 ( .Y(n81), .A(n80) );
  inv02 U1_3_1_4 ( .Y(pog_array_2__4_), .A(n81) );
  xor2 U71 ( .Y(n82), .A0(part_sum_8_), .A1(n55) );
  inv02 U72 ( .Y(SUM[8]), .A(n82) );
  xor2 U73 ( .Y(n84), .A0(part_sum_4_), .A1(n64) );
  inv02 U74 ( .Y(SUM[4]), .A(n84) );
  xor2 U75 ( .Y(n86), .A0(part_sum_6_), .A1(g_array_4__5_) );
  inv02 U76 ( .Y(SUM[6]), .A(n86) );
  xor2 U77 ( .Y(n88), .A0(part_sum_2_), .A1(g_array_4__1_) );
  inv02 U78 ( .Y(SUM[2]), .A(n88) );
  xor2 U79 ( .Y(n90), .A0(part_sum_9_), .A1(n57) );
  inv02 U80 ( .Y(SUM[9]), .A(n90) );
  xor2 U81 ( .Y(n92), .A0(part_sum_7_), .A1(g_array_4__6_) );
  inv02 U82 ( .Y(SUM[7]), .A(n92) );
  xor2 U83 ( .Y(n94), .A0(part_sum_5_), .A1(n66) );
  inv02 U84 ( .Y(SUM[5]), .A(n94) );
  xor2 U85 ( .Y(n96), .A0(part_sum_3_), .A1(g_array_4__2_) );
  inv02 U86 ( .Y(SUM[3]), .A(n96) );
  xor2 U87 ( .Y(n98), .A0(part_sum_1_), .A1(g_array_4__0_) );
  inv02 U88 ( .Y(SUM[1]), .A(n98) );
  nand02 U89 ( .Y(g_array_2__2_), .A0(n100), .A1(n101) );
  inv01 U90 ( .Y(n102), .A(g_array_1__2_) );
  inv01 U91 ( .Y(n103), .A(g_array_1__0_) );
  inv01 U92 ( .Y(n104), .A(pog_array_1__2_) );
  nand02 U93 ( .Y(n100), .A0(n102), .A1(n103) );
  nand02 U94 ( .Y(n101), .A0(n102), .A1(n104) );
  inv02 U1_2_2_2 ( .Y(g_array_3__2_), .A(g_array_2__2_) );
  inv02 U95 ( .Y(g_array_1__0_), .A(g_array_0__0_) );
  or02 U96 ( .Y(n105), .A0(A[2]), .A1(B[2]) );
  inv02 U97 ( .Y(n106), .A(n105) );
  inv01 U98 ( .Y(n128), .A(n106) );
  or02 U99 ( .Y(n107), .A0(A[4]), .A1(B[4]) );
  inv02 U100 ( .Y(n108), .A(n107) );
  or02 U101 ( .Y(n109), .A0(A[8]), .A1(B[8]) );
  inv02 U102 ( .Y(n110), .A(n109) );
  inv01 U103 ( .Y(n129), .A(n108) );
  inv01 U104 ( .Y(n131), .A(n110) );
  or02 U105 ( .Y(n111), .A0(A[6]), .A1(B[6]) );
  inv01 U106 ( .Y(n112), .A(n111) );
  inv01 U107 ( .Y(n113), .A(n111) );
  inv01 U108 ( .Y(n130), .A(n112) );
  inv02 U109 ( .Y(g_array_3__6_), .A(n114) );
  nor02 U110 ( .Y(n115), .A0(pog_array_2__6_), .A1(g_array_2__2_) );
  inv01 U111 ( .Y(n116), .A(g_array_2__6_) );
  nor02 U112 ( .Y(n114), .A0(n115), .A1(n116) );
  inv01 U1_2_3_6 ( .Y(g_array_4__6_), .A(g_array_3__6_) );
  inv04 U113 ( .Y(part_sum_9_), .A(n117) );
  inv04 U114 ( .Y(part_sum_8_), .A(n118) );
  inv04 U115 ( .Y(part_sum_6_), .A(n120) );
  inv04 U116 ( .Y(part_sum_4_), .A(n122) );
  inv04 U117 ( .Y(part_sum_3_), .A(n123) );
  inv04 U118 ( .Y(part_sum_2_), .A(n124) );
  inv04 U119 ( .Y(part_sum_1_), .A(n125) );
  inv04 U120 ( .Y(SUM[0]), .A(n126) );
  nand02 U0_1_0 ( .Y(g_array_0__0_), .A0(A[0]), .A1(B[0]) );
  nor02 U0_2_0 ( .Y(pog_array_0__0_), .A0(A[0]), .A1(B[0]) );
  nand02 U0_3_0 ( .Y(n126), .A0(g_array_0__0_), .A1(n127) );
  nand02 U0_1_1 ( .Y(g_array_0__1_), .A0(A[1]), .A1(B[1]) );
  nand02 U0_3_1 ( .Y(n125), .A0(g_array_0__1_), .A1(pog_array_1__1_) );
  nand02 U0_1_2 ( .Y(g_array_0__2_), .A0(A[2]), .A1(B[2]) );
  nand02 U0_3_2 ( .Y(n124), .A0(g_array_0__2_), .A1(n128) );
  nand02 U0_1_3 ( .Y(g_array_0__3_), .A0(A[3]), .A1(B[3]) );
  nand02 U0_3_3 ( .Y(n123), .A0(g_array_0__3_), .A1(pog_array_1__3_) );
  nand02 U0_1_4 ( .Y(g_array_0__4_), .A0(A[4]), .A1(B[4]) );
  nand02 U0_3_4 ( .Y(n122), .A0(g_array_0__4_), .A1(n129) );
  nand02 U0_1_5 ( .Y(g_array_0__5_), .A0(A[5]), .A1(B[5]) );
  nand02 U0_3_5 ( .Y(n121), .A0(g_array_0__5_), .A1(pog_array_1__5_) );
  nand02 U0_1_6 ( .Y(g_array_0__6_), .A0(A[6]), .A1(B[6]) );
  nand02 U0_3_6 ( .Y(n120), .A0(g_array_0__6_), .A1(n130) );
  nand02 U0_1_7 ( .Y(g_array_0__7_), .A0(A[7]), .A1(B[7]) );
  nand02 U0_3_7 ( .Y(n119), .A0(g_array_0__7_), .A1(pog_array_1__7_) );
  nand02 U0_1_8 ( .Y(g_array_0__8_), .A0(A[8]), .A1(B[8]) );
  nand02 U0_3_8 ( .Y(n118), .A0(g_array_0__8_), .A1(n131) );
  nand02 U0_1_9 ( .Y(g_array_0__9_), .A0(A[9]), .A1(B[9]) );
  nor02 U0_2_9 ( .Y(pog_array_0__9_), .A0(A[9]), .A1(B[9]) );
  nand02 U0_3_9 ( .Y(n117), .A0(g_array_0__9_), .A1(pog_array_1__9_) );
  nor02 U1_5_0_2 ( .Y(pog_array_1__2_), .A0(n79), .A1(n106) );
  nor02 U1_5_0_6 ( .Y(pog_array_1__6_), .A0(n74), .A1(n113) );
  nor02 U1_5_0_8 ( .Y(pog_array_1__8_), .A0(n77), .A1(n110) );
  inv04 U1_2_1_3 ( .Y(g_array_2__3_), .A(g_array_1__3_) );
  inv04 U1_3_1_3 ( .Y(pog_array_2__3_), .A(pog_array_1__3_) );
  aoi21 U1_4_1_6 ( .Y(g_array_2__6_), .A0(pog_array_1__6_), .A1(g_array_1__4_), 
        .B0(g_array_1__6_) );
  nand02 U1_5_1_6 ( .Y(pog_array_2__6_), .A0(pog_array_1__6_), .A1(n81) );
  inv04 U1_2_1_7 ( .Y(g_array_2__7_), .A(g_array_1__7_) );
  inv04 U1_3_1_7 ( .Y(pog_array_2__7_), .A(pog_array_1__7_) );
  inv04 U1_2_2_0 ( .Y(g_array_3__0_), .A(g_array_2__0_) );
  inv04 U1_2_2_3 ( .Y(g_array_3__3_), .A(g_array_2__3_) );
  inv04 U1_3_2_3 ( .Y(pog_array_3__3_), .A(pog_array_2__3_) );
  inv04 U1_2_2_4 ( .Y(g_array_3__4_), .A(g_array_2__4_) );
  inv04 U1_3_2_4 ( .Y(pog_array_3__4_), .A(pog_array_2__4_) );
  nor02 U1_5_2_5 ( .Y(pog_array_3__5_), .A0(pog_array_2__4_), .A1(
        pog_array_2__5_) );
  inv04 U1_2_2_7 ( .Y(g_array_3__7_), .A(g_array_2__7_) );
  inv04 U1_3_2_7 ( .Y(pog_array_3__7_), .A(pog_array_2__7_) );
  inv04 U1_2_2_8 ( .Y(g_array_3__8_), .A(g_array_2__8_) );
  inv04 U1_3_2_8 ( .Y(pog_array_3__8_), .A(pog_array_2__8_) );
  nor02 U1_5_2_9 ( .Y(pog_array_3__9_), .A0(pog_array_2__8_), .A1(
        pog_array_2__9_) );
  inv04 U1_2_3_0 ( .Y(g_array_4__0_), .A(g_array_3__0_) );
  inv04 U1_2_3_2 ( .Y(g_array_4__2_), .A(g_array_3__2_) );
endmodule


module mul_24_DW02_mult_6_6_1 ( A, B, TC, PRODUCT );
  input [5:0] A;
  input [5:0] B;
  output [11:0] PRODUCT;
  input TC;
  wire   U1_level_node_0__5__3_, U1_level_node_0__6__1_,
         U1_level_node_1__4__0_, U1_level_node_1__5__0_,
         U1_level_node_1__5__1_, U1_level_node_1__5__2_,
         U1_level_node_1__6__0_, U1_level_node_1__6__1_,
         U1_level_node_1__6__2_, U1_level_node_1__7__0_,
         U1_level_node_1__7__1_, U1_level_node_1__8__0_,
         U1_level_node_2__3__0_, U1_level_node_2__4__0_,
         U1_level_node_2__4__1_, U1_level_node_2__5__0_,
         U1_level_node_2__5__1_, U1_level_node_2__6__0_,
         U1_level_node_2__6__1_, U1_level_node_2__7__0_,
         U1_level_node_2__7__1_, U1_level_node_2__8__0_,
         U1_level_node_2__8__1_, U1_level_node_2__9__0_,
         U1_level_node_3__2__0_, U1_level_node_3__3__0_,
         U1_level_node_3__3__1_, U1_level_node_3__4__0_,
         U1_level_node_3__4__1_, U1_level_node_3__5__0_,
         U1_level_node_3__5__1_, U1_level_node_3__6__0_,
         U1_level_node_3__6__1_, U1_level_node_3__7__0_,
         U1_level_node_3__7__1_, U1_level_node_3__8__0_,
         U1_level_node_3__8__1_, U1_level_node_3__9__0_,
         U1_level_node_3__9__1_, U1_level_node_3__10__0_,
         U1_B_neg_correction_1_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303;

  nor02 U5 ( .Y(n1), .A0(n294), .A1(n295) );
  inv04 U6 ( .Y(n294), .A(A[3]) );
  or02 U7 ( .Y(n2), .A0(n298), .A1(n301) );
  inv01 U8 ( .Y(n3), .A(n2) );
  or02 U9 ( .Y(n4), .A0(n297), .A1(n300) );
  inv01 U10 ( .Y(n5), .A(n4) );
  or02 U11 ( .Y(n6), .A0(n299), .A1(n300) );
  inv01 U12 ( .Y(n7), .A(n6) );
  or02 U13 ( .Y(n8), .A0(n302), .A1(n303) );
  inv01 U14 ( .Y(n9), .A(n8) );
  or02 U15 ( .Y(n10), .A0(n292), .A1(n301) );
  inv01 U16 ( .Y(n11), .A(n10) );
  or02 U17 ( .Y(n12), .A0(n294), .A1(n301) );
  inv01 U18 ( .Y(n13), .A(n12) );
  or02 U19 ( .Y(n14), .A0(n296), .A1(n301) );
  inv01 U20 ( .Y(n15), .A(n14) );
  or02 U21 ( .Y(n16), .A0(n296), .A1(n299) );
  inv02 U22 ( .Y(n17), .A(n16) );
  or02 U23 ( .Y(n18), .A0(n298), .A1(n299) );
  inv02 U24 ( .Y(n19), .A(n18) );
  or02 U25 ( .Y(n20), .A0(n294), .A1(n299) );
  inv02 U26 ( .Y(n21), .A(n20) );
  nand02 U27 ( .Y(n22), .A0(n51), .A1(n45) );
  inv02 U28 ( .Y(n23), .A(n22) );
  nand02 U29 ( .Y(n24), .A0(n49), .A1(n47) );
  inv02 U30 ( .Y(n25), .A(n24) );
  inv01 U31 ( .Y(n26), .A(n118) );
  inv01 U32 ( .Y(n27), .A(n174) );
  inv01 U33 ( .Y(n28), .A(n176) );
  inv01 U34 ( .Y(n29), .A(n93) );
  or02 U35 ( .Y(n30), .A0(n293), .A1(n302) );
  inv02 U36 ( .Y(n31), .A(n30) );
  or02 U37 ( .Y(n32), .A0(n297), .A1(n302) );
  inv02 U38 ( .Y(n33), .A(n32) );
  or02 U39 ( .Y(n34), .A0(n301), .A1(n302) );
  inv02 U40 ( .Y(n35), .A(n34) );
  or02 U41 ( .Y(n36), .A0(n293), .A1(n300) );
  inv02 U42 ( .Y(n37), .A(n36) );
  or02 U43 ( .Y(n38), .A0(n295), .A1(n300) );
  inv02 U44 ( .Y(n39), .A(n38) );
  or02 U45 ( .Y(n40), .A0(n295), .A1(n302) );
  inv02 U46 ( .Y(n41), .A(n40) );
  buf02 U47 ( .Y(n42), .A(U1_level_node_2__4__1_) );
  buf02 U48 ( .Y(n43), .A(U1_level_node_2__3__0_) );
  buf02 U49 ( .Y(n44), .A(U1_level_node_0__5__3_) );
  buf02 U50 ( .Y(n45), .A(U1_level_node_0__5__3_) );
  buf02 U51 ( .Y(n46), .A(U1_B_neg_correction_1_) );
  buf02 U52 ( .Y(n47), .A(U1_B_neg_correction_1_) );
  or02 U53 ( .Y(n48), .A0(n299), .A1(n302) );
  inv02 U54 ( .Y(n49), .A(n48) );
  or02 U55 ( .Y(n50), .A0(n300), .A1(n303) );
  inv02 U56 ( .Y(n51), .A(n50) );
  or02 U57 ( .Y(n52), .A0(n297), .A1(n298) );
  inv02 U58 ( .Y(n53), .A(n52) );
  or02 U59 ( .Y(n54), .A0(n294), .A1(n303) );
  inv02 U60 ( .Y(n55), .A(n54) );
  or02 U61 ( .Y(n56), .A0(n292), .A1(n293) );
  inv02 U62 ( .Y(n57), .A(n56) );
  inv02 U63 ( .Y(U1_level_node_2__8__0_), .A(n58) );
  inv02 U64 ( .Y(U1_level_node_2__9__0_), .A(n59) );
  inv02 U65 ( .Y(n60), .A(n57) );
  inv02 U66 ( .Y(n61), .A(U1_level_node_1__8__0_) );
  inv02 U67 ( .Y(n62), .A(n55) );
  nor02 U68 ( .Y(n63), .A0(n60), .A1(n64) );
  nor02 U69 ( .Y(n65), .A0(n61), .A1(n66) );
  nor02 U70 ( .Y(n67), .A0(n62), .A1(n68) );
  nor02 U71 ( .Y(n69), .A0(n62), .A1(n70) );
  nor02 U72 ( .Y(n58), .A0(n71), .A1(n72) );
  nor02 U73 ( .Y(n73), .A0(n61), .A1(n62) );
  nor02 U74 ( .Y(n74), .A0(n60), .A1(n62) );
  nor02 U75 ( .Y(n75), .A0(n60), .A1(n61) );
  nor02 U76 ( .Y(n59), .A0(n75), .A1(n76) );
  nor02 U77 ( .Y(n77), .A0(U1_level_node_1__8__0_), .A1(n55) );
  inv01 U78 ( .Y(n64), .A(n77) );
  nor02 U79 ( .Y(n78), .A0(n57), .A1(n55) );
  inv01 U80 ( .Y(n66), .A(n78) );
  nor02 U81 ( .Y(n79), .A0(n57), .A1(U1_level_node_1__8__0_) );
  inv01 U82 ( .Y(n68), .A(n79) );
  nor02 U83 ( .Y(n80), .A0(n60), .A1(n61) );
  inv01 U84 ( .Y(n70), .A(n80) );
  nor02 U85 ( .Y(n81), .A0(n63), .A1(n65) );
  inv01 U86 ( .Y(n71), .A(n81) );
  nor02 U87 ( .Y(n82), .A0(n67), .A1(n69) );
  inv01 U88 ( .Y(n72), .A(n82) );
  nor02 U89 ( .Y(n83), .A0(n73), .A1(n74) );
  inv01 U90 ( .Y(n76), .A(n83) );
  or02 U91 ( .Y(n84), .A0(n292), .A1(n303) );
  inv02 U92 ( .Y(n85), .A(n84) );
  or02 U93 ( .Y(n86), .A0(n296), .A1(n297) );
  inv02 U94 ( .Y(n87), .A(n86) );
  or02 U95 ( .Y(n88), .A0(n295), .A1(n298) );
  inv02 U96 ( .Y(n89), .A(n88) );
  inv02 U97 ( .Y(U1_level_node_2__4__0_), .A(n90) );
  inv02 U98 ( .Y(U1_level_node_2__5__1_), .A(n91) );
  inv02 U99 ( .Y(n92), .A(n87) );
  inv02 U100 ( .Y(n93), .A(U1_level_node_1__4__0_) );
  inv02 U101 ( .Y(n94), .A(n89) );
  nor02 U102 ( .Y(n95), .A0(n92), .A1(n96) );
  nor02 U103 ( .Y(n97), .A0(n93), .A1(n98) );
  nor02 U104 ( .Y(n99), .A0(n94), .A1(n100) );
  nor02 U105 ( .Y(n101), .A0(n94), .A1(n102) );
  nor02 U106 ( .Y(n90), .A0(n103), .A1(n104) );
  nor02 U107 ( .Y(n105), .A0(n93), .A1(n94) );
  nor02 U108 ( .Y(n106), .A0(n92), .A1(n94) );
  nor02 U109 ( .Y(n107), .A0(n92), .A1(n93) );
  nor02 U110 ( .Y(n91), .A0(n107), .A1(n108) );
  nor02 U111 ( .Y(n109), .A0(U1_level_node_1__4__0_), .A1(n89) );
  inv01 U112 ( .Y(n96), .A(n109) );
  nor02 U113 ( .Y(n110), .A0(n87), .A1(n89) );
  inv01 U114 ( .Y(n98), .A(n110) );
  nor02 U115 ( .Y(n111), .A0(n87), .A1(n29) );
  inv01 U116 ( .Y(n100), .A(n111) );
  nor02 U117 ( .Y(n112), .A0(n92), .A1(n93) );
  inv01 U118 ( .Y(n102), .A(n112) );
  nor02 U119 ( .Y(n113), .A0(n95), .A1(n97) );
  inv01 U120 ( .Y(n103), .A(n113) );
  nor02 U121 ( .Y(n114), .A0(n99), .A1(n101) );
  inv01 U122 ( .Y(n104), .A(n114) );
  nor02 U123 ( .Y(n115), .A0(n105), .A1(n106) );
  inv01 U124 ( .Y(n108), .A(n115) );
  inv02 U125 ( .Y(U1_level_node_2__6__0_), .A(n116) );
  inv02 U126 ( .Y(U1_level_node_2__7__1_), .A(n117) );
  inv02 U127 ( .Y(n118), .A(U1_level_node_1__6__1_) );
  inv02 U128 ( .Y(n119), .A(U1_level_node_1__6__0_) );
  inv02 U129 ( .Y(n120), .A(U1_level_node_1__6__2_) );
  nor02 U130 ( .Y(n121), .A0(n118), .A1(n122) );
  nor02 U131 ( .Y(n123), .A0(n119), .A1(n124) );
  nor02 U132 ( .Y(n125), .A0(n120), .A1(n126) );
  nor02 U133 ( .Y(n127), .A0(n120), .A1(n128) );
  nor02 U134 ( .Y(n116), .A0(n129), .A1(n130) );
  nor02 U135 ( .Y(n131), .A0(n119), .A1(n120) );
  nor02 U136 ( .Y(n132), .A0(n118), .A1(n120) );
  nor02 U137 ( .Y(n133), .A0(n118), .A1(n119) );
  nor02 U138 ( .Y(n117), .A0(n133), .A1(n134) );
  nor02 U139 ( .Y(n135), .A0(U1_level_node_1__6__0_), .A1(
        U1_level_node_1__6__2_) );
  inv01 U140 ( .Y(n122), .A(n135) );
  nor02 U141 ( .Y(n136), .A0(n26), .A1(U1_level_node_1__6__2_) );
  inv01 U142 ( .Y(n124), .A(n136) );
  nor02 U143 ( .Y(n137), .A0(U1_level_node_1__6__1_), .A1(
        U1_level_node_1__6__0_) );
  inv01 U144 ( .Y(n126), .A(n137) );
  nor02 U145 ( .Y(n138), .A0(n118), .A1(n119) );
  inv01 U146 ( .Y(n128), .A(n138) );
  nor02 U147 ( .Y(n139), .A0(n121), .A1(n123) );
  inv01 U148 ( .Y(n129), .A(n139) );
  nor02 U149 ( .Y(n140), .A0(n125), .A1(n127) );
  inv01 U150 ( .Y(n130), .A(n140) );
  nor02 U151 ( .Y(n141), .A0(n131), .A1(n132) );
  inv01 U152 ( .Y(n134), .A(n141) );
  or02 U153 ( .Y(n142), .A0(n295), .A1(n296) );
  inv02 U154 ( .Y(n143), .A(n142) );
  or02 U155 ( .Y(n144), .A0(n294), .A1(n297) );
  inv02 U156 ( .Y(n145), .A(n144) );
  inv02 U157 ( .Y(U1_level_node_1__5__0_), .A(n146) );
  inv02 U158 ( .Y(U1_level_node_1__6__2_), .A(n147) );
  inv02 U159 ( .Y(n148), .A(n145) );
  inv02 U160 ( .Y(n149), .A(n288) );
  inv02 U161 ( .Y(n150), .A(n143) );
  nor02 U162 ( .Y(n151), .A0(n148), .A1(n152) );
  nor02 U163 ( .Y(n153), .A0(n149), .A1(n154) );
  nor02 U164 ( .Y(n155), .A0(n150), .A1(n156) );
  nor02 U165 ( .Y(n157), .A0(n150), .A1(n158) );
  nor02 U166 ( .Y(n146), .A0(n159), .A1(n160) );
  nor02 U167 ( .Y(n161), .A0(n149), .A1(n150) );
  nor02 U168 ( .Y(n162), .A0(n148), .A1(n150) );
  nor02 U169 ( .Y(n163), .A0(n148), .A1(n149) );
  nor02 U170 ( .Y(n147), .A0(n163), .A1(n164) );
  nor02 U171 ( .Y(n165), .A0(n288), .A1(n143) );
  inv01 U172 ( .Y(n152), .A(n165) );
  nor02 U173 ( .Y(n166), .A0(n145), .A1(n143) );
  inv01 U174 ( .Y(n154), .A(n166) );
  nor02 U175 ( .Y(n167), .A0(n145), .A1(n288) );
  inv01 U176 ( .Y(n156), .A(n167) );
  nor02 U177 ( .Y(n168), .A0(n148), .A1(n149) );
  inv01 U178 ( .Y(n158), .A(n168) );
  nor02 U179 ( .Y(n169), .A0(n151), .A1(n153) );
  inv01 U180 ( .Y(n159), .A(n169) );
  nor02 U181 ( .Y(n170), .A0(n155), .A1(n157) );
  inv01 U182 ( .Y(n160), .A(n170) );
  nor02 U183 ( .Y(n171), .A0(n161), .A1(n162) );
  inv01 U184 ( .Y(n164), .A(n171) );
  inv02 U185 ( .Y(U1_level_node_2__5__0_), .A(n172) );
  inv02 U186 ( .Y(U1_level_node_2__6__1_), .A(n173) );
  inv02 U187 ( .Y(n174), .A(U1_level_node_1__5__1_) );
  inv02 U188 ( .Y(n175), .A(U1_level_node_1__5__0_) );
  inv02 U189 ( .Y(n176), .A(U1_level_node_1__5__2_) );
  nor02 U190 ( .Y(n177), .A0(n174), .A1(n178) );
  nor02 U191 ( .Y(n179), .A0(n175), .A1(n180) );
  nor02 U192 ( .Y(n181), .A0(n176), .A1(n182) );
  nor02 U193 ( .Y(n183), .A0(n176), .A1(n184) );
  nor02 U194 ( .Y(n172), .A0(n185), .A1(n186) );
  nor02 U195 ( .Y(n187), .A0(n175), .A1(n176) );
  nor02 U196 ( .Y(n188), .A0(n174), .A1(n176) );
  nor02 U197 ( .Y(n189), .A0(n174), .A1(n175) );
  nor02 U198 ( .Y(n173), .A0(n189), .A1(n190) );
  nor02 U199 ( .Y(n191), .A0(U1_level_node_1__5__0_), .A1(
        U1_level_node_1__5__2_) );
  inv01 U200 ( .Y(n178), .A(n191) );
  nor02 U201 ( .Y(n192), .A0(n27), .A1(n28) );
  inv01 U202 ( .Y(n180), .A(n192) );
  nor02 U203 ( .Y(n193), .A0(U1_level_node_1__5__1_), .A1(
        U1_level_node_1__5__0_) );
  inv01 U204 ( .Y(n182), .A(n193) );
  nor02 U205 ( .Y(n194), .A0(n174), .A1(n175) );
  inv01 U206 ( .Y(n184), .A(n194) );
  nor02 U207 ( .Y(n195), .A0(n177), .A1(n179) );
  inv01 U208 ( .Y(n185), .A(n195) );
  nor02 U209 ( .Y(n196), .A0(n181), .A1(n183) );
  inv01 U210 ( .Y(n186), .A(n196) );
  nor02 U211 ( .Y(n197), .A0(n187), .A1(n188) );
  inv01 U212 ( .Y(n190), .A(n197) );
  or02 U213 ( .Y(n198), .A0(n293), .A1(n296) );
  inv02 U214 ( .Y(n199), .A(n198) );
  or02 U215 ( .Y(n200), .A0(n296), .A1(n303) );
  inv02 U216 ( .Y(n201), .A(n200) );
  nor02 U217 ( .Y(n202), .A0(n294), .A1(n295) );
  or02 U218 ( .Y(n203), .A0(n293), .A1(n294) );
  inv02 U219 ( .Y(n204), .A(n203) );
  inv04 U220 ( .Y(n295), .A(B[3]) );
  inv02 U221 ( .Y(U1_level_node_1__7__0_), .A(n205) );
  inv02 U222 ( .Y(U1_level_node_1__8__0_), .A(n206) );
  inv02 U223 ( .Y(n207), .A(n204) );
  inv02 U224 ( .Y(n208), .A(n286) );
  inv02 U225 ( .Y(n209), .A(n201) );
  nor02 U226 ( .Y(n210), .A0(n207), .A1(n211) );
  nor02 U227 ( .Y(n212), .A0(n208), .A1(n213) );
  nor02 U228 ( .Y(n214), .A0(n209), .A1(n215) );
  nor02 U229 ( .Y(n216), .A0(n209), .A1(n217) );
  nor02 U230 ( .Y(n205), .A0(n218), .A1(n219) );
  nor02 U231 ( .Y(n220), .A0(n208), .A1(n209) );
  nor02 U232 ( .Y(n221), .A0(n207), .A1(n209) );
  nor02 U233 ( .Y(n222), .A0(n207), .A1(n208) );
  nor02 U234 ( .Y(n206), .A0(n222), .A1(n223) );
  nor02 U235 ( .Y(n224), .A0(n286), .A1(n201) );
  inv01 U236 ( .Y(n211), .A(n224) );
  nor02 U237 ( .Y(n225), .A0(n204), .A1(n201) );
  inv01 U238 ( .Y(n213), .A(n225) );
  nor02 U239 ( .Y(n226), .A0(n204), .A1(n286) );
  inv01 U240 ( .Y(n215), .A(n226) );
  nor02 U241 ( .Y(n227), .A0(n207), .A1(n208) );
  inv01 U242 ( .Y(n217), .A(n227) );
  nor02 U243 ( .Y(n228), .A0(n210), .A1(n212) );
  inv01 U244 ( .Y(n218), .A(n228) );
  nor02 U245 ( .Y(n229), .A0(n214), .A1(n216) );
  inv01 U246 ( .Y(n219), .A(n229) );
  nor02 U247 ( .Y(n230), .A0(n220), .A1(n221) );
  inv01 U248 ( .Y(n223), .A(n230) );
  inv02 U249 ( .Y(U1_level_node_1__6__0_), .A(n231) );
  inv02 U250 ( .Y(U1_level_node_1__7__1_), .A(n232) );
  inv02 U251 ( .Y(n233), .A(U1_level_node_0__6__1_) );
  inv02 U252 ( .Y(n234), .A(n284) );
  inv02 U253 ( .Y(n235), .A(n199) );
  nor02 U254 ( .Y(n236), .A0(n233), .A1(n237) );
  nor02 U255 ( .Y(n238), .A0(n234), .A1(n239) );
  nor02 U256 ( .Y(n240), .A0(n235), .A1(n241) );
  nor02 U257 ( .Y(n242), .A0(n235), .A1(n243) );
  nor02 U258 ( .Y(n231), .A0(n244), .A1(n245) );
  nor02 U259 ( .Y(n246), .A0(n234), .A1(n235) );
  nor02 U260 ( .Y(n247), .A0(n233), .A1(n235) );
  nor02 U261 ( .Y(n248), .A0(n233), .A1(n234) );
  nor02 U262 ( .Y(n232), .A0(n248), .A1(n249) );
  nor02 U263 ( .Y(n250), .A0(n284), .A1(n199) );
  inv01 U264 ( .Y(n237), .A(n250) );
  nor02 U265 ( .Y(n251), .A0(n202), .A1(n199) );
  inv01 U266 ( .Y(n239), .A(n251) );
  nor02 U267 ( .Y(n252), .A0(n1), .A1(n284) );
  inv01 U268 ( .Y(n241), .A(n252) );
  nor02 U269 ( .Y(n253), .A0(n233), .A1(n234) );
  inv01 U270 ( .Y(n243), .A(n253) );
  nor02 U271 ( .Y(n254), .A0(n236), .A1(n238) );
  inv01 U272 ( .Y(n244), .A(n254) );
  nor02 U273 ( .Y(n255), .A0(n240), .A1(n242) );
  inv01 U274 ( .Y(n245), .A(n255) );
  nor02 U275 ( .Y(n256), .A0(n246), .A1(n247) );
  inv01 U276 ( .Y(n249), .A(n256) );
  inv02 U277 ( .Y(U1_level_node_2__7__0_), .A(n257) );
  inv02 U278 ( .Y(U1_level_node_2__8__1_), .A(n258) );
  inv02 U279 ( .Y(n259), .A(U1_level_node_1__7__1_) );
  inv02 U280 ( .Y(n260), .A(U1_level_node_1__7__0_) );
  inv02 U281 ( .Y(n261), .A(n25) );
  nor02 U282 ( .Y(n262), .A0(n259), .A1(n263) );
  nor02 U283 ( .Y(n264), .A0(n260), .A1(n265) );
  nor02 U284 ( .Y(n266), .A0(n261), .A1(n267) );
  nor02 U285 ( .Y(n268), .A0(n261), .A1(n269) );
  nor02 U286 ( .Y(n257), .A0(n270), .A1(n271) );
  nor02 U287 ( .Y(n272), .A0(n260), .A1(n261) );
  nor02 U288 ( .Y(n273), .A0(n259), .A1(n261) );
  nor02 U289 ( .Y(n274), .A0(n259), .A1(n260) );
  nor02 U290 ( .Y(n258), .A0(n274), .A1(n275) );
  nor02 U291 ( .Y(n276), .A0(U1_level_node_1__7__0_), .A1(n25) );
  inv01 U292 ( .Y(n263), .A(n276) );
  nor02 U293 ( .Y(n277), .A0(U1_level_node_1__7__1_), .A1(n25) );
  inv01 U294 ( .Y(n265), .A(n277) );
  nor02 U295 ( .Y(n278), .A0(U1_level_node_1__7__1_), .A1(
        U1_level_node_1__7__0_) );
  inv01 U296 ( .Y(n267), .A(n278) );
  nor02 U297 ( .Y(n279), .A0(n259), .A1(n260) );
  inv01 U298 ( .Y(n269), .A(n279) );
  nor02 U299 ( .Y(n280), .A0(n262), .A1(n264) );
  inv01 U300 ( .Y(n270), .A(n280) );
  nor02 U301 ( .Y(n281), .A0(n266), .A1(n268) );
  inv01 U302 ( .Y(n271), .A(n281) );
  nor02 U303 ( .Y(n282), .A0(n272), .A1(n273) );
  inv01 U304 ( .Y(n275), .A(n282) );
  or02 U305 ( .Y(n283), .A0(n292), .A1(n297) );
  inv02 U306 ( .Y(n284), .A(n283) );
  or02 U307 ( .Y(n285), .A0(n292), .A1(n295) );
  inv02 U308 ( .Y(n286), .A(n285) );
  or02 U309 ( .Y(n287), .A0(n292), .A1(n299) );
  inv02 U310 ( .Y(n288), .A(n287) );
  or02 U311 ( .Y(n289), .A0(n300), .A1(n301) );
  inv02 U312 ( .Y(PRODUCT[0]), .A(n289) );
  inv02 U313 ( .Y(n293), .A(B[4]) );
  inv02 U314 ( .Y(n299), .A(B[1]) );
  inv02 U315 ( .Y(n298), .A(A[1]) );
  inv02 U316 ( .Y(n297), .A(B[2]) );
  inv02 U317 ( .Y(n301), .A(B[0]) );
  inv02 U318 ( .Y(n303), .A(B[5]) );
  inv02 U319 ( .Y(n292), .A(A[4]) );
  inv02 U320 ( .Y(n296), .A(A[2]) );
  inv02 U321 ( .Y(n300), .A(A[0]) );
  inv02 U322 ( .Y(n302), .A(A[5]) );
  xor2 U323 ( .Y(U1_level_node_1__5__1_), .A0(n44), .A1(n51) );
  xor2 U324 ( .Y(U1_level_node_1__6__1_), .A0(n46), .A1(n49) );
  mul_24_DW01_add_11_1 U1_U9720 ( .A({1'b0, U1_level_node_3__10__0_, 
        U1_level_node_3__9__0_, U1_level_node_3__8__0_, U1_level_node_3__7__0_, 
        U1_level_node_3__6__0_, U1_level_node_3__5__0_, U1_level_node_3__4__0_, 
        U1_level_node_3__3__0_, U1_level_node_3__2__0_, n3}), .B({1'b0, n9, 
        U1_level_node_3__9__1_, U1_level_node_3__8__1_, U1_level_node_3__7__1_, 
        U1_level_node_3__6__1_, U1_level_node_3__5__1_, U1_level_node_3__4__1_, 
        U1_level_node_3__3__1_, n5, n7}), .CI(1'b0), .SUM(PRODUCT[11:1]) );
  nor02 U325 ( .Y(U1_level_node_0__6__1_), .A0(n294), .A1(n295) );
  nor02 U326 ( .Y(U1_level_node_0__5__3_), .A0(n293), .A1(n298) );
  nor02 U327 ( .Y(U1_B_neg_correction_1_), .A0(n298), .A1(n303) );
  hadd1 U1_U3220_1_4 ( .S(U1_level_node_1__4__0_), .CO(U1_level_node_1__5__2_), 
        .A(n11), .B(n21) );
  hadd1 U1_U3220_2_3 ( .S(U1_level_node_2__3__0_), .CO(U1_level_node_2__4__1_), 
        .A(n13), .B(n17) );
  fadd1 U1_U3140_3_9_0 ( .S(U1_level_node_3__9__0_), .CO(
        U1_level_node_3__10__0_), .A(U1_level_node_2__9__0_), .B(n85), .CI(n31) );
  fadd1 U1_U3140_3_8_0 ( .S(U1_level_node_3__8__0_), .CO(
        U1_level_node_3__9__1_), .A(U1_level_node_2__8__0_), .B(
        U1_level_node_2__8__1_), .CI(n41) );
  fadd1 U1_U3140_3_7_0 ( .S(U1_level_node_3__7__0_), .CO(
        U1_level_node_3__8__1_), .A(U1_level_node_2__7__0_), .B(
        U1_level_node_2__7__1_), .CI(n33) );
  fadd1 U1_U3140_3_6_0 ( .S(U1_level_node_3__6__0_), .CO(
        U1_level_node_3__7__1_), .A(U1_level_node_2__6__0_), .B(
        U1_level_node_2__6__1_), .CI(n23) );
  fadd1 U1_U3140_3_5_0 ( .S(U1_level_node_3__5__0_), .CO(
        U1_level_node_3__6__1_), .A(U1_level_node_2__5__0_), .B(
        U1_level_node_2__5__1_), .CI(n35) );
  fadd1 U1_U3140_3_4_0 ( .S(U1_level_node_3__4__0_), .CO(
        U1_level_node_3__5__1_), .A(U1_level_node_2__4__0_), .B(n42), .CI(n37)
         );
  fadd1 U1_U3140_3_3_0 ( .S(U1_level_node_3__3__0_), .CO(
        U1_level_node_3__4__1_), .A(n43), .B(n53), .CI(n39) );
  hadd1 U1_U3220_3_2 ( .S(U1_level_node_3__2__0_), .CO(U1_level_node_3__3__1_), 
        .A(n15), .B(n19) );
endmodule


module mul_24_DW01_add_11_0 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   g_array_0__9_, g_array_0__8_, g_array_0__7_, g_array_0__6_,
         g_array_0__5_, g_array_0__4_, g_array_0__3_, g_array_0__2_,
         g_array_0__1_, g_array_0__0_, g_array_1__9_, g_array_1__8_,
         g_array_1__7_, g_array_1__6_, g_array_1__5_, g_array_1__4_,
         g_array_1__3_, g_array_1__2_, g_array_1__1_, g_array_1__0_,
         g_array_2__9_, g_array_2__8_, g_array_2__7_, g_array_2__6_,
         g_array_2__5_, g_array_2__4_, g_array_2__3_, g_array_2__2_,
         g_array_2__1_, g_array_2__0_, g_array_3__9_, g_array_3__8_,
         g_array_3__7_, g_array_3__6_, g_array_3__5_, g_array_3__4_,
         g_array_3__3_, g_array_3__2_, g_array_3__1_, g_array_3__0_,
         g_array_4__9_, g_array_4__6_, g_array_4__5_, g_array_4__3_,
         g_array_4__2_, g_array_4__1_, g_array_4__0_, pog_array_0__9_,
         pog_array_0__0_, pog_array_1__9_, pog_array_1__8_, pog_array_1__7_,
         pog_array_1__6_, pog_array_1__5_, pog_array_1__3_, pog_array_1__2_,
         pog_array_1__1_, pog_array_2__9_, pog_array_2__8_, pog_array_2__7_,
         pog_array_2__6_, pog_array_2__5_, pog_array_2__4_, pog_array_2__3_,
         pog_array_2__1_, pog_array_3__9_, pog_array_3__8_, pog_array_3__7_,
         pog_array_3__5_, pog_array_3__4_, pog_array_3__3_, part_sum_9_,
         part_sum_8_, part_sum_7_, part_sum_6_, part_sum_5_, part_sum_4_,
         part_sum_3_, part_sum_2_, part_sum_1_, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n87, n89, n91, n93, n95, n97, n99,
         n101, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134;

  inv02 U1_2_0_5 ( .Y(g_array_1__5_), .A(g_array_0__5_) );
  inv02 U1_2_0_7 ( .Y(g_array_1__7_), .A(g_array_0__7_) );
  inv02 U7 ( .Y(part_sum_5_), .A(n124) );
  inv02 U8 ( .Y(part_sum_7_), .A(n122) );
  inv01 U9 ( .Y(g_array_3__9_), .A(n31) );
  nor02 U10 ( .Y(n32), .A0(pog_array_2__9_), .A1(g_array_2__8_) );
  inv01 U11 ( .Y(n33), .A(g_array_2__9_) );
  nor02 U12 ( .Y(n31), .A0(n32), .A1(n33) );
  inv01 U13 ( .Y(g_array_3__5_), .A(n34) );
  nor02 U14 ( .Y(n35), .A0(pog_array_2__5_), .A1(g_array_2__4_) );
  inv01 U15 ( .Y(n36), .A(g_array_2__5_) );
  nor02 U16 ( .Y(n34), .A0(n35), .A1(n36) );
  inv02 U1_3_1_9 ( .Y(pog_array_2__9_), .A(pog_array_1__9_) );
  inv02 U1_2_1_9 ( .Y(g_array_2__9_), .A(g_array_1__9_) );
  inv02 U1_3_1_5 ( .Y(pog_array_2__5_), .A(pog_array_1__5_) );
  inv02 U1_2_1_5 ( .Y(g_array_2__5_), .A(g_array_1__5_) );
  inv01 U17 ( .Y(g_array_1__2_), .A(n37) );
  nor02 U18 ( .Y(n38), .A0(n109), .A1(g_array_0__1_) );
  inv01 U19 ( .Y(n39), .A(g_array_0__2_) );
  nor02 U20 ( .Y(n37), .A0(n38), .A1(n39) );
  nand02 U21 ( .Y(g_array_1__6_), .A0(n40), .A1(g_array_0__6_) );
  inv01 U22 ( .Y(n41), .A(g_array_0__5_) );
  inv01 U23 ( .Y(n42), .A(n115) );
  nand02 U24 ( .Y(n40), .A0(n41), .A1(n42) );
  nand02 U25 ( .Y(g_array_4__9_), .A0(n43), .A1(n44) );
  inv01 U26 ( .Y(n45), .A(g_array_3__9_) );
  inv01 U27 ( .Y(n46), .A(g_array_3__6_) );
  inv01 U28 ( .Y(n47), .A(pog_array_3__9_) );
  nand02 U29 ( .Y(n43), .A0(n45), .A1(n46) );
  nand02 U30 ( .Y(n44), .A0(n45), .A1(n47) );
  inv02 U1_2_0_9 ( .Y(g_array_1__9_), .A(g_array_0__9_) );
  inv02 U1_3_1_8 ( .Y(pog_array_2__8_), .A(pog_array_1__8_) );
  inv02 U1_3_0_9 ( .Y(pog_array_1__9_), .A(pog_array_0__9_) );
  inv02 U31 ( .Y(g_array_3__1_), .A(n48) );
  nor02 U32 ( .Y(n49), .A0(pog_array_2__1_), .A1(g_array_2__0_) );
  inv01 U33 ( .Y(n50), .A(g_array_2__1_) );
  nor02 U34 ( .Y(n48), .A0(n49), .A1(n50) );
  inv02 U1_3_1_1 ( .Y(pog_array_2__1_), .A(pog_array_1__1_) );
  inv02 U1_2_1_0 ( .Y(g_array_2__0_), .A(g_array_1__0_) );
  inv02 U1_2_1_1 ( .Y(g_array_2__1_), .A(g_array_1__1_) );
  inv02 U35 ( .Y(n130), .A(pog_array_0__0_) );
  nand02 U36 ( .Y(g_array_1__8_), .A0(n51), .A1(g_array_0__8_) );
  inv01 U37 ( .Y(n52), .A(g_array_0__7_) );
  inv01 U38 ( .Y(n53), .A(n113) );
  nand02 U39 ( .Y(n51), .A0(n52), .A1(n53) );
  inv02 U1_2_1_8 ( .Y(g_array_2__8_), .A(g_array_1__8_) );
  nand02 U40 ( .Y(g_array_4__3_), .A0(n54), .A1(n55) );
  inv01 U41 ( .Y(n56), .A(g_array_3__3_) );
  inv01 U42 ( .Y(n57), .A(g_array_3__2_) );
  inv01 U43 ( .Y(n58), .A(pog_array_3__3_) );
  nand02 U44 ( .Y(n54), .A0(n56), .A1(n57) );
  nand02 U45 ( .Y(n55), .A0(n56), .A1(n58) );
  ao21 U46 ( .Y(n59), .A0(pog_array_3__4_), .A1(g_array_3__2_), .B0(
        g_array_3__4_) );
  inv01 U47 ( .Y(n60), .A(n59) );
  inv02 U48 ( .Y(SUM[10]), .A(g_array_4__9_) );
  inv02 U1_3_2_3 ( .Y(pog_array_3__3_), .A(pog_array_2__3_) );
  inv02 U1_2_2_3 ( .Y(g_array_3__3_), .A(g_array_2__3_) );
  nand02 U49 ( .Y(g_array_4__5_), .A0(n61), .A1(n62) );
  inv01 U50 ( .Y(n63), .A(g_array_3__5_) );
  inv01 U51 ( .Y(n64), .A(g_array_3__2_) );
  inv01 U52 ( .Y(n65), .A(pog_array_3__5_) );
  nand02 U53 ( .Y(n61), .A0(n63), .A1(n64) );
  nand02 U54 ( .Y(n62), .A0(n63), .A1(n65) );
  ao21 U55 ( .Y(n66), .A0(pog_array_3__7_), .A1(g_array_3__6_), .B0(
        g_array_3__7_) );
  inv01 U56 ( .Y(n67), .A(n66) );
  ao21 U57 ( .Y(n68), .A0(pog_array_3__8_), .A1(g_array_3__6_), .B0(
        g_array_3__8_) );
  inv01 U58 ( .Y(n69), .A(n68) );
  inv02 U1_2_0_3 ( .Y(g_array_1__3_), .A(g_array_0__3_) );
  inv01 U1_2_0_1 ( .Y(g_array_1__1_), .A(g_array_0__1_) );
  nand02 U59 ( .Y(g_array_1__4_), .A0(n70), .A1(g_array_0__4_) );
  inv01 U60 ( .Y(n71), .A(g_array_0__3_) );
  inv01 U61 ( .Y(n72), .A(n111) );
  nand02 U62 ( .Y(n70), .A0(n71), .A1(n72) );
  inv02 U1_2_1_4 ( .Y(g_array_2__4_), .A(g_array_1__4_) );
  or02 U63 ( .Y(n73), .A0(A[5]), .A1(B[5]) );
  inv01 U64 ( .Y(n74), .A(n73) );
  inv01 U65 ( .Y(n75), .A(n73) );
  or02 U66 ( .Y(n76), .A0(A[3]), .A1(B[3]) );
  inv01 U67 ( .Y(n77), .A(n76) );
  inv02 U1_3_0_5 ( .Y(pog_array_1__5_), .A(n74) );
  inv02 U1_3_0_3 ( .Y(pog_array_1__3_), .A(n77) );
  or02 U68 ( .Y(n78), .A0(A[7]), .A1(B[7]) );
  inv01 U69 ( .Y(n79), .A(n78) );
  inv01 U70 ( .Y(n80), .A(n78) );
  inv02 U1_3_0_7 ( .Y(pog_array_1__7_), .A(n79) );
  or02 U71 ( .Y(n81), .A0(A[1]), .A1(B[1]) );
  inv01 U72 ( .Y(n82), .A(n81) );
  inv02 U1_3_0_1 ( .Y(pog_array_1__1_), .A(n82) );
  or02 U73 ( .Y(n83), .A0(n77), .A1(n111) );
  inv01 U74 ( .Y(n84), .A(n83) );
  inv02 U1_3_1_4 ( .Y(pog_array_2__4_), .A(n84) );
  xor2 U75 ( .Y(n85), .A0(part_sum_4_), .A1(g_array_4__3_) );
  inv02 U76 ( .Y(SUM[4]), .A(n85) );
  xor2 U77 ( .Y(n87), .A0(part_sum_8_), .A1(n67) );
  inv02 U78 ( .Y(SUM[8]), .A(n87) );
  xor2 U79 ( .Y(n89), .A0(part_sum_6_), .A1(g_array_4__5_) );
  inv02 U80 ( .Y(SUM[6]), .A(n89) );
  xor2 U81 ( .Y(n91), .A0(part_sum_9_), .A1(n69) );
  inv02 U82 ( .Y(SUM[9]), .A(n91) );
  xor2 U83 ( .Y(n93), .A0(part_sum_2_), .A1(g_array_4__1_) );
  inv02 U84 ( .Y(SUM[2]), .A(n93) );
  xor2 U85 ( .Y(n95), .A0(part_sum_3_), .A1(g_array_4__2_) );
  inv02 U86 ( .Y(SUM[3]), .A(n95) );
  xor2 U87 ( .Y(n97), .A0(part_sum_5_), .A1(n60) );
  inv02 U88 ( .Y(SUM[5]), .A(n97) );
  xor2 U89 ( .Y(n99), .A0(part_sum_7_), .A1(g_array_4__6_) );
  inv02 U90 ( .Y(SUM[7]), .A(n99) );
  xor2 U91 ( .Y(n101), .A0(part_sum_1_), .A1(g_array_4__0_) );
  inv02 U92 ( .Y(SUM[1]), .A(n101) );
  nand02 U93 ( .Y(g_array_2__2_), .A0(n103), .A1(n104) );
  inv01 U94 ( .Y(n105), .A(g_array_1__2_) );
  inv01 U95 ( .Y(n106), .A(g_array_1__0_) );
  inv01 U96 ( .Y(n107), .A(pog_array_1__2_) );
  nand02 U97 ( .Y(n103), .A0(n105), .A1(n106) );
  nand02 U98 ( .Y(n104), .A0(n105), .A1(n107) );
  inv02 U1_2_2_2 ( .Y(g_array_3__2_), .A(g_array_2__2_) );
  inv02 U99 ( .Y(g_array_1__0_), .A(g_array_0__0_) );
  or02 U100 ( .Y(n108), .A0(A[2]), .A1(B[2]) );
  inv02 U101 ( .Y(n109), .A(n108) );
  inv01 U102 ( .Y(n131), .A(n109) );
  or02 U103 ( .Y(n110), .A0(A[4]), .A1(B[4]) );
  inv02 U104 ( .Y(n111), .A(n110) );
  or02 U105 ( .Y(n112), .A0(A[8]), .A1(B[8]) );
  inv02 U106 ( .Y(n113), .A(n112) );
  inv01 U107 ( .Y(n132), .A(n111) );
  inv01 U108 ( .Y(n134), .A(n113) );
  or02 U109 ( .Y(n114), .A0(A[6]), .A1(B[6]) );
  inv01 U110 ( .Y(n115), .A(n114) );
  inv01 U111 ( .Y(n116), .A(n114) );
  inv01 U112 ( .Y(n133), .A(n115) );
  inv02 U113 ( .Y(g_array_3__6_), .A(n117) );
  nor02 U114 ( .Y(n118), .A0(pog_array_2__6_), .A1(g_array_2__2_) );
  inv01 U115 ( .Y(n119), .A(g_array_2__6_) );
  nor02 U116 ( .Y(n117), .A0(n118), .A1(n119) );
  inv04 U117 ( .Y(part_sum_9_), .A(n120) );
  inv04 U118 ( .Y(part_sum_8_), .A(n121) );
  inv04 U119 ( .Y(part_sum_6_), .A(n123) );
  inv04 U120 ( .Y(part_sum_4_), .A(n125) );
  inv04 U121 ( .Y(part_sum_3_), .A(n126) );
  inv04 U122 ( .Y(part_sum_2_), .A(n127) );
  inv04 U123 ( .Y(part_sum_1_), .A(n128) );
  inv04 U124 ( .Y(SUM[0]), .A(n129) );
  nand02 U0_1_0 ( .Y(g_array_0__0_), .A0(A[0]), .A1(B[0]) );
  nor02 U0_2_0 ( .Y(pog_array_0__0_), .A0(A[0]), .A1(B[0]) );
  nand02 U0_3_0 ( .Y(n129), .A0(g_array_0__0_), .A1(n130) );
  nand02 U0_1_1 ( .Y(g_array_0__1_), .A0(A[1]), .A1(B[1]) );
  nand02 U0_3_1 ( .Y(n128), .A0(g_array_0__1_), .A1(pog_array_1__1_) );
  nand02 U0_1_2 ( .Y(g_array_0__2_), .A0(A[2]), .A1(B[2]) );
  nand02 U0_3_2 ( .Y(n127), .A0(g_array_0__2_), .A1(n131) );
  nand02 U0_1_3 ( .Y(g_array_0__3_), .A0(A[3]), .A1(B[3]) );
  nand02 U0_3_3 ( .Y(n126), .A0(g_array_0__3_), .A1(pog_array_1__3_) );
  nand02 U0_1_4 ( .Y(g_array_0__4_), .A0(A[4]), .A1(B[4]) );
  nand02 U0_3_4 ( .Y(n125), .A0(g_array_0__4_), .A1(n132) );
  nand02 U0_1_5 ( .Y(g_array_0__5_), .A0(A[5]), .A1(B[5]) );
  nand02 U0_3_5 ( .Y(n124), .A0(g_array_0__5_), .A1(pog_array_1__5_) );
  nand02 U0_1_6 ( .Y(g_array_0__6_), .A0(A[6]), .A1(B[6]) );
  nand02 U0_3_6 ( .Y(n123), .A0(g_array_0__6_), .A1(n133) );
  nand02 U0_1_7 ( .Y(g_array_0__7_), .A0(A[7]), .A1(B[7]) );
  nand02 U0_3_7 ( .Y(n122), .A0(g_array_0__7_), .A1(pog_array_1__7_) );
  nand02 U0_1_8 ( .Y(g_array_0__8_), .A0(A[8]), .A1(B[8]) );
  nand02 U0_3_8 ( .Y(n121), .A0(g_array_0__8_), .A1(n134) );
  nand02 U0_1_9 ( .Y(g_array_0__9_), .A0(A[9]), .A1(B[9]) );
  nor02 U0_2_9 ( .Y(pog_array_0__9_), .A0(A[9]), .A1(B[9]) );
  nand02 U0_3_9 ( .Y(n120), .A0(g_array_0__9_), .A1(pog_array_1__9_) );
  nor02 U1_5_0_2 ( .Y(pog_array_1__2_), .A0(n82), .A1(n109) );
  nor02 U1_5_0_6 ( .Y(pog_array_1__6_), .A0(n75), .A1(n116) );
  nor02 U1_5_0_8 ( .Y(pog_array_1__8_), .A0(n80), .A1(n113) );
  inv04 U1_2_1_3 ( .Y(g_array_2__3_), .A(g_array_1__3_) );
  inv04 U1_3_1_3 ( .Y(pog_array_2__3_), .A(pog_array_1__3_) );
  aoi21 U1_4_1_6 ( .Y(g_array_2__6_), .A0(pog_array_1__6_), .A1(g_array_1__4_), 
        .B0(g_array_1__6_) );
  nand02 U1_5_1_6 ( .Y(pog_array_2__6_), .A0(pog_array_1__6_), .A1(n84) );
  inv04 U1_2_1_7 ( .Y(g_array_2__7_), .A(g_array_1__7_) );
  inv04 U1_3_1_7 ( .Y(pog_array_2__7_), .A(pog_array_1__7_) );
  inv04 U1_2_2_0 ( .Y(g_array_3__0_), .A(g_array_2__0_) );
  inv04 U1_2_2_4 ( .Y(g_array_3__4_), .A(g_array_2__4_) );
  inv04 U1_3_2_4 ( .Y(pog_array_3__4_), .A(pog_array_2__4_) );
  nor02 U1_5_2_5 ( .Y(pog_array_3__5_), .A0(pog_array_2__4_), .A1(
        pog_array_2__5_) );
  inv04 U1_2_2_7 ( .Y(g_array_3__7_), .A(g_array_2__7_) );
  inv04 U1_3_2_7 ( .Y(pog_array_3__7_), .A(pog_array_2__7_) );
  inv04 U1_2_2_8 ( .Y(g_array_3__8_), .A(g_array_2__8_) );
  inv04 U1_3_2_8 ( .Y(pog_array_3__8_), .A(pog_array_2__8_) );
  nor02 U1_5_2_9 ( .Y(pog_array_3__9_), .A0(pog_array_2__8_), .A1(
        pog_array_2__9_) );
  inv04 U1_2_3_0 ( .Y(g_array_4__0_), .A(g_array_3__0_) );
  inv04 U1_2_3_1 ( .Y(g_array_4__1_), .A(g_array_3__1_) );
  inv04 U1_2_3_2 ( .Y(g_array_4__2_), .A(g_array_3__2_) );
  inv04 U1_2_3_6 ( .Y(g_array_4__6_), .A(g_array_3__6_) );
endmodule


module mul_24_DW02_mult_6_6_0 ( A, B, TC, PRODUCT );
  input [5:0] A;
  input [5:0] B;
  output [11:0] PRODUCT;
  input TC;
  wire   U1_level_node_1__4__0_, U1_level_node_1__5__0_,
         U1_level_node_1__5__1_, U1_level_node_1__5__2_,
         U1_level_node_1__6__0_, U1_level_node_1__6__1_,
         U1_level_node_1__6__2_, U1_level_node_1__7__0_,
         U1_level_node_1__7__1_, U1_level_node_1__8__0_,
         U1_level_node_2__3__0_, U1_level_node_2__4__0_,
         U1_level_node_2__4__1_, U1_level_node_2__5__0_,
         U1_level_node_2__5__1_, U1_level_node_2__6__0_,
         U1_level_node_2__6__1_, U1_level_node_2__7__0_,
         U1_level_node_2__7__1_, U1_level_node_2__8__0_,
         U1_level_node_2__8__1_, U1_level_node_2__9__0_,
         U1_level_node_3__2__0_, U1_level_node_3__3__0_,
         U1_level_node_3__3__1_, U1_level_node_3__4__0_,
         U1_level_node_3__4__1_, U1_level_node_3__5__0_,
         U1_level_node_3__5__1_, U1_level_node_3__6__0_,
         U1_level_node_3__6__1_, U1_level_node_3__7__0_,
         U1_level_node_3__7__1_, U1_level_node_3__8__0_,
         U1_level_node_3__8__1_, U1_level_node_3__9__0_,
         U1_level_node_3__9__1_, U1_level_node_3__10__0_,
         U1_B_neg_correction_2_, U1_B_neg_correction_1_, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303;

  or02 U5 ( .Y(n1), .A0(n298), .A1(n301) );
  inv01 U6 ( .Y(n2), .A(n1) );
  nor02 U7 ( .Y(n3), .A0(n296), .A1(n303) );
  inv04 U8 ( .Y(n296), .A(A[2]) );
  or02 U9 ( .Y(n4), .A0(n297), .A1(n300) );
  inv01 U10 ( .Y(n5), .A(n4) );
  or02 U11 ( .Y(n6), .A0(n299), .A1(n300) );
  inv01 U12 ( .Y(n7), .A(n6) );
  or02 U13 ( .Y(n8), .A0(n302), .A1(n303) );
  inv01 U14 ( .Y(n9), .A(n8) );
  or02 U15 ( .Y(n10), .A0(n296), .A1(n301) );
  inv01 U16 ( .Y(n11), .A(n10) );
  or02 U17 ( .Y(n12), .A0(n292), .A1(n301) );
  inv01 U18 ( .Y(n13), .A(n12) );
  or02 U19 ( .Y(n14), .A0(n294), .A1(n301) );
  inv01 U20 ( .Y(n15), .A(n14) );
  or02 U21 ( .Y(n16), .A0(n294), .A1(n299) );
  inv02 U22 ( .Y(n17), .A(n16) );
  or02 U23 ( .Y(n18), .A0(n296), .A1(n299) );
  inv02 U24 ( .Y(n19), .A(n18) );
  or02 U25 ( .Y(n20), .A0(n298), .A1(n299) );
  inv02 U26 ( .Y(n21), .A(n20) );
  nand02 U27 ( .Y(n22), .A0(n47), .A1(n49) );
  inv02 U28 ( .Y(n23), .A(n22) );
  nand02 U29 ( .Y(n24), .A0(n51), .A1(n45) );
  inv02 U30 ( .Y(n25), .A(n24) );
  inv01 U31 ( .Y(n26), .A(n118) );
  inv01 U32 ( .Y(n27), .A(n174) );
  inv01 U33 ( .Y(n28), .A(n176) );
  inv01 U34 ( .Y(n29), .A(n63) );
  or02 U35 ( .Y(n30), .A0(n293), .A1(n300) );
  inv02 U36 ( .Y(n31), .A(n30) );
  or02 U37 ( .Y(n32), .A0(n293), .A1(n302) );
  inv02 U38 ( .Y(n33), .A(n32) );
  or02 U39 ( .Y(n34), .A0(n297), .A1(n302) );
  inv02 U40 ( .Y(n35), .A(n34) );
  or02 U41 ( .Y(n36), .A0(n301), .A1(n302) );
  inv02 U42 ( .Y(n37), .A(n36) );
  or02 U43 ( .Y(n38), .A0(n295), .A1(n300) );
  inv02 U44 ( .Y(n39), .A(n38) );
  or02 U45 ( .Y(n40), .A0(n295), .A1(n302) );
  inv02 U46 ( .Y(n41), .A(n40) );
  buf02 U47 ( .Y(n42), .A(U1_level_node_2__4__1_) );
  buf02 U48 ( .Y(n43), .A(U1_level_node_2__3__0_) );
  buf02 U49 ( .Y(n44), .A(U1_B_neg_correction_1_) );
  buf02 U50 ( .Y(n45), .A(U1_B_neg_correction_1_) );
  or02 U51 ( .Y(n46), .A0(n300), .A1(n303) );
  inv02 U52 ( .Y(n47), .A(n46) );
  or02 U53 ( .Y(n48), .A0(n293), .A1(n298) );
  inv02 U54 ( .Y(n49), .A(n48) );
  or02 U55 ( .Y(n50), .A0(n299), .A1(n302) );
  inv02 U56 ( .Y(n51), .A(n50) );
  or02 U57 ( .Y(n52), .A0(n292), .A1(n303) );
  inv02 U58 ( .Y(n53), .A(n52) );
  or02 U59 ( .Y(n54), .A0(n297), .A1(n298) );
  inv02 U60 ( .Y(n55), .A(n54) );
  or02 U61 ( .Y(n56), .A0(n296), .A1(n297) );
  inv02 U62 ( .Y(n57), .A(n56) );
  or02 U63 ( .Y(n58), .A0(n295), .A1(n298) );
  inv02 U64 ( .Y(n59), .A(n58) );
  inv02 U65 ( .Y(U1_level_node_2__4__0_), .A(n60) );
  inv02 U66 ( .Y(U1_level_node_2__5__1_), .A(n61) );
  inv02 U67 ( .Y(n62), .A(n57) );
  inv02 U68 ( .Y(n63), .A(U1_level_node_1__4__0_) );
  inv02 U69 ( .Y(n64), .A(n59) );
  nor02 U70 ( .Y(n65), .A0(n62), .A1(n66) );
  nor02 U71 ( .Y(n67), .A0(n63), .A1(n68) );
  nor02 U72 ( .Y(n69), .A0(n64), .A1(n70) );
  nor02 U73 ( .Y(n71), .A0(n64), .A1(n72) );
  nor02 U74 ( .Y(n60), .A0(n73), .A1(n74) );
  nor02 U75 ( .Y(n75), .A0(n63), .A1(n64) );
  nor02 U76 ( .Y(n76), .A0(n62), .A1(n64) );
  nor02 U77 ( .Y(n77), .A0(n62), .A1(n63) );
  nor02 U78 ( .Y(n61), .A0(n77), .A1(n78) );
  nor02 U79 ( .Y(n79), .A0(U1_level_node_1__4__0_), .A1(n59) );
  inv01 U80 ( .Y(n66), .A(n79) );
  nor02 U81 ( .Y(n80), .A0(n57), .A1(n59) );
  inv01 U82 ( .Y(n68), .A(n80) );
  nor02 U83 ( .Y(n81), .A0(n57), .A1(n29) );
  inv01 U84 ( .Y(n70), .A(n81) );
  nor02 U85 ( .Y(n82), .A0(n62), .A1(n63) );
  inv01 U86 ( .Y(n72), .A(n82) );
  nor02 U87 ( .Y(n83), .A0(n65), .A1(n67) );
  inv01 U88 ( .Y(n73), .A(n83) );
  nor02 U89 ( .Y(n84), .A0(n69), .A1(n71) );
  inv01 U90 ( .Y(n74), .A(n84) );
  nor02 U91 ( .Y(n85), .A0(n75), .A1(n76) );
  inv01 U92 ( .Y(n78), .A(n85) );
  or02 U93 ( .Y(n86), .A0(n292), .A1(n293) );
  inv02 U94 ( .Y(n87), .A(n86) );
  or02 U95 ( .Y(n88), .A0(n294), .A1(n303) );
  inv02 U96 ( .Y(n89), .A(n88) );
  inv02 U97 ( .Y(U1_level_node_2__8__0_), .A(n90) );
  inv02 U98 ( .Y(U1_level_node_2__9__0_), .A(n91) );
  inv02 U99 ( .Y(n92), .A(n87) );
  inv02 U100 ( .Y(n93), .A(U1_level_node_1__8__0_) );
  inv02 U101 ( .Y(n94), .A(n89) );
  nor02 U102 ( .Y(n95), .A0(n92), .A1(n96) );
  nor02 U103 ( .Y(n97), .A0(n93), .A1(n98) );
  nor02 U104 ( .Y(n99), .A0(n94), .A1(n100) );
  nor02 U105 ( .Y(n101), .A0(n94), .A1(n102) );
  nor02 U106 ( .Y(n90), .A0(n103), .A1(n104) );
  nor02 U107 ( .Y(n105), .A0(n93), .A1(n94) );
  nor02 U108 ( .Y(n106), .A0(n92), .A1(n94) );
  nor02 U109 ( .Y(n107), .A0(n92), .A1(n93) );
  nor02 U110 ( .Y(n91), .A0(n107), .A1(n108) );
  nor02 U111 ( .Y(n109), .A0(U1_level_node_1__8__0_), .A1(n89) );
  inv01 U112 ( .Y(n96), .A(n109) );
  nor02 U113 ( .Y(n110), .A0(n87), .A1(n89) );
  inv01 U114 ( .Y(n98), .A(n110) );
  nor02 U115 ( .Y(n111), .A0(n87), .A1(U1_level_node_1__8__0_) );
  inv01 U116 ( .Y(n100), .A(n111) );
  nor02 U117 ( .Y(n112), .A0(n92), .A1(n93) );
  inv01 U118 ( .Y(n102), .A(n112) );
  nor02 U119 ( .Y(n113), .A0(n95), .A1(n97) );
  inv01 U120 ( .Y(n103), .A(n113) );
  nor02 U121 ( .Y(n114), .A0(n99), .A1(n101) );
  inv01 U122 ( .Y(n104), .A(n114) );
  nor02 U123 ( .Y(n115), .A0(n105), .A1(n106) );
  inv01 U124 ( .Y(n108), .A(n115) );
  inv02 U125 ( .Y(U1_level_node_2__6__0_), .A(n116) );
  inv02 U126 ( .Y(U1_level_node_2__7__1_), .A(n117) );
  inv02 U127 ( .Y(n118), .A(U1_level_node_1__6__1_) );
  inv02 U128 ( .Y(n119), .A(U1_level_node_1__6__0_) );
  inv02 U129 ( .Y(n120), .A(U1_level_node_1__6__2_) );
  nor02 U130 ( .Y(n121), .A0(n118), .A1(n122) );
  nor02 U131 ( .Y(n123), .A0(n119), .A1(n124) );
  nor02 U132 ( .Y(n125), .A0(n120), .A1(n126) );
  nor02 U133 ( .Y(n127), .A0(n120), .A1(n128) );
  nor02 U134 ( .Y(n116), .A0(n129), .A1(n130) );
  nor02 U135 ( .Y(n131), .A0(n119), .A1(n120) );
  nor02 U136 ( .Y(n132), .A0(n118), .A1(n120) );
  nor02 U137 ( .Y(n133), .A0(n118), .A1(n119) );
  nor02 U138 ( .Y(n117), .A0(n133), .A1(n134) );
  nor02 U139 ( .Y(n135), .A0(U1_level_node_1__6__0_), .A1(
        U1_level_node_1__6__2_) );
  inv01 U140 ( .Y(n122), .A(n135) );
  nor02 U141 ( .Y(n136), .A0(n26), .A1(U1_level_node_1__6__2_) );
  inv01 U142 ( .Y(n124), .A(n136) );
  nor02 U143 ( .Y(n137), .A0(U1_level_node_1__6__1_), .A1(
        U1_level_node_1__6__0_) );
  inv01 U144 ( .Y(n126), .A(n137) );
  nor02 U145 ( .Y(n138), .A0(n118), .A1(n119) );
  inv01 U146 ( .Y(n128), .A(n138) );
  nor02 U147 ( .Y(n139), .A0(n121), .A1(n123) );
  inv01 U148 ( .Y(n129), .A(n139) );
  nor02 U149 ( .Y(n140), .A0(n125), .A1(n127) );
  inv01 U150 ( .Y(n130), .A(n140) );
  nor02 U151 ( .Y(n141), .A0(n131), .A1(n132) );
  inv01 U152 ( .Y(n134), .A(n141) );
  or02 U153 ( .Y(n142), .A0(n294), .A1(n297) );
  inv02 U154 ( .Y(n143), .A(n142) );
  or02 U155 ( .Y(n144), .A0(n295), .A1(n296) );
  inv02 U156 ( .Y(n145), .A(n144) );
  inv02 U157 ( .Y(U1_level_node_1__5__0_), .A(n146) );
  inv02 U158 ( .Y(U1_level_node_1__6__2_), .A(n147) );
  inv02 U159 ( .Y(n148), .A(n143) );
  inv02 U160 ( .Y(n149), .A(n288) );
  inv02 U161 ( .Y(n150), .A(n145) );
  nor02 U162 ( .Y(n151), .A0(n148), .A1(n152) );
  nor02 U163 ( .Y(n153), .A0(n149), .A1(n154) );
  nor02 U164 ( .Y(n155), .A0(n150), .A1(n156) );
  nor02 U165 ( .Y(n157), .A0(n150), .A1(n158) );
  nor02 U166 ( .Y(n146), .A0(n159), .A1(n160) );
  nor02 U167 ( .Y(n161), .A0(n149), .A1(n150) );
  nor02 U168 ( .Y(n162), .A0(n148), .A1(n150) );
  nor02 U169 ( .Y(n163), .A0(n148), .A1(n149) );
  nor02 U170 ( .Y(n147), .A0(n163), .A1(n164) );
  nor02 U171 ( .Y(n165), .A0(n288), .A1(n145) );
  inv01 U172 ( .Y(n152), .A(n165) );
  nor02 U173 ( .Y(n166), .A0(n143), .A1(n145) );
  inv01 U174 ( .Y(n154), .A(n166) );
  nor02 U175 ( .Y(n167), .A0(n143), .A1(n288) );
  inv01 U176 ( .Y(n156), .A(n167) );
  nor02 U177 ( .Y(n168), .A0(n148), .A1(n149) );
  inv01 U178 ( .Y(n158), .A(n168) );
  nor02 U179 ( .Y(n169), .A0(n151), .A1(n153) );
  inv01 U180 ( .Y(n159), .A(n169) );
  nor02 U181 ( .Y(n170), .A0(n155), .A1(n157) );
  inv01 U182 ( .Y(n160), .A(n170) );
  nor02 U183 ( .Y(n171), .A0(n161), .A1(n162) );
  inv01 U184 ( .Y(n164), .A(n171) );
  inv02 U185 ( .Y(U1_level_node_2__5__0_), .A(n172) );
  inv02 U186 ( .Y(U1_level_node_2__6__1_), .A(n173) );
  inv02 U187 ( .Y(n174), .A(U1_level_node_1__5__1_) );
  inv02 U188 ( .Y(n175), .A(U1_level_node_1__5__0_) );
  inv02 U189 ( .Y(n176), .A(U1_level_node_1__5__2_) );
  nor02 U190 ( .Y(n177), .A0(n174), .A1(n178) );
  nor02 U191 ( .Y(n179), .A0(n175), .A1(n180) );
  nor02 U192 ( .Y(n181), .A0(n176), .A1(n182) );
  nor02 U193 ( .Y(n183), .A0(n176), .A1(n184) );
  nor02 U194 ( .Y(n172), .A0(n185), .A1(n186) );
  nor02 U195 ( .Y(n187), .A0(n175), .A1(n176) );
  nor02 U196 ( .Y(n188), .A0(n174), .A1(n176) );
  nor02 U197 ( .Y(n189), .A0(n174), .A1(n175) );
  nor02 U198 ( .Y(n173), .A0(n189), .A1(n190) );
  nor02 U199 ( .Y(n191), .A0(U1_level_node_1__5__0_), .A1(
        U1_level_node_1__5__2_) );
  inv01 U200 ( .Y(n178), .A(n191) );
  nor02 U201 ( .Y(n192), .A0(n27), .A1(n28) );
  inv01 U202 ( .Y(n180), .A(n192) );
  nor02 U203 ( .Y(n193), .A0(U1_level_node_1__5__1_), .A1(
        U1_level_node_1__5__0_) );
  inv01 U204 ( .Y(n182), .A(n193) );
  nor02 U205 ( .Y(n194), .A0(n174), .A1(n175) );
  inv01 U206 ( .Y(n184), .A(n194) );
  nor02 U207 ( .Y(n195), .A0(n177), .A1(n179) );
  inv01 U208 ( .Y(n185), .A(n195) );
  nor02 U209 ( .Y(n196), .A0(n181), .A1(n183) );
  inv01 U210 ( .Y(n186), .A(n196) );
  nor02 U211 ( .Y(n197), .A0(n187), .A1(n188) );
  inv01 U212 ( .Y(n190), .A(n197) );
  nor02 U213 ( .Y(n198), .A0(n296), .A1(n303) );
  or02 U214 ( .Y(n199), .A0(n293), .A1(n296) );
  inv02 U215 ( .Y(n200), .A(n199) );
  or02 U216 ( .Y(n201), .A0(n293), .A1(n294) );
  inv02 U217 ( .Y(n202), .A(n201) );
  or02 U218 ( .Y(n203), .A0(n294), .A1(n295) );
  inv02 U219 ( .Y(n204), .A(n203) );
  inv04 U220 ( .Y(n303), .A(B[5]) );
  inv02 U221 ( .Y(U1_level_node_1__7__0_), .A(n205) );
  inv02 U222 ( .Y(U1_level_node_1__8__0_), .A(n206) );
  inv02 U223 ( .Y(n207), .A(n202) );
  inv02 U224 ( .Y(n208), .A(n284) );
  inv02 U225 ( .Y(n209), .A(U1_B_neg_correction_2_) );
  nor02 U226 ( .Y(n210), .A0(n207), .A1(n211) );
  nor02 U227 ( .Y(n212), .A0(n208), .A1(n213) );
  nor02 U228 ( .Y(n214), .A0(n209), .A1(n215) );
  nor02 U229 ( .Y(n216), .A0(n209), .A1(n217) );
  nor02 U230 ( .Y(n205), .A0(n218), .A1(n219) );
  nor02 U231 ( .Y(n220), .A0(n208), .A1(n209) );
  nor02 U232 ( .Y(n221), .A0(n207), .A1(n209) );
  nor02 U233 ( .Y(n222), .A0(n207), .A1(n208) );
  nor02 U234 ( .Y(n206), .A0(n222), .A1(n223) );
  nor02 U235 ( .Y(n224), .A0(n284), .A1(n198) );
  inv01 U236 ( .Y(n211), .A(n224) );
  nor02 U237 ( .Y(n225), .A0(n202), .A1(n3) );
  inv01 U238 ( .Y(n213), .A(n225) );
  nor02 U239 ( .Y(n226), .A0(n202), .A1(n284) );
  inv01 U240 ( .Y(n215), .A(n226) );
  nor02 U241 ( .Y(n227), .A0(n207), .A1(n208) );
  inv01 U242 ( .Y(n217), .A(n227) );
  nor02 U243 ( .Y(n228), .A0(n210), .A1(n212) );
  inv01 U244 ( .Y(n218), .A(n228) );
  nor02 U245 ( .Y(n229), .A0(n214), .A1(n216) );
  inv01 U246 ( .Y(n219), .A(n229) );
  nor02 U247 ( .Y(n230), .A0(n220), .A1(n221) );
  inv01 U248 ( .Y(n223), .A(n230) );
  inv02 U249 ( .Y(U1_level_node_1__6__0_), .A(n231) );
  inv02 U250 ( .Y(U1_level_node_1__7__1_), .A(n232) );
  inv02 U251 ( .Y(n233), .A(n204) );
  inv02 U252 ( .Y(n234), .A(n286) );
  inv02 U253 ( .Y(n235), .A(n200) );
  nor02 U254 ( .Y(n236), .A0(n233), .A1(n237) );
  nor02 U255 ( .Y(n238), .A0(n234), .A1(n239) );
  nor02 U256 ( .Y(n240), .A0(n235), .A1(n241) );
  nor02 U257 ( .Y(n242), .A0(n235), .A1(n243) );
  nor02 U258 ( .Y(n231), .A0(n244), .A1(n245) );
  nor02 U259 ( .Y(n246), .A0(n234), .A1(n235) );
  nor02 U260 ( .Y(n247), .A0(n233), .A1(n235) );
  nor02 U261 ( .Y(n248), .A0(n233), .A1(n234) );
  nor02 U262 ( .Y(n232), .A0(n248), .A1(n249) );
  nor02 U263 ( .Y(n250), .A0(n286), .A1(n200) );
  inv01 U264 ( .Y(n237), .A(n250) );
  nor02 U265 ( .Y(n251), .A0(n204), .A1(n200) );
  inv01 U266 ( .Y(n239), .A(n251) );
  nor02 U267 ( .Y(n252), .A0(n204), .A1(n286) );
  inv01 U268 ( .Y(n241), .A(n252) );
  nor02 U269 ( .Y(n253), .A0(n233), .A1(n234) );
  inv01 U270 ( .Y(n243), .A(n253) );
  nor02 U271 ( .Y(n254), .A0(n236), .A1(n238) );
  inv01 U272 ( .Y(n244), .A(n254) );
  nor02 U273 ( .Y(n255), .A0(n240), .A1(n242) );
  inv01 U274 ( .Y(n245), .A(n255) );
  nor02 U275 ( .Y(n256), .A0(n246), .A1(n247) );
  inv01 U276 ( .Y(n249), .A(n256) );
  inv02 U277 ( .Y(U1_level_node_2__7__0_), .A(n257) );
  inv02 U278 ( .Y(U1_level_node_2__8__1_), .A(n258) );
  inv02 U279 ( .Y(n259), .A(U1_level_node_1__7__1_) );
  inv02 U280 ( .Y(n260), .A(U1_level_node_1__7__0_) );
  inv02 U281 ( .Y(n261), .A(n25) );
  nor02 U282 ( .Y(n262), .A0(n259), .A1(n263) );
  nor02 U283 ( .Y(n264), .A0(n260), .A1(n265) );
  nor02 U284 ( .Y(n266), .A0(n261), .A1(n267) );
  nor02 U285 ( .Y(n268), .A0(n261), .A1(n269) );
  nor02 U286 ( .Y(n257), .A0(n270), .A1(n271) );
  nor02 U287 ( .Y(n272), .A0(n260), .A1(n261) );
  nor02 U288 ( .Y(n273), .A0(n259), .A1(n261) );
  nor02 U289 ( .Y(n274), .A0(n259), .A1(n260) );
  nor02 U290 ( .Y(n258), .A0(n274), .A1(n275) );
  nor02 U291 ( .Y(n276), .A0(U1_level_node_1__7__0_), .A1(n25) );
  inv01 U292 ( .Y(n263), .A(n276) );
  nor02 U293 ( .Y(n277), .A0(U1_level_node_1__7__1_), .A1(n25) );
  inv01 U294 ( .Y(n265), .A(n277) );
  nor02 U295 ( .Y(n278), .A0(U1_level_node_1__7__1_), .A1(
        U1_level_node_1__7__0_) );
  inv01 U296 ( .Y(n267), .A(n278) );
  nor02 U297 ( .Y(n279), .A0(n259), .A1(n260) );
  inv01 U298 ( .Y(n269), .A(n279) );
  nor02 U299 ( .Y(n280), .A0(n262), .A1(n264) );
  inv01 U300 ( .Y(n270), .A(n280) );
  nor02 U301 ( .Y(n281), .A0(n266), .A1(n268) );
  inv01 U302 ( .Y(n271), .A(n281) );
  nor02 U303 ( .Y(n282), .A0(n272), .A1(n273) );
  inv01 U304 ( .Y(n275), .A(n282) );
  or02 U305 ( .Y(n283), .A0(n292), .A1(n295) );
  inv02 U306 ( .Y(n284), .A(n283) );
  or02 U307 ( .Y(n285), .A0(n292), .A1(n297) );
  inv02 U308 ( .Y(n286), .A(n285) );
  or02 U309 ( .Y(n287), .A0(n292), .A1(n299) );
  inv02 U310 ( .Y(n288), .A(n287) );
  or02 U311 ( .Y(n289), .A0(n300), .A1(n301) );
  inv02 U312 ( .Y(PRODUCT[0]), .A(n289) );
  inv02 U313 ( .Y(n299), .A(B[1]) );
  inv02 U314 ( .Y(n295), .A(B[3]) );
  inv02 U315 ( .Y(n294), .A(A[3]) );
  inv02 U316 ( .Y(n297), .A(B[2]) );
  inv02 U317 ( .Y(n301), .A(B[0]) );
  inv02 U318 ( .Y(n298), .A(A[1]) );
  inv02 U319 ( .Y(n293), .A(B[4]) );
  inv02 U320 ( .Y(n292), .A(A[4]) );
  inv02 U321 ( .Y(n300), .A(A[0]) );
  inv02 U322 ( .Y(n302), .A(A[5]) );
  xor2 U323 ( .Y(U1_level_node_1__5__1_), .A0(n49), .A1(n47) );
  xor2 U324 ( .Y(U1_level_node_1__6__1_), .A0(n44), .A1(n51) );
  mul_24_DW01_add_11_0 U1_U9720 ( .A({1'b0, U1_level_node_3__10__0_, 
        U1_level_node_3__9__0_, U1_level_node_3__8__0_, U1_level_node_3__7__0_, 
        U1_level_node_3__6__0_, U1_level_node_3__5__0_, U1_level_node_3__4__0_, 
        U1_level_node_3__3__0_, U1_level_node_3__2__0_, n2}), .B({1'b0, n9, 
        U1_level_node_3__9__1_, U1_level_node_3__8__1_, U1_level_node_3__7__1_, 
        U1_level_node_3__6__1_, U1_level_node_3__5__1_, U1_level_node_3__4__1_, 
        U1_level_node_3__3__1_, n5, n7}), .CI(1'b0), .SUM(PRODUCT[11:1]) );
  nor02 U325 ( .Y(U1_B_neg_correction_2_), .A0(n296), .A1(n303) );
  nor02 U326 ( .Y(U1_B_neg_correction_1_), .A0(n298), .A1(n303) );
  hadd1 U1_U3220_1_4 ( .S(U1_level_node_1__4__0_), .CO(U1_level_node_1__5__2_), 
        .A(n13), .B(n17) );
  hadd1 U1_U3220_2_3 ( .S(U1_level_node_2__3__0_), .CO(U1_level_node_2__4__1_), 
        .A(n15), .B(n19) );
  fadd1 U1_U3140_3_9_0 ( .S(U1_level_node_3__9__0_), .CO(
        U1_level_node_3__10__0_), .A(U1_level_node_2__9__0_), .B(n53), .CI(n33) );
  fadd1 U1_U3140_3_8_0 ( .S(U1_level_node_3__8__0_), .CO(
        U1_level_node_3__9__1_), .A(U1_level_node_2__8__0_), .B(
        U1_level_node_2__8__1_), .CI(n41) );
  fadd1 U1_U3140_3_7_0 ( .S(U1_level_node_3__7__0_), .CO(
        U1_level_node_3__8__1_), .A(U1_level_node_2__7__0_), .B(
        U1_level_node_2__7__1_), .CI(n35) );
  fadd1 U1_U3140_3_6_0 ( .S(U1_level_node_3__6__0_), .CO(
        U1_level_node_3__7__1_), .A(U1_level_node_2__6__0_), .B(
        U1_level_node_2__6__1_), .CI(n23) );
  fadd1 U1_U3140_3_5_0 ( .S(U1_level_node_3__5__0_), .CO(
        U1_level_node_3__6__1_), .A(U1_level_node_2__5__0_), .B(
        U1_level_node_2__5__1_), .CI(n37) );
  fadd1 U1_U3140_3_4_0 ( .S(U1_level_node_3__4__0_), .CO(
        U1_level_node_3__5__1_), .A(U1_level_node_2__4__0_), .B(n42), .CI(n31)
         );
  fadd1 U1_U3140_3_3_0 ( .S(U1_level_node_3__3__0_), .CO(
        U1_level_node_3__4__1_), .A(n43), .B(n55), .CI(n39) );
  hadd1 U1_U3220_3_2 ( .S(U1_level_node_3__2__0_), .CO(U1_level_node_3__3__1_), 
        .A(n11), .B(n21) );
endmodule


module mul_24 ( clk_i, fracta_i, fractb_i, signa_i, signb_i, start_i, fract_o, 
        sign_o, ready_o );
  input [23:0] fracta_i;
  input [23:0] fractb_i;
  output [47:0] fract_o;
  input clk_i, signa_i, signb_i, start_i;
  output sign_o, ready_o;
  wire   s_signb_i, prod_a_b_3__23_, prod_a_b_3__22_, prod_a_b_3__21_,
         prod_a_b_3__20_, prod_a_b_3__19_, prod_a_b_3__18_, prod_a_b_3__17_,
         prod_a_b_3__16_, prod_a_b_3__15_, prod_a_b_3__14_, prod_a_b_3__13_,
         prod_a_b_3__12_, prod_a_b_3__11_, prod_a_b_3__10_, prod_a_b_3__9_,
         prod_a_b_3__8_, prod_a_b_3__7_, prod_a_b_3__6_, prod_a_b_3__5_,
         prod_a_b_3__4_, prod_a_b_3__3_, prod_a_b_3__2_, prod_a_b_3__1_,
         prod_a_b_3__0_, prod_a_b_2__35_, prod_a_b_2__34_, prod_a_b_2__33_,
         prod_a_b_2__32_, prod_a_b_2__31_, prod_a_b_2__30_, prod_a_b_2__29_,
         prod_a_b_2__28_, prod_a_b_2__27_, prod_a_b_2__26_, prod_a_b_2__25_,
         prod_a_b_2__24_, prod_a_b_2__23_, prod_a_b_2__22_, prod_a_b_2__21_,
         prod_a_b_2__20_, prod_a_b_2__19_, prod_a_b_2__18_, prod_a_b_2__17_,
         prod_a_b_2__16_, prod_a_b_2__15_, prod_a_b_2__14_, prod_a_b_2__13_,
         prod_a_b_2__12_, prod_a_b_1__35_, prod_a_b_1__34_, prod_a_b_1__33_,
         prod_a_b_1__32_, prod_a_b_1__31_, prod_a_b_1__30_, prod_a_b_1__29_,
         prod_a_b_1__28_, prod_a_b_1__27_, prod_a_b_1__26_, prod_a_b_1__25_,
         prod_a_b_1__24_, prod_a_b_1__23_, prod_a_b_1__22_, prod_a_b_1__21_,
         prod_a_b_1__20_, prod_a_b_1__19_, prod_a_b_1__18_, prod_a_b_1__17_,
         prod_a_b_1__16_, prod_a_b_1__15_, prod_a_b_1__14_, prod_a_b_1__13_,
         prod_a_b_1__12_, prod_a_b_0__47_, prod_a_b_0__46_, prod_a_b_0__45_,
         prod_a_b_0__44_, prod_a_b_0__43_, prod_a_b_0__42_, prod_a_b_0__41_,
         prod_a_b_0__40_, prod_a_b_0__39_, prod_a_b_0__38_, prod_a_b_0__37_,
         prod_a_b_0__36_, prod_a_b_0__35_, prod_a_b_0__34_, prod_a_b_0__33_,
         prod_a_b_0__32_, prod_a_b_0__31_, prod_a_b_0__30_, prod_a_b_0__29_,
         prod_a_b_0__28_, prod_a_b_0__27_, prod_a_b_0__26_, prod_a_b_0__25_,
         prod_a_b_0__24_, s_state, s_state83, count_2_, count_1_, count_0_,
         n____return437_11_, n____return437_10_, n____return437_9_,
         n____return437_8_, n____return437_7_, n____return437_6_,
         n____return437_5_, n____return437_4_, n____return437_3_,
         n____return437_2_, n____return437_1_, n____return437_0_,
         member360_1__3_, member360_1__1_, n____return792_11_,
         n____return792_10_, n____return792_9_, n____return792_8_,
         n____return792_7_, n____return792_6_, n____return792_5_,
         n____return792_4_, n____return792_3_, n____return792_2_,
         n____return792_1_, n____return792_0_, member638_2__3_,
         n____return1150_11_, n____return1150_10_, n____return1150_9_,
         n____return1150_8_, n____return1150_7_, n____return1150_6_,
         n____return1150_5_, n____return1150_4_, n____return1150_3_,
         n____return1150_2_, n____return1150_1_, n____return1150_0_,
         member996_4__4_, member996_4__2_, member996_4__1_,
         n____return1508_11_, n____return1508_10_, n____return1508_9_,
         n____return1508_8_, n____return1508_7_, n____return1508_6_,
         n____return1508_5_, n____return1508_4_, n____return1508_3_,
         n____return1508_2_, n____return1508_1_, n____return1508_0_,
         n____return2214_23_, n____return2214_22_, n____return2214_21_,
         n____return2214_20_, n____return2214_19_, n____return2214_18_,
         n____return2214_17_, n____return2214_16_, n____return2214_15_,
         n____return2214_14_, n____return2214_13_, n____return2214_12_,
         n____return2214_11_, n____return2214_10_, n____return2214_9_,
         n____return2214_8_, n____return2214_7_, n____return2214_6_,
         n____return2214_5_, n____return2214_4_, n____return2214_3_,
         n____return2214_2_, n____return2214_1_, n____return2214_0_,
         member1796_0__23_, member1796_0__22_, member1796_0__21_,
         member1796_0__20_, member1796_0__19_, member1796_0__18_,
         member1796_0__17_, member1796_0__16_, member1796_0__15_,
         member1796_0__14_, member1796_0__13_, member1796_0__12_,
         member1796_0__11_, member1796_0__10_, member1796_0__9_,
         member1796_0__8_, member1796_0__7_, member1796_0__6_,
         member1796_0__5_, member1796_0__4_, member1796_0__3_,
         member1796_0__2_, member1796_0__1_, member1796_0__0_,
         member1883_1__23_, member1883_1__22_, member1883_1__21_,
         member1883_1__20_, member1883_1__19_, member1883_1__18_,
         member1883_1__17_, member1883_1__16_, member1883_1__15_,
         member1883_1__14_, member1883_1__13_, member1883_1__12_,
         member1883_1__11_, member1883_1__10_, member1883_1__9_,
         member1883_1__8_, member1883_1__7_, member1883_1__6_,
         member1883_1__5_, member1883_1__4_, member1883_1__3_,
         member1883_1__2_, member1883_1__1_, member1883_1__0_,
         member2010_2__23_, member2010_2__22_, member2010_2__21_,
         member2010_2__20_, member2010_2__19_, member2010_2__18_,
         member2010_2__17_, member2010_2__16_, member2010_2__15_,
         member2010_2__14_, member2010_2__13_, member2010_2__12_,
         member2010_2__11_, member2010_2__10_, member2010_2__9_,
         member2010_2__8_, member2010_2__7_, member2010_2__6_,
         member2010_2__5_, member2010_2__4_, member2010_2__3_,
         member2010_2__2_, member2010_2__1_, member2010_2__0_,
         member2137_3__23_, member2137_3__22_, member2137_3__21_,
         member2137_3__20_, member2137_3__19_, member2137_3__18_,
         member2137_3__17_, member2137_3__16_, member2137_3__15_,
         member2137_3__14_, member2137_3__13_, member2137_3__12_,
         member2137_3__11_, member2137_3__10_, member2137_3__9_,
         member2137_3__8_, member2137_3__7_, member2137_3__6_,
         member2137_3__5_, member2137_3__4_, member2137_3__3_,
         member2137_3__2_, member2137_3__1_, member2137_3__0_,
         n____return2087_23_, n____return2087_22_, n____return2087_21_,
         n____return2087_20_, n____return2087_19_, n____return2087_18_,
         n____return2087_17_, n____return2087_16_, n____return2087_15_,
         n____return2087_14_, n____return2087_13_, n____return2087_12_,
         n____return2087_11_, n____return2087_10_, n____return2087_9_,
         n____return2087_8_, n____return2087_7_, n____return2087_6_,
         n____return2087_5_, n____return2087_4_, n____return2087_3_,
         n____return2087_2_, n____return2087_1_, n____return2087_0_,
         n____return1960_23_, n____return1960_22_, n____return1960_21_,
         n____return1960_20_, n____return1960_19_, n____return1960_18_,
         n____return1960_17_, n____return1960_16_, n____return1960_15_,
         n____return1960_14_, n____return1960_13_, n____return1960_12_,
         n____return1960_11_, n____return1960_10_, n____return1960_9_,
         n____return1960_8_, n____return1960_7_, n____return1960_6_,
         n____return1960_5_, n____return1960_4_, n____return1960_3_,
         n____return1960_2_, n____return1960_1_, n____return1960_0_,
         n____return2414_36_, n____return2414_35_, n____return2414_34_,
         n____return2414_33_, n____return2414_32_, n____return2414_31_,
         n____return2414_30_, n____return2414_29_, n____return2414_28_,
         n____return2414_27_, n____return2414_26_, n____return2414_25_,
         n____return2414_24_, n____return2414_23_, n____return2414_22_,
         n____return2414_21_, n____return2414_20_, n____return2414_19_,
         n____return2414_18_, n____return2414_17_, n____return2414_16_,
         n____return2414_15_, n____return2414_14_, n____return2414_13_,
         n____return2414_12_, n____return2414_11_, n____return2414_10_,
         n____return2414_9_, n____return2414_8_, n____return2414_7_,
         n____return2414_6_, n____return2414_5_, n____return2414_4_,
         n____return2414_3_, n____return2414_2_, n____return2414_1_,
         n____return2414_0_, n____return2374_47_, n____return2374_46_,
         n____return2374_45_, n____return2374_44_, n____return2374_43_,
         n____return2374_42_, n____return2374_41_, n____return2374_40_,
         n____return2374_39_, n____return2374_38_, n____return2374_37_,
         n____return2374_36_, n____return2374_35_, n____return2374_34_,
         n____return2374_33_, n____return2374_32_, n____return2374_31_,
         n____return2374_30_, n____return2374_29_, n____return2374_28_,
         n____return2374_27_, n____return2374_26_, n____return2374_25_,
         n____return2374_24_, n____return2374_23_, n____return2374_22_,
         n____return2374_21_, n____return2374_20_, n____return2374_19_,
         n____return2374_18_, n____return2374_17_, n____return2374_16_,
         n____return2374_15_, n____return2374_14_, n____return2374_13_,
         n____return2374_12_, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23;
  wire   [383:0] larray;

  dff count_reg_0_ ( .Q(count_0_), .D(n6283), .CLK(clk_i) );
  dff count_reg_1_ ( .Q(count_1_), .D(n6285), .CLK(clk_i) );
  dff count_reg_2_ ( .Q(count_2_), .D(n5808), .CLK(clk_i) );
  dff prod2_reg_3__3__23_ ( .Q(larray[383]), .D(n5938), .CLK(clk_i) );
  dff prod2_reg_3__3__22_ ( .Q(larray[382]), .D(n5834), .CLK(clk_i) );
  dff prod2_reg_3__3__21_ ( .Q(larray[381]), .D(n5996), .CLK(clk_i) );
  dff prod2_reg_3__3__20_ ( .Q(larray[380]), .D(n5966), .CLK(clk_i) );
  dff prod2_reg_3__3__19_ ( .Q(larray[379]), .D(n5962), .CLK(clk_i) );
  dff prod2_reg_3__3__18_ ( .Q(larray[378]), .D(n5980), .CLK(clk_i) );
  dff prod2_reg_3__3__17_ ( .Q(larray[377]), .D(n5900), .CLK(clk_i) );
  dff prod2_reg_3__3__16_ ( .Q(larray[376]), .D(n5866), .CLK(clk_i) );
  dff prod2_reg_3__3__15_ ( .Q(larray[375]), .D(n5992), .CLK(clk_i) );
  dff prod2_reg_3__3__14_ ( .Q(larray[374]), .D(n5978), .CLK(clk_i) );
  dff prod2_reg_3__3__13_ ( .Q(larray[373]), .D(n5942), .CLK(clk_i) );
  dff prod2_reg_3__3__12_ ( .Q(larray[372]), .D(n5902), .CLK(clk_i) );
  dff prod2_reg_3__3__11_ ( .Q(larray[371]), .D(n4301), .CLK(clk_i) );
  dff prod2_reg_3__3__10_ ( .Q(larray[370]), .D(n6232), .CLK(clk_i) );
  dff prod2_reg_3__3__9_ ( .Q(larray[369]), .D(n6200), .CLK(clk_i) );
  dff prod2_reg_3__3__8_ ( .Q(larray[368]), .D(n6197), .CLK(clk_i) );
  dff prod2_reg_3__3__7_ ( .Q(larray[367]), .D(n6195), .CLK(clk_i) );
  dff prod2_reg_3__3__6_ ( .Q(larray[366]), .D(n6259), .CLK(clk_i) );
  dff prod2_reg_3__3__5_ ( .Q(larray[365]), .D(n6227), .CLK(clk_i) );
  dff prod2_reg_3__3__4_ ( .Q(larray[364]), .D(n6174), .CLK(clk_i) );
  dff prod2_reg_3__3__3_ ( .Q(larray[363]), .D(n6196), .CLK(clk_i) );
  dff prod2_reg_3__3__2_ ( .Q(larray[362]), .D(n6175), .CLK(clk_i) );
  dff prod2_reg_3__3__1_ ( .Q(larray[361]), .D(n6143), .CLK(clk_i) );
  dff prod2_reg_3__3__0_ ( .Q(larray[360]), .D(n6274), .CLK(clk_i) );
  dff prod2_reg_3__2__23_ ( .Q(larray[359]), .D(n5986), .CLK(clk_i) );
  dff prod2_reg_3__2__22_ ( .Q(larray[358]), .D(n5990), .CLK(clk_i) );
  dff prod2_reg_3__2__21_ ( .Q(larray[357]), .D(n5998), .CLK(clk_i) );
  dff prod2_reg_3__2__20_ ( .Q(larray[356]), .D(n5956), .CLK(clk_i) );
  dff prod2_reg_3__2__19_ ( .Q(larray[355]), .D(n5988), .CLK(clk_i) );
  dff prod2_reg_3__2__18_ ( .Q(larray[354]), .D(n6000), .CLK(clk_i) );
  dff prod2_reg_3__2__17_ ( .Q(larray[353]), .D(n6144), .CLK(clk_i) );
  dff prod2_reg_3__2__16_ ( .Q(larray[352]), .D(n6205), .CLK(clk_i) );
  dff prod2_reg_3__2__15_ ( .Q(larray[351]), .D(n6247), .CLK(clk_i) );
  dff prod2_reg_3__2__14_ ( .Q(larray[350]), .D(n6226), .CLK(clk_i) );
  dff prod2_reg_3__2__13_ ( .Q(larray[349]), .D(n6186), .CLK(clk_i) );
  dff prod2_reg_3__2__12_ ( .Q(larray[348]), .D(n6231), .CLK(clk_i) );
  dff prod2_reg_3__2__11_ ( .Q(larray[347]), .D(n6222), .CLK(clk_i) );
  dff prod2_reg_3__2__10_ ( .Q(larray[346]), .D(n6194), .CLK(clk_i) );
  dff prod2_reg_3__2__9_ ( .Q(larray[345]), .D(n6198), .CLK(clk_i) );
  dff prod2_reg_3__2__8_ ( .Q(larray[344]), .D(n4328), .CLK(clk_i) );
  dff prod2_reg_3__2__7_ ( .Q(larray[343]), .D(n6137), .CLK(clk_i) );
  dff prod2_reg_3__2__6_ ( .Q(larray[342]), .D(n4330), .CLK(clk_i) );
  dff prod2_reg_3__2__5_ ( .Q(larray[341]), .D(n5904), .CLK(clk_i) );
  dff prod2_reg_3__2__4_ ( .Q(larray[340]), .D(n5912), .CLK(clk_i) );
  dff prod2_reg_3__2__3_ ( .Q(larray[339]), .D(n5870), .CLK(clk_i) );
  dff prod2_reg_3__2__2_ ( .Q(larray[338]), .D(n5908), .CLK(clk_i) );
  dff prod2_reg_3__2__1_ ( .Q(larray[337]), .D(n5982), .CLK(clk_i) );
  dff prod2_reg_3__2__0_ ( .Q(larray[336]), .D(n5910), .CLK(clk_i) );
  dff prod2_reg_3__1__23_ ( .Q(larray[335]), .D(n5868), .CLK(clk_i) );
  dff prod2_reg_3__1__22_ ( .Q(larray[334]), .D(n5972), .CLK(clk_i) );
  dff prod2_reg_3__1__21_ ( .Q(larray[333]), .D(n5906), .CLK(clk_i) );
  dff prod2_reg_3__1__20_ ( .Q(larray[332]), .D(n5994), .CLK(clk_i) );
  dff prod2_reg_3__1__19_ ( .Q(larray[331]), .D(n5946), .CLK(clk_i) );
  dff prod2_reg_3__1__18_ ( .Q(larray[330]), .D(n5898), .CLK(clk_i) );
  dff prod2_reg_3__1__17_ ( .Q(larray[329]), .D(n6159), .CLK(clk_i) );
  dff prod2_reg_3__1__16_ ( .Q(larray[328]), .D(n6201), .CLK(clk_i) );
  dff prod2_reg_3__1__15_ ( .Q(larray[327]), .D(n6184), .CLK(clk_i) );
  dff prod2_reg_3__1__14_ ( .Q(larray[326]), .D(n6185), .CLK(clk_i) );
  dff prod2_reg_3__1__13_ ( .Q(larray[325]), .D(n6245), .CLK(clk_i) );
  dff prod2_reg_3__1__12_ ( .Q(larray[324]), .D(n6224), .CLK(clk_i) );
  dff prod2_reg_3__1__11_ ( .Q(larray[323]), .D(n6230), .CLK(clk_i) );
  dff prod2_reg_3__1__10_ ( .Q(larray[322]), .D(n4350), .CLK(clk_i) );
  dff prod2_reg_3__1__9_ ( .Q(larray[321]), .D(n6207), .CLK(clk_i) );
  dff prod2_reg_3__1__8_ ( .Q(larray[320]), .D(n6182), .CLK(clk_i) );
  dff prod2_reg_3__1__7_ ( .Q(larray[319]), .D(n6138), .CLK(clk_i) );
  dff prod2_reg_3__1__6_ ( .Q(larray[318]), .D(n6266), .CLK(clk_i) );
  dff prod2_reg_3__1__5_ ( .Q(larray[317]), .D(n5948), .CLK(clk_i) );
  dff prod2_reg_3__1__4_ ( .Q(larray[316]), .D(n5940), .CLK(clk_i) );
  dff prod2_reg_3__1__3_ ( .Q(larray[315]), .D(n5960), .CLK(clk_i) );
  dff prod2_reg_3__1__2_ ( .Q(larray[314]), .D(n5954), .CLK(clk_i) );
  dff prod2_reg_3__1__1_ ( .Q(larray[313]), .D(n5874), .CLK(clk_i) );
  dff prod2_reg_3__1__0_ ( .Q(larray[312]), .D(n5976), .CLK(clk_i) );
  dff prod2_reg_3__0__23_ ( .Q(larray[311]), .D(n4361), .CLK(clk_i) );
  dff prod2_reg_3__0__22_ ( .Q(larray[310]), .D(n6209), .CLK(clk_i) );
  dff prod2_reg_3__0__21_ ( .Q(larray[309]), .D(n6236), .CLK(clk_i) );
  dff prod2_reg_3__0__20_ ( .Q(larray[308]), .D(n6225), .CLK(clk_i) );
  dff prod2_reg_3__0__19_ ( .Q(larray[307]), .D(n6239), .CLK(clk_i) );
  dff prod2_reg_3__0__18_ ( .Q(larray[306]), .D(n6234), .CLK(clk_i) );
  dff prod2_reg_3__0__17_ ( .Q(larray[305]), .D(n6215), .CLK(clk_i) );
  dff prod2_reg_3__0__16_ ( .Q(larray[304]), .D(n6256), .CLK(clk_i) );
  dff prod2_reg_3__0__15_ ( .Q(larray[303]), .D(n6166), .CLK(clk_i) );
  dff prod2_reg_3__0__14_ ( .Q(larray[302]), .D(n6167), .CLK(clk_i) );
  dff prod2_reg_3__0__13_ ( .Q(larray[301]), .D(n6136), .CLK(clk_i) );
  dff prod2_reg_3__0__12_ ( .Q(larray[300]), .D(n6265), .CLK(clk_i) );
  dff prod2_reg_3__0__11_ ( .Q(larray[299]), .D(n5876), .CLK(clk_i) );
  dff prod2_reg_3__0__10_ ( .Q(larray[298]), .D(n5964), .CLK(clk_i) );
  dff prod2_reg_3__0__9_ ( .Q(larray[297]), .D(n5970), .CLK(clk_i) );
  dff prod2_reg_3__0__8_ ( .Q(larray[296]), .D(n5842), .CLK(clk_i) );
  dff prod2_reg_3__0__7_ ( .Q(larray[295]), .D(n5950), .CLK(clk_i) );
  dff prod2_reg_3__0__6_ ( .Q(larray[294]), .D(n5968), .CLK(clk_i) );
  dff prod2_reg_3__0__5_ ( .Q(larray[293]), .D(n5944), .CLK(clk_i) );
  dff prod2_reg_3__0__4_ ( .Q(larray[292]), .D(n5974), .CLK(clk_i) );
  dff prod2_reg_3__0__3_ ( .Q(larray[291]), .D(n5958), .CLK(clk_i) );
  dff prod2_reg_3__0__2_ ( .Q(larray[290]), .D(n5984), .CLK(clk_i) );
  dff prod2_reg_3__0__1_ ( .Q(larray[289]), .D(n5872), .CLK(clk_i) );
  dff prod2_reg_3__0__0_ ( .Q(larray[288]), .D(n5952), .CLK(clk_i) );
  dff prod2_reg_2__3__23_ ( .Q(larray[287]), .D(n5626), .CLK(clk_i) );
  dff prod2_reg_2__3__22_ ( .Q(larray[286]), .D(n5678), .CLK(clk_i) );
  dff prod2_reg_2__3__21_ ( .Q(larray[285]), .D(n5764), .CLK(clk_i) );
  dff prod2_reg_2__3__20_ ( .Q(larray[284]), .D(n5650), .CLK(clk_i) );
  dff prod2_reg_2__3__19_ ( .Q(larray[283]), .D(n5654), .CLK(clk_i) );
  dff prod2_reg_2__3__18_ ( .Q(larray[282]), .D(n5772), .CLK(clk_i) );
  dff prod2_reg_2__3__17_ ( .Q(larray[281]), .D(n5634), .CLK(clk_i) );
  dff prod2_reg_2__3__16_ ( .Q(larray[280]), .D(n5640), .CLK(clk_i) );
  dff prod2_reg_2__3__15_ ( .Q(larray[279]), .D(n5760), .CLK(clk_i) );
  dff prod2_reg_2__3__14_ ( .Q(larray[278]), .D(n5648), .CLK(clk_i) );
  dff prod2_reg_2__3__13_ ( .Q(larray[277]), .D(n5652), .CLK(clk_i) );
  dff prod2_reg_2__3__12_ ( .Q(larray[276]), .D(n5776), .CLK(clk_i) );
  dff prod2_reg_2__3__11_ ( .Q(larray[275]), .D(n6151), .CLK(clk_i) );
  dff prod2_reg_2__3__10_ ( .Q(larray[274]), .D(n6193), .CLK(clk_i) );
  dff prod2_reg_2__3__9_ ( .Q(larray[273]), .D(n6250), .CLK(clk_i) );
  dff prod2_reg_2__3__8_ ( .Q(larray[272]), .D(n6258), .CLK(clk_i) );
  dff prod2_reg_2__3__7_ ( .Q(larray[271]), .D(n4401), .CLK(clk_i) );
  dff prod2_reg_2__3__6_ ( .Q(larray[270]), .D(n6216), .CLK(clk_i) );
  dff prod2_reg_2__3__5_ ( .Q(larray[269]), .D(n6251), .CLK(clk_i) );
  dff prod2_reg_2__3__4_ ( .Q(larray[268]), .D(n4404), .CLK(clk_i) );
  dff prod2_reg_2__3__3_ ( .Q(larray[267]), .D(n6228), .CLK(clk_i) );
  dff prod2_reg_2__3__2_ ( .Q(larray[266]), .D(n6176), .CLK(clk_i) );
  dff prod2_reg_2__3__1_ ( .Q(larray[265]), .D(n6141), .CLK(clk_i) );
  dff prod2_reg_2__3__0_ ( .Q(larray[264]), .D(n4408), .CLK(clk_i) );
  dff prod2_reg_2__2__23_ ( .Q(larray[263]), .D(n5660), .CLK(clk_i) );
  dff prod2_reg_2__2__22_ ( .Q(larray[262]), .D(n5682), .CLK(clk_i) );
  dff prod2_reg_2__2__21_ ( .Q(larray[261]), .D(n5750), .CLK(clk_i) );
  dff prod2_reg_2__2__20_ ( .Q(larray[260]), .D(n5632), .CLK(clk_i) );
  dff prod2_reg_2__2__19_ ( .Q(larray[259]), .D(n5674), .CLK(clk_i) );
  dff prod2_reg_2__2__18_ ( .Q(larray[258]), .D(n5758), .CLK(clk_i) );
  dff prod2_reg_2__2__17_ ( .Q(larray[257]), .D(n6158), .CLK(clk_i) );
  dff prod2_reg_2__2__16_ ( .Q(larray[256]), .D(n6252), .CLK(clk_i) );
  dff prod2_reg_2__2__15_ ( .Q(larray[255]), .D(n6199), .CLK(clk_i) );
  dff prod2_reg_2__2__14_ ( .Q(larray[254]), .D(n6223), .CLK(clk_i) );
  dff prod2_reg_2__2__13_ ( .Q(larray[253]), .D(n6257), .CLK(clk_i) );
  dff prod2_reg_2__2__12_ ( .Q(larray[252]), .D(n6204), .CLK(clk_i) );
  dff prod2_reg_2__2__11_ ( .Q(larray[251]), .D(n4421), .CLK(clk_i) );
  dff prod2_reg_2__2__10_ ( .Q(larray[250]), .D(n6254), .CLK(clk_i) );
  dff prod2_reg_2__2__9_ ( .Q(larray[249]), .D(n6229), .CLK(clk_i) );
  dff prod2_reg_2__2__8_ ( .Q(larray[248]), .D(n6165), .CLK(clk_i) );
  dff prod2_reg_2__2__7_ ( .Q(larray[247]), .D(n6139), .CLK(clk_i) );
  dff prod2_reg_2__2__6_ ( .Q(larray[246]), .D(n6267), .CLK(clk_i) );
  dff prod2_reg_2__2__5_ ( .Q(larray[245]), .D(n5662), .CLK(clk_i) );
  dff prod2_reg_2__2__4_ ( .Q(larray[244]), .D(n5672), .CLK(clk_i) );
  dff prod2_reg_2__2__3_ ( .Q(larray[243]), .D(n5792), .CLK(clk_i) );
  dff prod2_reg_2__2__2_ ( .Q(larray[242]), .D(n5628), .CLK(clk_i) );
  dff prod2_reg_2__2__1_ ( .Q(larray[241]), .D(n5680), .CLK(clk_i) );
  dff prod2_reg_2__2__0_ ( .Q(larray[240]), .D(n5744), .CLK(clk_i) );
  dff prod2_reg_2__1__23_ ( .Q(larray[239]), .D(n5630), .CLK(clk_i) );
  dff prod2_reg_2__1__22_ ( .Q(larray[238]), .D(n5622), .CLK(clk_i) );
  dff prod2_reg_2__1__21_ ( .Q(larray[237]), .D(n5746), .CLK(clk_i) );
  dff prod2_reg_2__1__20_ ( .Q(larray[236]), .D(n5664), .CLK(clk_i) );
  dff prod2_reg_2__1__19_ ( .Q(larray[235]), .D(n5656), .CLK(clk_i) );
  dff prod2_reg_2__1__18_ ( .Q(larray[234]), .D(n5774), .CLK(clk_i) );
  dff prod2_reg_2__1__17_ ( .Q(larray[233]), .D(n6145), .CLK(clk_i) );
  dff prod2_reg_2__1__16_ ( .Q(larray[232]), .D(n6238), .CLK(clk_i) );
  dff prod2_reg_2__1__15_ ( .Q(larray[231]), .D(n6208), .CLK(clk_i) );
  dff prod2_reg_2__1__14_ ( .Q(larray[230]), .D(n6237), .CLK(clk_i) );
  dff prod2_reg_2__1__13_ ( .Q(larray[229]), .D(n6255), .CLK(clk_i) );
  dff prod2_reg_2__1__12_ ( .Q(larray[228]), .D(n6253), .CLK(clk_i) );
  dff prod2_reg_2__1__11_ ( .Q(larray[227]), .D(n6233), .CLK(clk_i) );
  dff prod2_reg_2__1__10_ ( .Q(larray[226]), .D(n6246), .CLK(clk_i) );
  dff prod2_reg_2__1__9_ ( .Q(larray[225]), .D(n6187), .CLK(clk_i) );
  dff prod2_reg_2__1__8_ ( .Q(larray[224]), .D(n4448), .CLK(clk_i) );
  dff prod2_reg_2__1__7_ ( .Q(larray[223]), .D(n6142), .CLK(clk_i) );
  dff prod2_reg_2__1__6_ ( .Q(larray[222]), .D(n6273), .CLK(clk_i) );
  dff prod2_reg_2__1__5_ ( .Q(larray[221]), .D(n5644), .CLK(clk_i) );
  dff prod2_reg_2__1__4_ ( .Q(larray[220]), .D(n5642), .CLK(clk_i) );
  dff prod2_reg_2__1__3_ ( .Q(larray[219]), .D(n5790), .CLK(clk_i) );
  dff prod2_reg_2__1__2_ ( .Q(larray[218]), .D(n5618), .CLK(clk_i) );
  dff prod2_reg_2__1__1_ ( .Q(larray[217]), .D(n5624), .CLK(clk_i) );
  dff prod2_reg_2__1__0_ ( .Q(larray[216]), .D(n5778), .CLK(clk_i) );
  dff prod2_reg_2__0__23_ ( .Q(larray[215]), .D(n6157), .CLK(clk_i) );
  dff prod2_reg_2__0__22_ ( .Q(larray[214]), .D(n6235), .CLK(clk_i) );
  dff prod2_reg_2__0__21_ ( .Q(larray[213]), .D(n6206), .CLK(clk_i) );
  dff prod2_reg_2__0__20_ ( .Q(larray[212]), .D(n6202), .CLK(clk_i) );
  dff prod2_reg_2__0__19_ ( .Q(larray[211]), .D(n6248), .CLK(clk_i) );
  dff prod2_reg_2__0__18_ ( .Q(larray[210]), .D(n6203), .CLK(clk_i) );
  dff prod2_reg_2__0__17_ ( .Q(larray[209]), .D(n4463), .CLK(clk_i) );
  dff prod2_reg_2__0__16_ ( .Q(larray[208]), .D(n6249), .CLK(clk_i) );
  dff prod2_reg_2__0__15_ ( .Q(larray[207]), .D(n6168), .CLK(clk_i) );
  dff prod2_reg_2__0__14_ ( .Q(larray[206]), .D(n6183), .CLK(clk_i) );
  dff prod2_reg_2__0__13_ ( .Q(larray[205]), .D(n6140), .CLK(clk_i) );
  dff prod2_reg_2__0__12_ ( .Q(larray[204]), .D(n6275), .CLK(clk_i) );
  dff prod2_reg_2__0__11_ ( .Q(larray[203]), .D(n5616), .CLK(clk_i) );
  dff prod2_reg_2__0__10_ ( .Q(larray[202]), .D(n5676), .CLK(clk_i) );
  dff prod2_reg_2__0__9_ ( .Q(larray[201]), .D(n5748), .CLK(clk_i) );
  dff prod2_reg_2__0__8_ ( .Q(larray[200]), .D(n5620), .CLK(clk_i) );
  dff prod2_reg_2__0__7_ ( .Q(larray[199]), .D(n5638), .CLK(clk_i) );
  dff prod2_reg_2__0__6_ ( .Q(larray[198]), .D(n5762), .CLK(clk_i) );
  dff prod2_reg_2__0__5_ ( .Q(larray[197]), .D(n5646), .CLK(clk_i) );
  dff prod2_reg_2__0__4_ ( .Q(larray[196]), .D(n5636), .CLK(clk_i) );
  dff prod2_reg_2__0__3_ ( .Q(larray[195]), .D(n5788), .CLK(clk_i) );
  dff prod2_reg_2__0__2_ ( .Q(larray[194]), .D(n5666), .CLK(clk_i) );
  dff prod2_reg_2__0__1_ ( .Q(larray[193]), .D(n5658), .CLK(clk_i) );
  dff prod2_reg_2__0__0_ ( .Q(larray[192]), .D(n5786), .CLK(clk_i) );
  dff prod2_reg_1__3__23_ ( .Q(larray[191]), .D(n5824), .CLK(clk_i) );
  dff prod2_reg_1__3__22_ ( .Q(larray[190]), .D(n5892), .CLK(clk_i) );
  dff prod2_reg_1__3__21_ ( .Q(larray[189]), .D(n5922), .CLK(clk_i) );
  dff prod2_reg_1__3__20_ ( .Q(larray[188]), .D(n5930), .CLK(clk_i) );
  dff prod2_reg_1__3__19_ ( .Q(larray[187]), .D(n5820), .CLK(clk_i) );
  dff prod2_reg_1__3__18_ ( .Q(larray[186]), .D(n5826), .CLK(clk_i) );
  dff prod2_reg_1__3__17_ ( .Q(larray[185]), .D(n5854), .CLK(clk_i) );
  dff prod2_reg_1__3__16_ ( .Q(larray[184]), .D(n5836), .CLK(clk_i) );
  dff prod2_reg_1__3__15_ ( .Q(larray[183]), .D(n5914), .CLK(clk_i) );
  dff prod2_reg_1__3__14_ ( .Q(larray[182]), .D(n5852), .CLK(clk_i) );
  dff prod2_reg_1__3__13_ ( .Q(larray[181]), .D(n5880), .CLK(clk_i) );
  dff prod2_reg_1__3__12_ ( .Q(larray[180]), .D(n5886), .CLK(clk_i) );
  dff prod2_reg_1__3__11_ ( .Q(larray[179]), .D(n4493), .CLK(clk_i) );
  dff prod2_reg_1__3__10_ ( .Q(larray[178]), .D(n4494), .CLK(clk_i) );
  dff prod2_reg_1__3__9_ ( .Q(larray[177]), .D(n4495), .CLK(clk_i) );
  dff prod2_reg_1__3__8_ ( .Q(larray[176]), .D(n4496), .CLK(clk_i) );
  dff prod2_reg_1__3__7_ ( .Q(larray[175]), .D(n4497), .CLK(clk_i) );
  dff prod2_reg_1__3__6_ ( .Q(larray[174]), .D(n4498), .CLK(clk_i) );
  dff prod2_reg_1__3__5_ ( .Q(larray[173]), .D(n4499), .CLK(clk_i) );
  dff prod2_reg_1__3__4_ ( .Q(larray[172]), .D(n4500), .CLK(clk_i) );
  dff prod2_reg_1__3__3_ ( .Q(larray[171]), .D(n4501), .CLK(clk_i) );
  dff prod2_reg_1__3__2_ ( .Q(larray[170]), .D(n4502), .CLK(clk_i) );
  dff prod2_reg_1__3__1_ ( .Q(larray[169]), .D(n4503), .CLK(clk_i) );
  dff prod2_reg_1__3__0_ ( .Q(larray[168]), .D(n4504), .CLK(clk_i) );
  dff prod2_reg_1__2__23_ ( .Q(larray[167]), .D(n5862), .CLK(clk_i) );
  dff prod2_reg_1__2__22_ ( .Q(larray[166]), .D(n5884), .CLK(clk_i) );
  dff prod2_reg_1__2__21_ ( .Q(larray[165]), .D(n5860), .CLK(clk_i) );
  dff prod2_reg_1__2__20_ ( .Q(larray[164]), .D(n5916), .CLK(clk_i) );
  dff prod2_reg_1__2__19_ ( .Q(larray[163]), .D(n5832), .CLK(clk_i) );
  dff prod2_reg_1__2__18_ ( .Q(larray[162]), .D(n5838), .CLK(clk_i) );
  dff prod2_reg_1__2__17_ ( .Q(larray[161]), .D(n4511), .CLK(clk_i) );
  dff prod2_reg_1__2__16_ ( .Q(larray[160]), .D(n4512), .CLK(clk_i) );
  dff prod2_reg_1__2__15_ ( .Q(larray[159]), .D(n4513), .CLK(clk_i) );
  dff prod2_reg_1__2__14_ ( .Q(larray[158]), .D(n4514), .CLK(clk_i) );
  dff prod2_reg_1__2__13_ ( .Q(larray[157]), .D(n4515), .CLK(clk_i) );
  dff prod2_reg_1__2__12_ ( .Q(larray[156]), .D(n4516), .CLK(clk_i) );
  dff prod2_reg_1__2__11_ ( .Q(larray[155]), .D(n4517), .CLK(clk_i) );
  dff prod2_reg_1__2__10_ ( .Q(larray[154]), .D(n4518), .CLK(clk_i) );
  dff prod2_reg_1__2__9_ ( .Q(larray[153]), .D(n4519), .CLK(clk_i) );
  dff prod2_reg_1__2__8_ ( .Q(larray[152]), .D(n4520), .CLK(clk_i) );
  dff prod2_reg_1__2__7_ ( .Q(larray[151]), .D(n4521), .CLK(clk_i) );
  dff prod2_reg_1__2__6_ ( .Q(larray[150]), .D(n4522), .CLK(clk_i) );
  dff prod2_reg_1__2__5_ ( .Q(larray[149]), .D(n5822), .CLK(clk_i) );
  dff prod2_reg_1__2__4_ ( .Q(larray[148]), .D(n5896), .CLK(clk_i) );
  dff prod2_reg_1__2__3_ ( .Q(larray[147]), .D(n5918), .CLK(clk_i) );
  dff prod2_reg_1__2__2_ ( .Q(larray[146]), .D(n5890), .CLK(clk_i) );
  dff prod2_reg_1__2__1_ ( .Q(larray[145]), .D(n5878), .CLK(clk_i) );
  dff prod2_reg_1__2__0_ ( .Q(larray[144]), .D(n5894), .CLK(clk_i) );
  dff prod2_reg_1__1__23_ ( .Q(larray[143]), .D(n5926), .CLK(clk_i) );
  dff prod2_reg_1__1__22_ ( .Q(larray[142]), .D(n5814), .CLK(clk_i) );
  dff prod2_reg_1__1__21_ ( .Q(larray[141]), .D(n5810), .CLK(clk_i) );
  dff prod2_reg_1__1__20_ ( .Q(larray[140]), .D(n5840), .CLK(clk_i) );
  dff prod2_reg_1__1__19_ ( .Q(larray[139]), .D(n5858), .CLK(clk_i) );
  dff prod2_reg_1__1__18_ ( .Q(larray[138]), .D(n5844), .CLK(clk_i) );
  dff prod2_reg_1__1__17_ ( .Q(larray[137]), .D(n4535), .CLK(clk_i) );
  dff prod2_reg_1__1__16_ ( .Q(larray[136]), .D(n4536), .CLK(clk_i) );
  dff prod2_reg_1__1__15_ ( .Q(larray[135]), .D(n4537), .CLK(clk_i) );
  dff prod2_reg_1__1__14_ ( .Q(larray[134]), .D(n4538), .CLK(clk_i) );
  dff prod2_reg_1__1__13_ ( .Q(larray[133]), .D(n4539), .CLK(clk_i) );
  dff prod2_reg_1__1__12_ ( .Q(larray[132]), .D(n4540), .CLK(clk_i) );
  dff prod2_reg_1__1__11_ ( .Q(larray[131]), .D(n4541), .CLK(clk_i) );
  dff prod2_reg_1__1__10_ ( .Q(larray[130]), .D(n4542), .CLK(clk_i) );
  dff prod2_reg_1__1__9_ ( .Q(larray[129]), .D(n4543), .CLK(clk_i) );
  dff prod2_reg_1__1__8_ ( .Q(larray[128]), .D(n4544), .CLK(clk_i) );
  dff prod2_reg_1__1__7_ ( .Q(larray[127]), .D(n4545), .CLK(clk_i) );
  dff prod2_reg_1__1__6_ ( .Q(larray[126]), .D(n4546), .CLK(clk_i) );
  dff prod2_reg_1__1__5_ ( .Q(larray[125]), .D(n5932), .CLK(clk_i) );
  dff prod2_reg_1__1__4_ ( .Q(larray[124]), .D(n5920), .CLK(clk_i) );
  dff prod2_reg_1__1__3_ ( .Q(larray[123]), .D(n5924), .CLK(clk_i) );
  dff prod2_reg_1__1__2_ ( .Q(larray[122]), .D(n5830), .CLK(clk_i) );
  dff prod2_reg_1__1__1_ ( .Q(larray[121]), .D(n5828), .CLK(clk_i) );
  dff prod2_reg_1__1__0_ ( .Q(larray[120]), .D(n5848), .CLK(clk_i) );
  dff prod2_reg_1__0__23_ ( .Q(larray[119]), .D(n4553), .CLK(clk_i) );
  dff prod2_reg_1__0__22_ ( .Q(larray[118]), .D(n4554), .CLK(clk_i) );
  dff prod2_reg_1__0__21_ ( .Q(larray[117]), .D(n4555), .CLK(clk_i) );
  dff prod2_reg_1__0__20_ ( .Q(larray[116]), .D(n4556), .CLK(clk_i) );
  dff prod2_reg_1__0__19_ ( .Q(larray[115]), .D(n4557), .CLK(clk_i) );
  dff prod2_reg_1__0__18_ ( .Q(larray[114]), .D(n4558), .CLK(clk_i) );
  dff prod2_reg_1__0__17_ ( .Q(larray[113]), .D(n4559), .CLK(clk_i) );
  dff prod2_reg_1__0__16_ ( .Q(larray[112]), .D(n4560), .CLK(clk_i) );
  dff prod2_reg_1__0__15_ ( .Q(larray[111]), .D(n4561), .CLK(clk_i) );
  dff prod2_reg_1__0__14_ ( .Q(larray[110]), .D(n4562), .CLK(clk_i) );
  dff prod2_reg_1__0__13_ ( .Q(larray[109]), .D(n4563), .CLK(clk_i) );
  dff prod2_reg_1__0__12_ ( .Q(larray[108]), .D(n4564), .CLK(clk_i) );
  dff prod2_reg_1__0__11_ ( .Q(larray[107]), .D(n5812), .CLK(clk_i) );
  dff prod2_reg_1__0__10_ ( .Q(larray[106]), .D(n5816), .CLK(clk_i) );
  dff prod2_reg_1__0__9_ ( .Q(larray[105]), .D(n5882), .CLK(clk_i) );
  dff prod2_reg_1__0__8_ ( .Q(larray[104]), .D(n5850), .CLK(clk_i) );
  dff prod2_reg_1__0__7_ ( .Q(larray[103]), .D(n5888), .CLK(clk_i) );
  dff prod2_reg_1__0__6_ ( .Q(larray[102]), .D(n5934), .CLK(clk_i) );
  dff prod2_reg_1__0__5_ ( .Q(larray[101]), .D(n5856), .CLK(clk_i) );
  dff prod2_reg_1__0__4_ ( .Q(larray[100]), .D(n5864), .CLK(clk_i) );
  dff prod2_reg_1__0__3_ ( .Q(larray[99]), .D(n5936), .CLK(clk_i) );
  dff prod2_reg_1__0__2_ ( .Q(larray[98]), .D(n5928), .CLK(clk_i) );
  dff prod2_reg_1__0__1_ ( .Q(larray[97]), .D(n5818), .CLK(clk_i) );
  dff prod2_reg_1__0__0_ ( .Q(larray[96]), .D(n5846), .CLK(clk_i) );
  dff prod2_reg_0__3__23_ ( .Q(larray[95]), .D(n5742), .CLK(clk_i) );
  dff prod2_reg_0__3__22_ ( .Q(larray[94]), .D(n5784), .CLK(clk_i) );
  dff prod2_reg_0__3__21_ ( .Q(larray[93]), .D(n5684), .CLK(clk_i) );
  dff prod2_reg_0__3__20_ ( .Q(larray[92]), .D(n5732), .CLK(clk_i) );
  dff prod2_reg_0__3__19_ ( .Q(larray[91]), .D(n5798), .CLK(clk_i) );
  dff prod2_reg_0__3__18_ ( .Q(larray[90]), .D(n5702), .CLK(clk_i) );
  dff prod2_reg_0__3__17_ ( .Q(larray[89]), .D(n5736), .CLK(clk_i) );
  dff prod2_reg_0__3__16_ ( .Q(larray[88]), .D(n5806), .CLK(clk_i) );
  dff prod2_reg_0__3__15_ ( .Q(larray[87]), .D(n5690), .CLK(clk_i) );
  dff prod2_reg_0__3__14_ ( .Q(larray[86]), .D(n5716), .CLK(clk_i) );
  dff prod2_reg_0__3__13_ ( .Q(larray[85]), .D(n5780), .CLK(clk_i) );
  dff prod2_reg_0__3__12_ ( .Q(larray[84]), .D(n5698), .CLK(clk_i) );
  dff prod2_reg_0__3__11_ ( .Q(larray[83]), .D(n4589), .CLK(clk_i) );
  dff prod2_reg_0__3__10_ ( .Q(larray[82]), .D(n4590), .CLK(clk_i) );
  dff prod2_reg_0__3__9_ ( .Q(larray[81]), .D(n4591), .CLK(clk_i) );
  dff prod2_reg_0__3__8_ ( .Q(larray[80]), .D(n4592), .CLK(clk_i) );
  dff prod2_reg_0__3__7_ ( .Q(larray[79]), .D(n4593), .CLK(clk_i) );
  dff prod2_reg_0__3__6_ ( .Q(larray[78]), .D(n4594), .CLK(clk_i) );
  dff prod2_reg_0__3__5_ ( .Q(larray[77]), .D(n4595), .CLK(clk_i) );
  dff prod2_reg_0__3__4_ ( .Q(larray[76]), .D(n4596), .CLK(clk_i) );
  dff prod2_reg_0__3__3_ ( .Q(larray[75]), .D(n4597), .CLK(clk_i) );
  dff prod2_reg_0__3__2_ ( .Q(larray[74]), .D(n4598), .CLK(clk_i) );
  dff prod2_reg_0__3__1_ ( .Q(larray[73]), .D(n4599), .CLK(clk_i) );
  dff prod2_reg_0__3__0_ ( .Q(larray[72]), .D(n4600), .CLK(clk_i) );
  dff prod2_reg_0__2__23_ ( .Q(larray[71]), .D(n5718), .CLK(clk_i) );
  dff prod2_reg_0__2__22_ ( .Q(larray[70]), .D(n5794), .CLK(clk_i) );
  dff prod2_reg_0__2__21_ ( .Q(larray[69]), .D(n5670), .CLK(clk_i) );
  dff prod2_reg_0__2__20_ ( .Q(larray[68]), .D(n5740), .CLK(clk_i) );
  dff prod2_reg_0__2__19_ ( .Q(larray[67]), .D(n5796), .CLK(clk_i) );
  dff prod2_reg_0__2__18_ ( .Q(larray[66]), .D(n5696), .CLK(clk_i) );
  dff prod2_reg_0__2__17_ ( .Q(larray[65]), .D(n4607), .CLK(clk_i) );
  dff prod2_reg_0__2__16_ ( .Q(larray[64]), .D(n4608), .CLK(clk_i) );
  dff prod2_reg_0__2__15_ ( .Q(larray[63]), .D(n4609), .CLK(clk_i) );
  dff prod2_reg_0__2__14_ ( .Q(larray[62]), .D(n4610), .CLK(clk_i) );
  dff prod2_reg_0__2__13_ ( .Q(larray[61]), .D(n4611), .CLK(clk_i) );
  dff prod2_reg_0__2__12_ ( .Q(larray[60]), .D(n4612), .CLK(clk_i) );
  dff prod2_reg_0__2__11_ ( .Q(larray[59]), .D(n4613), .CLK(clk_i) );
  dff prod2_reg_0__2__10_ ( .Q(larray[58]), .D(n4614), .CLK(clk_i) );
  dff prod2_reg_0__2__9_ ( .Q(larray[57]), .D(n4615), .CLK(clk_i) );
  dff prod2_reg_0__2__8_ ( .Q(larray[56]), .D(n4616), .CLK(clk_i) );
  dff prod2_reg_0__2__7_ ( .Q(larray[55]), .D(n4617), .CLK(clk_i) );
  dff prod2_reg_0__2__6_ ( .Q(larray[54]), .D(n4618), .CLK(clk_i) );
  dff prod2_reg_0__2__5_ ( .Q(larray[53]), .D(n5720), .CLK(clk_i) );
  dff prod2_reg_0__2__4_ ( .Q(larray[52]), .D(n5768), .CLK(clk_i) );
  dff prod2_reg_0__2__3_ ( .Q(larray[51]), .D(n5686), .CLK(clk_i) );
  dff prod2_reg_0__2__2_ ( .Q(larray[50]), .D(n5724), .CLK(clk_i) );
  dff prod2_reg_0__2__1_ ( .Q(larray[49]), .D(n5766), .CLK(clk_i) );
  dff prod2_reg_0__2__0_ ( .Q(larray[48]), .D(n5708), .CLK(clk_i) );
  dff prod2_reg_0__1__23_ ( .Q(larray[47]), .D(n5712), .CLK(clk_i) );
  dff prod2_reg_0__1__22_ ( .Q(larray[46]), .D(n5782), .CLK(clk_i) );
  dff prod2_reg_0__1__21_ ( .Q(larray[45]), .D(n5710), .CLK(clk_i) );
  dff prod2_reg_0__1__20_ ( .Q(larray[44]), .D(n5728), .CLK(clk_i) );
  dff prod2_reg_0__1__19_ ( .Q(larray[43]), .D(n5800), .CLK(clk_i) );
  dff prod2_reg_0__1__18_ ( .Q(larray[42]), .D(n5704), .CLK(clk_i) );
  dff prod2_reg_0__1__17_ ( .Q(larray[41]), .D(n4631), .CLK(clk_i) );
  dff prod2_reg_0__1__16_ ( .Q(larray[40]), .D(n4632), .CLK(clk_i) );
  dff prod2_reg_0__1__15_ ( .Q(larray[39]), .D(n4633), .CLK(clk_i) );
  dff prod2_reg_0__1__14_ ( .Q(larray[38]), .D(n4634), .CLK(clk_i) );
  dff prod2_reg_0__1__13_ ( .Q(larray[37]), .D(n4635), .CLK(clk_i) );
  dff prod2_reg_0__1__12_ ( .Q(larray[36]), .D(n4636), .CLK(clk_i) );
  dff prod2_reg_0__1__11_ ( .Q(larray[35]), .D(n4637), .CLK(clk_i) );
  dff prod2_reg_0__1__10_ ( .Q(larray[34]), .D(n4638), .CLK(clk_i) );
  dff prod2_reg_0__1__9_ ( .Q(larray[33]), .D(n4639), .CLK(clk_i) );
  dff prod2_reg_0__1__8_ ( .Q(larray[32]), .D(n4640), .CLK(clk_i) );
  dff prod2_reg_0__1__7_ ( .Q(larray[31]), .D(n4641), .CLK(clk_i) );
  dff prod2_reg_0__1__6_ ( .Q(larray[30]), .D(n4642), .CLK(clk_i) );
  dff prod2_reg_0__1__5_ ( .Q(larray[29]), .D(n5726), .CLK(clk_i) );
  dff prod2_reg_0__1__4_ ( .Q(larray[28]), .D(n5754), .CLK(clk_i) );
  dff prod2_reg_0__1__3_ ( .Q(larray[27]), .D(n5700), .CLK(clk_i) );
  dff prod2_reg_0__1__2_ ( .Q(larray[26]), .D(n5722), .CLK(clk_i) );
  dff prod2_reg_0__1__1_ ( .Q(larray[25]), .D(n5756), .CLK(clk_i) );
  dff prod2_reg_0__1__0_ ( .Q(larray[24]), .D(n5706), .CLK(clk_i) );
  dff prod2_reg_0__0__23_ ( .Q(larray[23]), .D(n4649), .CLK(clk_i) );
  dff prod2_reg_0__0__22_ ( .Q(larray[22]), .D(n4650), .CLK(clk_i) );
  dff prod2_reg_0__0__21_ ( .Q(larray[21]), .D(n4651), .CLK(clk_i) );
  dff prod2_reg_0__0__20_ ( .Q(larray[20]), .D(n4652), .CLK(clk_i) );
  dff prod2_reg_0__0__19_ ( .Q(larray[19]), .D(n4653), .CLK(clk_i) );
  dff prod2_reg_0__0__18_ ( .Q(larray[18]), .D(n4654), .CLK(clk_i) );
  dff prod2_reg_0__0__17_ ( .Q(larray[17]), .D(n4655), .CLK(clk_i) );
  dff prod2_reg_0__0__16_ ( .Q(larray[16]), .D(n4656), .CLK(clk_i) );
  dff prod2_reg_0__0__15_ ( .Q(larray[15]), .D(n4657), .CLK(clk_i) );
  dff prod2_reg_0__0__14_ ( .Q(larray[14]), .D(n4658), .CLK(clk_i) );
  dff prod2_reg_0__0__13_ ( .Q(larray[13]), .D(n4659), .CLK(clk_i) );
  dff prod2_reg_0__0__12_ ( .Q(larray[12]), .D(n4660), .CLK(clk_i) );
  dff prod2_reg_0__0__11_ ( .Q(larray[11]), .D(n5730), .CLK(clk_i) );
  dff prod2_reg_0__0__10_ ( .Q(larray[10]), .D(n5804), .CLK(clk_i) );
  dff prod2_reg_0__0__9_ ( .Q(larray[9]), .D(n5688), .CLK(clk_i) );
  dff prod2_reg_0__0__8_ ( .Q(larray[8]), .D(n5734), .CLK(clk_i) );
  dff prod2_reg_0__0__7_ ( .Q(larray[7]), .D(n5770), .CLK(clk_i) );
  dff prod2_reg_0__0__6_ ( .Q(larray[6]), .D(n5668), .CLK(clk_i) );
  dff prod2_reg_0__0__5_ ( .Q(larray[5]), .D(n5714), .CLK(clk_i) );
  dff prod2_reg_0__0__4_ ( .Q(larray[4]), .D(n5752), .CLK(clk_i) );
  dff prod2_reg_0__0__3_ ( .Q(larray[3]), .D(n5692), .CLK(clk_i) );
  dff prod2_reg_0__0__2_ ( .Q(larray[2]), .D(n5738), .CLK(clk_i) );
  dff prod2_reg_0__0__1_ ( .Q(larray[1]), .D(n5802), .CLK(clk_i) );
  dff prod2_reg_0__0__0_ ( .Q(larray[0]), .D(n5694), .CLK(clk_i) );
  dff sum_reg_3__23_ ( .Q(prod_a_b_3__23_), .QB(n4277), .D(n6128), .CLK(clk_i)
         );
  dff sum_reg_3__22_ ( .Q(prod_a_b_3__22_), .QB(n4276), .D(n4674), .CLK(clk_i)
         );
  dff sum_reg_3__21_ ( .Q(prod_a_b_3__21_), .QB(n4275), .D(n6064), .CLK(clk_i)
         );
  dff sum_reg_3__20_ ( .Q(prod_a_b_3__20_), .QB(n4274), .D(n6040), .CLK(clk_i)
         );
  dff sum_reg_3__19_ ( .Q(prod_a_b_3__19_), .QB(n4272), .D(n6025), .CLK(clk_i)
         );
  dff sum_reg_3__18_ ( .Q(prod_a_b_3__18_), .QB(n4271), .D(n6076), .CLK(clk_i)
         );
  dff sum_reg_3__17_ ( .Q(prod_a_b_3__17_), .QB(n4270), .D(n6093), .CLK(clk_i)
         );
  dff sum_reg_3__16_ ( .Q(prod_a_b_3__16_), .QB(n4269), .D(n6104), .CLK(clk_i)
         );
  dff sum_reg_3__15_ ( .Q(prod_a_b_3__15_), .QB(n4268), .D(n6062), .CLK(clk_i)
         );
  dff sum_reg_3__14_ ( .Q(prod_a_b_3__14_), .QB(n4267), .D(n6105), .CLK(clk_i)
         );
  dff sum_reg_3__13_ ( .Q(prod_a_b_3__13_), .QB(n4266), .D(n6108), .CLK(clk_i)
         );
  dff sum_reg_3__12_ ( .Q(prod_a_b_3__12_), .QB(n4265), .D(n6051), .CLK(clk_i)
         );
  dff sum_reg_3__11_ ( .Q(prod_a_b_3__11_), .QB(n4264), .D(n6112), .CLK(clk_i)
         );
  dff sum_reg_3__10_ ( .Q(prod_a_b_3__10_), .QB(n4263), .D(n6082), .CLK(clk_i)
         );
  dff sum_reg_3__9_ ( .Q(prod_a_b_3__9_), .QB(n4285), .D(n6091), .CLK(clk_i)
         );
  dff sum_reg_3__8_ ( .Q(prod_a_b_3__8_), .QB(n4284), .D(n6069), .CLK(clk_i)
         );
  dff sum_reg_3__7_ ( .Q(prod_a_b_3__7_), .QB(n4283), .D(n6114), .CLK(clk_i)
         );
  dff sum_reg_3__6_ ( .Q(prod_a_b_3__6_), .QB(n4282), .D(n6075), .CLK(clk_i)
         );
  dff sum_reg_3__5_ ( .Q(prod_a_b_3__5_), .QB(n4281), .D(n6036), .CLK(clk_i)
         );
  dff sum_reg_3__4_ ( .Q(prod_a_b_3__4_), .QB(n4280), .D(n6023), .CLK(clk_i)
         );
  dff sum_reg_3__3_ ( .Q(prod_a_b_3__3_), .QB(n4279), .D(n6016), .CLK(clk_i)
         );
  dff sum_reg_3__2_ ( .Q(prod_a_b_3__2_), .QB(n4278), .D(n6101), .CLK(clk_i)
         );
  dff sum_reg_3__1_ ( .Q(prod_a_b_3__1_), .QB(n4273), .D(n6109), .CLK(clk_i)
         );
  dff sum_reg_3__0_ ( .Q(prod_a_b_3__0_), .QB(n4262), .D(n4696), .CLK(clk_i)
         );
  dff sum_reg_2__23_ ( .Q(prod_a_b_2__35_), .QB(n4253), .D(n4697), .CLK(clk_i)
         );
  dff sum_reg_2__22_ ( .Q(prod_a_b_2__34_), .QB(n4252), .D(n6134), .CLK(clk_i)
         );
  dff sum_reg_2__21_ ( .Q(prod_a_b_2__33_), .QB(n4251), .D(n6037), .CLK(clk_i)
         );
  dff sum_reg_2__20_ ( .Q(prod_a_b_2__32_), .QB(n4250), .D(n6038), .CLK(clk_i)
         );
  dff sum_reg_2__19_ ( .Q(prod_a_b_2__31_), .QB(n4248), .D(n6096), .CLK(clk_i)
         );
  dff sum_reg_2__18_ ( .Q(prod_a_b_2__30_), .QB(n4247), .D(n6033), .CLK(clk_i)
         );
  dff sum_reg_2__17_ ( .Q(prod_a_b_2__29_), .QB(n4246), .D(n6039), .CLK(clk_i)
         );
  dff sum_reg_2__16_ ( .Q(prod_a_b_2__28_), .QB(n4245), .D(n6098), .CLK(clk_i)
         );
  dff sum_reg_2__15_ ( .Q(prod_a_b_2__27_), .QB(n4244), .D(n6032), .CLK(clk_i)
         );
  dff sum_reg_2__14_ ( .Q(prod_a_b_2__26_), .QB(n4243), .D(n6063), .CLK(clk_i)
         );
  dff sum_reg_2__13_ ( .Q(prod_a_b_2__25_), .QB(n4242), .D(n6024), .CLK(clk_i)
         );
  dff sum_reg_2__12_ ( .Q(prod_a_b_2__24_), .QB(n4241), .D(n4708), .CLK(clk_i)
         );
  dff sum_reg_2__11_ ( .Q(prod_a_b_2__23_), .QB(n4240), .D(n6073), .CLK(clk_i)
         );
  dff sum_reg_2__10_ ( .Q(prod_a_b_2__22_), .QB(n4239), .D(n6089), .CLK(clk_i)
         );
  dff sum_reg_2__9_ ( .Q(prod_a_b_2__21_), .QB(n4261), .D(n6066), .CLK(clk_i)
         );
  dff sum_reg_2__8_ ( .Q(prod_a_b_2__20_), .QB(n4260), .D(n6065), .CLK(clk_i)
         );
  dff sum_reg_2__7_ ( .Q(prod_a_b_2__19_), .QB(n4259), .D(n6058), .CLK(clk_i)
         );
  dff sum_reg_2__6_ ( .Q(prod_a_b_2__18_), .QB(n4258), .D(n6077), .CLK(clk_i)
         );
  dff sum_reg_2__5_ ( .Q(prod_a_b_2__17_), .QB(n4257), .D(n6092), .CLK(clk_i)
         );
  dff sum_reg_2__4_ ( .Q(prod_a_b_2__16_), .QB(n4256), .D(n6068), .CLK(clk_i)
         );
  dff sum_reg_2__3_ ( .Q(prod_a_b_2__15_), .QB(n4255), .D(n4717), .CLK(clk_i)
         );
  dff sum_reg_2__2_ ( .Q(prod_a_b_2__14_), .QB(n4254), .D(n6110), .CLK(clk_i)
         );
  dff sum_reg_2__1_ ( .Q(prod_a_b_2__13_), .QB(n4249), .D(n6031), .CLK(clk_i)
         );
  dff sum_reg_2__0_ ( .Q(prod_a_b_2__12_), .QB(n4238), .D(n6011), .CLK(clk_i)
         );
  dff sum_reg_1__23_ ( .Q(prod_a_b_1__35_), .QB(n4229), .D(n6135), .CLK(clk_i)
         );
  dff sum_reg_1__22_ ( .Q(prod_a_b_1__34_), .QB(n4228), .D(n6022), .CLK(clk_i)
         );
  dff sum_reg_1__21_ ( .Q(prod_a_b_1__33_), .QB(n4227), .D(n6097), .CLK(clk_i)
         );
  dff sum_reg_1__20_ ( .Q(prod_a_b_1__32_), .QB(n4226), .D(n6106), .CLK(clk_i)
         );
  dff sum_reg_1__19_ ( .Q(prod_a_b_1__31_), .QB(n4224), .D(n6102), .CLK(clk_i)
         );
  dff sum_reg_1__18_ ( .Q(prod_a_b_1__30_), .QB(n4223), .D(n6081), .CLK(clk_i)
         );
  dff sum_reg_1__17_ ( .Q(prod_a_b_1__29_), .QB(n4222), .D(n6052), .CLK(clk_i)
         );
  dff sum_reg_1__16_ ( .Q(prod_a_b_1__28_), .QB(n4221), .D(n6115), .CLK(clk_i)
         );
  dff sum_reg_1__15_ ( .Q(prod_a_b_1__27_), .QB(n4220), .D(n6078), .CLK(clk_i)
         );
  dff sum_reg_1__14_ ( .Q(prod_a_b_1__26_), .QB(n4219), .D(n6044), .CLK(clk_i)
         );
  dff sum_reg_1__13_ ( .Q(prod_a_b_1__25_), .QB(n4218), .D(n6041), .CLK(clk_i)
         );
  dff sum_reg_1__12_ ( .Q(prod_a_b_1__24_), .QB(n4217), .D(n6116), .CLK(clk_i)
         );
  dff sum_reg_1__11_ ( .Q(prod_a_b_1__23_), .QB(n4216), .D(n6100), .CLK(clk_i)
         );
  dff sum_reg_1__10_ ( .Q(prod_a_b_1__22_), .QB(n4215), .D(n6061), .CLK(clk_i)
         );
  dff sum_reg_1__9_ ( .Q(prod_a_b_1__21_), .QB(n4237), .D(n6059), .CLK(clk_i)
         );
  dff sum_reg_1__8_ ( .Q(prod_a_b_1__20_), .QB(n4236), .D(n6054), .CLK(clk_i)
         );
  dff sum_reg_1__7_ ( .Q(prod_a_b_1__19_), .QB(n4235), .D(n6060), .CLK(clk_i)
         );
  dff sum_reg_1__6_ ( .Q(prod_a_b_1__18_), .QB(n4234), .D(n6034), .CLK(clk_i)
         );
  dff sum_reg_1__5_ ( .Q(prod_a_b_1__17_), .QB(n4233), .D(n6113), .CLK(clk_i)
         );
  dff sum_reg_1__4_ ( .Q(prod_a_b_1__16_), .QB(n4232), .D(n6053), .CLK(clk_i)
         );
  dff sum_reg_1__3_ ( .Q(prod_a_b_1__15_), .QB(n4231), .D(n6094), .CLK(clk_i)
         );
  dff sum_reg_1__2_ ( .Q(prod_a_b_1__14_), .QB(n4230), .D(n6071), .CLK(clk_i)
         );
  dff sum_reg_1__1_ ( .Q(prod_a_b_1__13_), .QB(n4225), .D(n6095), .CLK(clk_i)
         );
  dff sum_reg_1__0_ ( .Q(prod_a_b_1__12_), .QB(n4214), .D(n4744), .CLK(clk_i)
         );
  dff sum_reg_0__23_ ( .Q(prod_a_b_0__47_), .QB(n4205), .D(n4745), .CLK(clk_i)
         );
  dff sum_reg_0__22_ ( .Q(prod_a_b_0__46_), .QB(n4204), .D(n4746), .CLK(clk_i)
         );
  dff sum_reg_0__21_ ( .Q(prod_a_b_0__45_), .QB(n4203), .D(n6056), .CLK(clk_i)
         );
  dff sum_reg_0__20_ ( .Q(prod_a_b_0__44_), .QB(n4202), .D(n6070), .CLK(clk_i)
         );
  dff sum_reg_0__19_ ( .Q(prod_a_b_0__43_), .QB(n4200), .D(n6043), .CLK(clk_i)
         );
  dff sum_reg_0__18_ ( .Q(prod_a_b_0__42_), .QB(n4199), .D(n6072), .CLK(clk_i)
         );
  dff sum_reg_0__17_ ( .Q(prod_a_b_0__41_), .QB(n4198), .D(n6067), .CLK(clk_i)
         );
  dff sum_reg_0__16_ ( .Q(prod_a_b_0__40_), .QB(n4197), .D(n6042), .CLK(clk_i)
         );
  dff sum_reg_0__15_ ( .Q(prod_a_b_0__39_), .QB(n4196), .D(n6111), .CLK(clk_i)
         );
  dff sum_reg_0__14_ ( .Q(prod_a_b_0__38_), .QB(n4195), .D(n6080), .CLK(clk_i)
         );
  dff sum_reg_0__13_ ( .Q(prod_a_b_0__37_), .QB(n4194), .D(n6035), .CLK(clk_i)
         );
  dff sum_reg_0__12_ ( .Q(prod_a_b_0__36_), .QB(n4193), .D(n6079), .CLK(clk_i)
         );
  dff sum_reg_0__11_ ( .Q(prod_a_b_0__35_), .QB(n4192), .D(n6055), .CLK(clk_i)
         );
  dff sum_reg_0__10_ ( .Q(prod_a_b_0__34_), .QB(n4191), .D(n6117), .CLK(clk_i)
         );
  dff sum_reg_0__9_ ( .Q(prod_a_b_0__33_), .QB(n4213), .D(n6074), .CLK(clk_i)
         );
  dff sum_reg_0__8_ ( .Q(prod_a_b_0__32_), .QB(n4212), .D(n6099), .CLK(clk_i)
         );
  dff sum_reg_0__7_ ( .Q(prod_a_b_0__31_), .QB(n4211), .D(n6107), .CLK(clk_i)
         );
  dff sum_reg_0__6_ ( .Q(prod_a_b_0__30_), .QB(n4210), .D(n6103), .CLK(clk_i)
         );
  dff sum_reg_0__5_ ( .Q(prod_a_b_0__29_), .QB(n4209), .D(n6057), .CLK(clk_i)
         );
  dff sum_reg_0__4_ ( .Q(prod_a_b_0__28_), .QB(n4208), .D(n6083), .CLK(clk_i)
         );
  dff sum_reg_0__3_ ( .Q(prod_a_b_0__27_), .QB(n4207), .D(n6090), .CLK(clk_i)
         );
  dff sum_reg_0__2_ ( .Q(prod_a_b_0__26_), .QB(n4206), .D(n6045), .CLK(clk_i)
         );
  dff sum_reg_0__1_ ( .Q(prod_a_b_0__25_), .QB(n4201), .D(n4767), .CLK(clk_i)
         );
  dff sum_reg_0__0_ ( .Q(prod_a_b_0__24_), .QB(n4190), .D(n4768), .CLK(clk_i)
         );
  dff s_state_reg ( .Q(s_state), .D(n4769), .CLK(clk_i) );
  dff s_ready_o_reg ( .Q(ready_o), .QB(n4189), .D(n4770), .CLK(clk_i) );
  dff s_fracta_i_reg_23_ ( .QB(n3583), .D(fracta_i[23]), .CLK(clk_i) );
  dff s_fracta_i_reg_22_ ( .QB(n3582), .D(fracta_i[22]), .CLK(clk_i) );
  dff s_fracta_i_reg_21_ ( .QB(n3581), .D(fracta_i[21]), .CLK(clk_i) );
  dff s_fracta_i_reg_20_ ( .QB(n3580), .D(fracta_i[20]), .CLK(clk_i) );
  dff s_fracta_i_reg_19_ ( .QB(n3579), .D(fracta_i[19]), .CLK(clk_i) );
  dff s_fracta_i_reg_18_ ( .QB(n3578), .D(fracta_i[18]), .CLK(clk_i) );
  dff s_fracta_i_reg_17_ ( .QB(n3577), .D(fracta_i[17]), .CLK(clk_i) );
  dff s_fracta_i_reg_16_ ( .QB(n3576), .D(fracta_i[16]), .CLK(clk_i) );
  dff s_fracta_i_reg_15_ ( .QB(n3575), .D(fracta_i[15]), .CLK(clk_i) );
  dff s_fracta_i_reg_14_ ( .QB(n3574), .D(fracta_i[14]), .CLK(clk_i) );
  dff s_fracta_i_reg_13_ ( .QB(n3573), .D(fracta_i[13]), .CLK(clk_i) );
  dff s_fracta_i_reg_12_ ( .QB(n3572), .D(fracta_i[12]), .CLK(clk_i) );
  dff s_fracta_i_reg_11_ ( .QB(n3571), .D(fracta_i[11]), .CLK(clk_i) );
  dff s_fracta_i_reg_10_ ( .QB(n3570), .D(fracta_i[10]), .CLK(clk_i) );
  dff s_fracta_i_reg_9_ ( .QB(n3569), .D(fracta_i[9]), .CLK(clk_i) );
  dff s_fracta_i_reg_8_ ( .QB(n3568), .D(fracta_i[8]), .CLK(clk_i) );
  dff s_fracta_i_reg_7_ ( .QB(n3567), .D(fracta_i[7]), .CLK(clk_i) );
  dff s_fracta_i_reg_6_ ( .QB(n3566), .D(fracta_i[6]), .CLK(clk_i) );
  dff s_fracta_i_reg_5_ ( .QB(n3565), .D(fracta_i[5]), .CLK(clk_i) );
  dff s_fracta_i_reg_4_ ( .QB(n3564), .D(fracta_i[4]), .CLK(clk_i) );
  dff s_fracta_i_reg_3_ ( .QB(n3563), .D(fracta_i[3]), .CLK(clk_i) );
  dff s_fracta_i_reg_2_ ( .QB(n3562), .D(fracta_i[2]), .CLK(clk_i) );
  dff s_fracta_i_reg_1_ ( .QB(n3561), .D(fracta_i[1]), .CLK(clk_i) );
  dff s_fracta_i_reg_0_ ( .QB(n3560), .D(fracta_i[0]), .CLK(clk_i) );
  dff s_fractb_i_reg_23_ ( .QB(n3559), .D(fractb_i[23]), .CLK(clk_i) );
  dff s_fractb_i_reg_22_ ( .QB(n3558), .D(fractb_i[22]), .CLK(clk_i) );
  dff s_fractb_i_reg_21_ ( .QB(n3557), .D(fractb_i[21]), .CLK(clk_i) );
  dff s_fractb_i_reg_20_ ( .QB(n3556), .D(fractb_i[20]), .CLK(clk_i) );
  dff s_fractb_i_reg_19_ ( .QB(n3555), .D(fractb_i[19]), .CLK(clk_i) );
  dff s_fractb_i_reg_18_ ( .QB(n3554), .D(fractb_i[18]), .CLK(clk_i) );
  dff s_fractb_i_reg_17_ ( .QB(n3553), .D(fractb_i[17]), .CLK(clk_i) );
  dff s_fractb_i_reg_16_ ( .QB(n3552), .D(fractb_i[16]), .CLK(clk_i) );
  dff s_fractb_i_reg_15_ ( .QB(n3551), .D(fractb_i[15]), .CLK(clk_i) );
  dff s_fractb_i_reg_14_ ( .QB(n3550), .D(fractb_i[14]), .CLK(clk_i) );
  dff s_fractb_i_reg_13_ ( .QB(n3549), .D(fractb_i[13]), .CLK(clk_i) );
  dff s_fractb_i_reg_12_ ( .QB(n3548), .D(fractb_i[12]), .CLK(clk_i) );
  dff s_fractb_i_reg_11_ ( .QB(n3547), .D(fractb_i[11]), .CLK(clk_i) );
  dff s_fractb_i_reg_10_ ( .QB(n3546), .D(fractb_i[10]), .CLK(clk_i) );
  dff s_fractb_i_reg_9_ ( .QB(n3545), .D(fractb_i[9]), .CLK(clk_i) );
  dff s_fractb_i_reg_8_ ( .QB(n3544), .D(fractb_i[8]), .CLK(clk_i) );
  dff s_fractb_i_reg_7_ ( .QB(n3543), .D(fractb_i[7]), .CLK(clk_i) );
  dff s_fractb_i_reg_6_ ( .QB(n3542), .D(fractb_i[6]), .CLK(clk_i) );
  dff s_fractb_i_reg_5_ ( .QB(n3541), .D(fractb_i[5]), .CLK(clk_i) );
  dff s_fractb_i_reg_4_ ( .QB(n3540), .D(fractb_i[4]), .CLK(clk_i) );
  dff s_fractb_i_reg_3_ ( .QB(n3539), .D(fractb_i[3]), .CLK(clk_i) );
  dff s_fractb_i_reg_2_ ( .QB(n3538), .D(fractb_i[2]), .CLK(clk_i) );
  dff s_fractb_i_reg_1_ ( .QB(n3537), .D(fractb_i[1]), .CLK(clk_i) );
  dff s_fractb_i_reg_0_ ( .QB(n3536), .D(fractb_i[0]), .CLK(clk_i) );
  dff s_signa_i_reg ( .QB(n3535), .D(signa_i), .CLK(clk_i) );
  dff s_signb_i_reg ( .Q(s_signb_i), .D(signb_i), .CLK(clk_i) );
  dff s_start_i_reg ( .Q(s_state83), .D(start_i), .CLK(clk_i) );
  ao21 U1504 ( .Y(n4771), .A0(n6994), .A1(n6995), .B0(n4189) );
  inv01 U1505 ( .Y(n4772), .A(n4771) );
  inv02 U1506 ( .Y(n6994), .A(s_state83) );
  inv01 U1507 ( .Y(member996_4__2_), .A(n4773) );
  nor02 U1508 ( .Y(n4774), .A0(n6940), .A1(n7366) );
  nor02 U1509 ( .Y(n4775), .A0(n3562), .A1(n7366) );
  nor02 U1510 ( .Y(n4776), .A0(n6940), .A1(n3574) );
  nor02 U1511 ( .Y(n4777), .A0(n3562), .A1(n3574) );
  nor02 U1512 ( .Y(n4773), .A0(n4778), .A1(n4779) );
  nor02 U1513 ( .Y(n4780), .A0(n4774), .A1(n4775) );
  inv01 U1514 ( .Y(n4778), .A(n4780) );
  nor02 U1515 ( .Y(n4781), .A0(n4776), .A1(n4777) );
  inv01 U1516 ( .Y(n4779), .A(n4781) );
  buf16 U1517 ( .Y(n6940), .A(count_1_) );
  buf02 U1518 ( .Y(n4782), .A(n7463) );
  nand02 U1519 ( .Y(n7474), .A0(n4783), .A1(n4784) );
  inv01 U1520 ( .Y(n4785), .A(n6970) );
  inv01 U1521 ( .Y(n4786), .A(n6975) );
  inv01 U1522 ( .Y(n4787), .A(larray[171]) );
  inv01 U1523 ( .Y(n4788), .A(larray[75]) );
  nand02 U1524 ( .Y(n4789), .A0(n4785), .A1(n4786) );
  nand02 U1525 ( .Y(n4790), .A0(n4785), .A1(n4787) );
  nand02 U1526 ( .Y(n4791), .A0(n4786), .A1(n4788) );
  nand02 U1527 ( .Y(n4792), .A0(n4787), .A1(n4788) );
  nand02 U1528 ( .Y(n4793), .A0(n4789), .A1(n4790) );
  inv01 U1529 ( .Y(n4783), .A(n4793) );
  nand02 U1530 ( .Y(n4794), .A0(n4791), .A1(n4792) );
  inv01 U1531 ( .Y(n4784), .A(n4794) );
  nand02 U1532 ( .Y(n7516), .A0(n4795), .A1(n4796) );
  inv01 U1533 ( .Y(n4797), .A(n6972) );
  inv01 U1534 ( .Y(n4798), .A(n6975) );
  inv01 U1535 ( .Y(n4799), .A(larray[104]) );
  inv01 U1536 ( .Y(n4800), .A(larray[8]) );
  nand02 U1537 ( .Y(n4801), .A0(n4797), .A1(n4798) );
  nand02 U1538 ( .Y(n4802), .A0(n4797), .A1(n4799) );
  nand02 U1539 ( .Y(n4803), .A0(n4798), .A1(n4800) );
  nand02 U1540 ( .Y(n4804), .A0(n4799), .A1(n4800) );
  nand02 U1541 ( .Y(n4805), .A0(n4801), .A1(n4802) );
  inv01 U1542 ( .Y(n4795), .A(n4805) );
  nand02 U1543 ( .Y(n4806), .A0(n4803), .A1(n4804) );
  inv01 U1544 ( .Y(n4796), .A(n4806) );
  ao22 U1545 ( .Y(n4807), .A0(larray[191]), .A1(n6975), .B0(larray[95]), .B1(
        n6971) );
  inv01 U1546 ( .Y(n4808), .A(n4807) );
  nand02 U1547 ( .Y(n7502), .A0(n4809), .A1(n4810) );
  inv01 U1548 ( .Y(n4811), .A(n6972) );
  inv01 U1549 ( .Y(n4812), .A(n6975) );
  inv01 U1550 ( .Y(n4813), .A(larray[128]) );
  inv01 U1551 ( .Y(n4814), .A(larray[32]) );
  nand02 U1552 ( .Y(n4815), .A0(n4811), .A1(n4812) );
  nand02 U1553 ( .Y(n4816), .A0(n4811), .A1(n4813) );
  nand02 U1554 ( .Y(n4817), .A0(n4812), .A1(n4814) );
  nand02 U1555 ( .Y(n4818), .A0(n4813), .A1(n4814) );
  nand02 U1556 ( .Y(n4819), .A0(n4815), .A1(n4816) );
  inv01 U1557 ( .Y(n4809), .A(n4819) );
  nand02 U1558 ( .Y(n4820), .A0(n4817), .A1(n4818) );
  inv01 U1559 ( .Y(n4810), .A(n4820) );
  nand02 U1560 ( .Y(n7527), .A0(n4821), .A1(n4822) );
  inv01 U1561 ( .Y(n4823), .A(n6972) );
  inv01 U1562 ( .Y(n4824), .A(n6975) );
  inv01 U1563 ( .Y(n4825), .A(larray[115]) );
  inv01 U1564 ( .Y(n4826), .A(larray[19]) );
  nand02 U1565 ( .Y(n4827), .A0(n4823), .A1(n4824) );
  nand02 U1566 ( .Y(n4828), .A0(n4823), .A1(n4825) );
  nand02 U1567 ( .Y(n4829), .A0(n4824), .A1(n4826) );
  nand02 U1568 ( .Y(n4830), .A0(n4825), .A1(n4826) );
  nand02 U1569 ( .Y(n4831), .A0(n4827), .A1(n4828) );
  inv01 U1570 ( .Y(n4821), .A(n4831) );
  nand02 U1571 ( .Y(n4832), .A0(n4829), .A1(n4830) );
  inv01 U1572 ( .Y(n4822), .A(n4832) );
  nand02 U1573 ( .Y(n7493), .A0(n4833), .A1(n4834) );
  inv01 U1574 ( .Y(n4835), .A(n6972) );
  inv01 U1575 ( .Y(n4836), .A(n6975) );
  inv01 U1576 ( .Y(n4837), .A(larray[163]) );
  inv01 U1577 ( .Y(n4838), .A(larray[67]) );
  nand02 U1578 ( .Y(n4839), .A0(n4835), .A1(n4836) );
  nand02 U1579 ( .Y(n4840), .A0(n4835), .A1(n4837) );
  nand02 U1580 ( .Y(n4841), .A0(n4836), .A1(n4838) );
  nand02 U1581 ( .Y(n4842), .A0(n4837), .A1(n4838) );
  nand02 U1582 ( .Y(n4843), .A0(n4839), .A1(n4840) );
  inv01 U1583 ( .Y(n4833), .A(n4843) );
  nand02 U1584 ( .Y(n4844), .A0(n4841), .A1(n4842) );
  inv01 U1585 ( .Y(n4834), .A(n4844) );
  ao22 U1586 ( .Y(n4845), .A0(larray[169]), .A1(n6975), .B0(larray[73]), .B1(
        n6970) );
  inv01 U1587 ( .Y(n4846), .A(n4845) );
  nand02 U1588 ( .Y(n7490), .A0(n4847), .A1(n4848) );
  inv01 U1589 ( .Y(n4849), .A(n6972) );
  inv01 U1590 ( .Y(n4850), .A(n6974) );
  inv01 U1591 ( .Y(n4851), .A(larray[165]) );
  inv01 U1592 ( .Y(n4852), .A(larray[69]) );
  nand02 U1593 ( .Y(n4853), .A0(n4849), .A1(n4850) );
  nand02 U1594 ( .Y(n4854), .A0(n4849), .A1(n4851) );
  nand02 U1595 ( .Y(n4855), .A0(n4850), .A1(n4852) );
  nand02 U1596 ( .Y(n4856), .A0(n4851), .A1(n4852) );
  nand02 U1597 ( .Y(n4857), .A0(n4853), .A1(n4854) );
  inv01 U1598 ( .Y(n4847), .A(n4857) );
  nand02 U1599 ( .Y(n4858), .A0(n4855), .A1(n4856) );
  inv01 U1600 ( .Y(n4848), .A(n4858) );
  nand02 U1601 ( .Y(n7477), .A0(n4859), .A1(n4860) );
  inv01 U1602 ( .Y(n4861), .A(n6972) );
  inv01 U1603 ( .Y(n4862), .A(n6974) );
  inv01 U1604 ( .Y(n4863), .A(larray[187]) );
  inv01 U1605 ( .Y(n4864), .A(larray[91]) );
  nand02 U1606 ( .Y(n4865), .A0(n4861), .A1(n4862) );
  nand02 U1607 ( .Y(n4866), .A0(n4861), .A1(n4863) );
  nand02 U1608 ( .Y(n4867), .A0(n4862), .A1(n4864) );
  nand02 U1609 ( .Y(n4868), .A0(n4863), .A1(n4864) );
  nand02 U1610 ( .Y(n4869), .A0(n4865), .A1(n4866) );
  inv01 U1611 ( .Y(n4859), .A(n4869) );
  nand02 U1612 ( .Y(n4870), .A0(n4867), .A1(n4868) );
  inv01 U1613 ( .Y(n4860), .A(n4870) );
  ao22 U1614 ( .Y(n4871), .A0(larray[160]), .A1(n6974), .B0(larray[64]), .B1(
        n6972) );
  inv01 U1615 ( .Y(n4872), .A(n4871) );
  nand02 U1616 ( .Y(n7503), .A0(n4873), .A1(n4874) );
  inv01 U1617 ( .Y(n4875), .A(n6971) );
  inv01 U1618 ( .Y(n4876), .A(n6975) );
  inv01 U1619 ( .Y(n4877), .A(larray[124]) );
  inv01 U1620 ( .Y(n4878), .A(larray[28]) );
  nand02 U1621 ( .Y(n4879), .A0(n4875), .A1(n4876) );
  nand02 U1622 ( .Y(n4880), .A0(n4875), .A1(n4877) );
  nand02 U1623 ( .Y(n4881), .A0(n4876), .A1(n4878) );
  nand02 U1624 ( .Y(n4882), .A0(n4877), .A1(n4878) );
  nand02 U1625 ( .Y(n4883), .A0(n4879), .A1(n4880) );
  inv01 U1626 ( .Y(n4873), .A(n4883) );
  nand02 U1627 ( .Y(n4884), .A0(n4881), .A1(n4882) );
  inv01 U1628 ( .Y(n4874), .A(n4884) );
  ao22 U1629 ( .Y(n4885), .A0(larray[189]), .A1(n6975), .B0(larray[93]), .B1(
        n6972) );
  inv01 U1630 ( .Y(n4886), .A(n4885) );
  nand02 U1631 ( .Y(n7485), .A0(n4887), .A1(n4888) );
  inv01 U1632 ( .Y(n4889), .A(n6972) );
  inv01 U1633 ( .Y(n4890), .A(n6974) );
  inv01 U1634 ( .Y(n4891), .A(larray[152]) );
  inv01 U1635 ( .Y(n4892), .A(larray[56]) );
  nand02 U1636 ( .Y(n4893), .A0(n4889), .A1(n4890) );
  nand02 U1637 ( .Y(n4894), .A0(n4889), .A1(n4891) );
  nand02 U1638 ( .Y(n4895), .A0(n4890), .A1(n4892) );
  nand02 U1639 ( .Y(n4896), .A0(n4891), .A1(n4892) );
  nand02 U1640 ( .Y(n4897), .A0(n4893), .A1(n4894) );
  inv01 U1641 ( .Y(n4887), .A(n4897) );
  nand02 U1642 ( .Y(n4898), .A0(n4895), .A1(n4896) );
  inv01 U1643 ( .Y(n4888), .A(n4898) );
  nand02 U1644 ( .Y(n7481), .A0(n4899), .A1(n4900) );
  inv01 U1645 ( .Y(n4901), .A(n6972) );
  inv01 U1646 ( .Y(n4902), .A(n6974) );
  inv01 U1647 ( .Y(n4903), .A(larray[181]) );
  inv01 U1648 ( .Y(n4904), .A(larray[85]) );
  nand02 U1649 ( .Y(n4905), .A0(n4901), .A1(n4902) );
  nand02 U1650 ( .Y(n4906), .A0(n4901), .A1(n4903) );
  nand02 U1651 ( .Y(n4907), .A0(n4902), .A1(n4904) );
  nand02 U1652 ( .Y(n4908), .A0(n4903), .A1(n4904) );
  nand02 U1653 ( .Y(n4909), .A0(n4905), .A1(n4906) );
  inv01 U1654 ( .Y(n4899), .A(n4909) );
  nand02 U1655 ( .Y(n4910), .A0(n4907), .A1(n4908) );
  inv01 U1656 ( .Y(n4900), .A(n4910) );
  ao22 U1657 ( .Y(n4911), .A0(larray[162]), .A1(n6974), .B0(larray[66]), .B1(
        n6971) );
  inv01 U1658 ( .Y(n4912), .A(n4911) );
  nand02 U1659 ( .Y(n7479), .A0(n4913), .A1(n4914) );
  inv01 U1660 ( .Y(n4915), .A(n6972) );
  inv01 U1661 ( .Y(n4916), .A(n6975) );
  inv01 U1662 ( .Y(n4917), .A(larray[184]) );
  inv01 U1663 ( .Y(n4918), .A(larray[88]) );
  nand02 U1664 ( .Y(n4919), .A0(n4915), .A1(n4916) );
  nand02 U1665 ( .Y(n4920), .A0(n4915), .A1(n4917) );
  nand02 U1666 ( .Y(n4921), .A0(n4916), .A1(n4918) );
  nand02 U1667 ( .Y(n4922), .A0(n4917), .A1(n4918) );
  nand02 U1668 ( .Y(n4923), .A0(n4919), .A1(n4920) );
  inv01 U1669 ( .Y(n4913), .A(n4923) );
  nand02 U1670 ( .Y(n4924), .A0(n4921), .A1(n4922) );
  inv01 U1671 ( .Y(n4914), .A(n4924) );
  nand02 U1672 ( .Y(n7511), .A0(n4925), .A1(n4926) );
  inv01 U1673 ( .Y(n4927), .A(n6972) );
  inv01 U1674 ( .Y(n4928), .A(n6975) );
  inv01 U1675 ( .Y(n4929), .A(larray[133]) );
  inv01 U1676 ( .Y(n4930), .A(larray[37]) );
  nand02 U1677 ( .Y(n4931), .A0(n4927), .A1(n4928) );
  nand02 U1678 ( .Y(n4932), .A0(n4927), .A1(n4929) );
  nand02 U1679 ( .Y(n4933), .A0(n4928), .A1(n4930) );
  nand02 U1680 ( .Y(n4934), .A0(n4929), .A1(n4930) );
  nand02 U1681 ( .Y(n4935), .A0(n4931), .A1(n4932) );
  inv01 U1682 ( .Y(n4925), .A(n4935) );
  nand02 U1683 ( .Y(n4936), .A0(n4933), .A1(n4934) );
  inv01 U1684 ( .Y(n4926), .A(n4936) );
  nand02 U1685 ( .Y(n7515), .A0(n4937), .A1(n4938) );
  inv01 U1686 ( .Y(n4939), .A(n6971) );
  inv01 U1687 ( .Y(n4940), .A(n6975) );
  inv01 U1688 ( .Y(n4941), .A(larray[120]) );
  inv01 U1689 ( .Y(n4942), .A(larray[24]) );
  nand02 U1690 ( .Y(n4943), .A0(n4939), .A1(n4940) );
  nand02 U1691 ( .Y(n4944), .A0(n4939), .A1(n4941) );
  nand02 U1692 ( .Y(n4945), .A0(n4940), .A1(n4942) );
  nand02 U1693 ( .Y(n4946), .A0(n4941), .A1(n4942) );
  nand02 U1694 ( .Y(n4947), .A0(n4943), .A1(n4944) );
  inv01 U1695 ( .Y(n4937), .A(n4947) );
  nand02 U1696 ( .Y(n4948), .A0(n4945), .A1(n4946) );
  inv01 U1697 ( .Y(n4938), .A(n4948) );
  ao22 U1698 ( .Y(n4949), .A0(larray[139]), .A1(n6975), .B0(larray[43]), .B1(
        n6972) );
  inv01 U1699 ( .Y(n4950), .A(n4949) );
  nand02 U1700 ( .Y(n7492), .A0(n4951), .A1(n4952) );
  inv01 U1701 ( .Y(n4953), .A(n6970) );
  inv01 U1702 ( .Y(n4954), .A(n6974) );
  inv01 U1703 ( .Y(n4955), .A(larray[145]) );
  inv01 U1704 ( .Y(n4956), .A(larray[49]) );
  nand02 U1705 ( .Y(n4957), .A0(n4953), .A1(n4954) );
  nand02 U1706 ( .Y(n4958), .A0(n4953), .A1(n4955) );
  nand02 U1707 ( .Y(n4959), .A0(n4954), .A1(n4956) );
  nand02 U1708 ( .Y(n4960), .A0(n4955), .A1(n4956) );
  nand02 U1709 ( .Y(n4961), .A0(n4957), .A1(n4958) );
  inv01 U1710 ( .Y(n4951), .A(n4961) );
  nand02 U1711 ( .Y(n4962), .A0(n4959), .A1(n4960) );
  inv01 U1712 ( .Y(n4952), .A(n4962) );
  nand02 U1713 ( .Y(n7517), .A0(n4963), .A1(n4964) );
  inv01 U1714 ( .Y(n4965), .A(n6971) );
  inv01 U1715 ( .Y(n4966), .A(n6974) );
  inv01 U1716 ( .Y(n4967), .A(larray[103]) );
  inv01 U1717 ( .Y(n4968), .A(larray[7]) );
  nand02 U1718 ( .Y(n4969), .A0(n4965), .A1(n4966) );
  nand02 U1719 ( .Y(n4970), .A0(n4965), .A1(n4967) );
  nand02 U1720 ( .Y(n4971), .A0(n4966), .A1(n4968) );
  nand02 U1721 ( .Y(n4972), .A0(n4967), .A1(n4968) );
  nand02 U1722 ( .Y(n4973), .A0(n4969), .A1(n4970) );
  inv01 U1723 ( .Y(n4963), .A(n4973) );
  nand02 U1724 ( .Y(n4974), .A0(n4971), .A1(n4972) );
  inv01 U1725 ( .Y(n4964), .A(n4974) );
  nand02 U1726 ( .Y(n7525), .A0(n4975), .A1(n4976) );
  inv01 U1727 ( .Y(n4977), .A(n6972) );
  inv01 U1728 ( .Y(n4978), .A(n6974) );
  inv01 U1729 ( .Y(n4979), .A(larray[117]) );
  inv01 U1730 ( .Y(n4980), .A(larray[21]) );
  nand02 U1731 ( .Y(n4981), .A0(n4977), .A1(n4978) );
  nand02 U1732 ( .Y(n4982), .A0(n4977), .A1(n4979) );
  nand02 U1733 ( .Y(n4983), .A0(n4978), .A1(n4980) );
  nand02 U1734 ( .Y(n4984), .A0(n4979), .A1(n4980) );
  nand02 U1735 ( .Y(n4985), .A0(n4981), .A1(n4982) );
  inv01 U1736 ( .Y(n4975), .A(n4985) );
  nand02 U1737 ( .Y(n4986), .A0(n4983), .A1(n4984) );
  inv01 U1738 ( .Y(n4976), .A(n4986) );
  ao22 U1739 ( .Y(n4987), .A0(larray[123]), .A1(n6974), .B0(larray[27]), .B1(
        n6970) );
  inv01 U1740 ( .Y(n4988), .A(n4987) );
  nand02 U1741 ( .Y(n7491), .A0(n4989), .A1(n4990) );
  inv01 U1742 ( .Y(n4991), .A(n6971) );
  inv01 U1743 ( .Y(n4992), .A(n6975) );
  inv01 U1744 ( .Y(n4993), .A(larray[164]) );
  inv01 U1745 ( .Y(n4994), .A(larray[68]) );
  nand02 U1746 ( .Y(n4995), .A0(n4991), .A1(n4992) );
  nand02 U1747 ( .Y(n4996), .A0(n4991), .A1(n4993) );
  nand02 U1748 ( .Y(n4997), .A0(n4992), .A1(n4994) );
  nand02 U1749 ( .Y(n4998), .A0(n4993), .A1(n4994) );
  nand02 U1750 ( .Y(n4999), .A0(n4995), .A1(n4996) );
  inv01 U1751 ( .Y(n4989), .A(n4999) );
  nand02 U1752 ( .Y(n5000), .A0(n4997), .A1(n4998) );
  inv01 U1753 ( .Y(n4990), .A(n5000) );
  nand02 U1754 ( .Y(n7489), .A0(n5001), .A1(n5002) );
  inv01 U1755 ( .Y(n5003), .A(n6970) );
  inv01 U1756 ( .Y(n5004), .A(n6975) );
  inv01 U1757 ( .Y(n5005), .A(larray[166]) );
  inv01 U1758 ( .Y(n5006), .A(larray[70]) );
  nand02 U1759 ( .Y(n5007), .A0(n5003), .A1(n5004) );
  nand02 U1760 ( .Y(n5008), .A0(n5003), .A1(n5005) );
  nand02 U1761 ( .Y(n5009), .A0(n5004), .A1(n5006) );
  nand02 U1762 ( .Y(n5010), .A0(n5005), .A1(n5006) );
  nand02 U1763 ( .Y(n5011), .A0(n5007), .A1(n5008) );
  inv01 U1764 ( .Y(n5001), .A(n5011) );
  nand02 U1765 ( .Y(n5012), .A0(n5009), .A1(n5010) );
  inv01 U1766 ( .Y(n5002), .A(n5012) );
  nand02 U1767 ( .Y(n7494), .A0(n5013), .A1(n5014) );
  inv01 U1768 ( .Y(n5015), .A(n6971) );
  inv01 U1769 ( .Y(n5016), .A(n6975) );
  inv01 U1770 ( .Y(n5017), .A(larray[159]) );
  inv01 U1771 ( .Y(n5018), .A(larray[63]) );
  nand02 U1772 ( .Y(n5019), .A0(n5015), .A1(n5016) );
  nand02 U1773 ( .Y(n5020), .A0(n5015), .A1(n5017) );
  nand02 U1774 ( .Y(n5021), .A0(n5016), .A1(n5018) );
  nand02 U1775 ( .Y(n5022), .A0(n5017), .A1(n5018) );
  nand02 U1776 ( .Y(n5023), .A0(n5019), .A1(n5020) );
  inv01 U1777 ( .Y(n5013), .A(n5023) );
  nand02 U1778 ( .Y(n5024), .A0(n5021), .A1(n5022) );
  inv01 U1779 ( .Y(n5014), .A(n5024) );
  ao22 U1780 ( .Y(n5025), .A0(larray[182]), .A1(n6975), .B0(larray[86]), .B1(
        n6970) );
  inv01 U1781 ( .Y(n5026), .A(n5025) );
  nand02 U1782 ( .Y(n7521), .A0(n5027), .A1(n5028) );
  inv01 U1783 ( .Y(n5029), .A(n6970) );
  inv01 U1784 ( .Y(n5030), .A(n6974) );
  inv01 U1785 ( .Y(n5031), .A(larray[99]) );
  inv01 U1786 ( .Y(n5032), .A(larray[3]) );
  nand02 U1787 ( .Y(n5033), .A0(n5029), .A1(n5030) );
  nand02 U1788 ( .Y(n5034), .A0(n5029), .A1(n5031) );
  nand02 U1789 ( .Y(n5035), .A0(n5030), .A1(n5032) );
  nand02 U1790 ( .Y(n5036), .A0(n5031), .A1(n5032) );
  nand02 U1791 ( .Y(n5037), .A0(n5033), .A1(n5034) );
  inv01 U1792 ( .Y(n5027), .A(n5037) );
  nand02 U1793 ( .Y(n5038), .A0(n5035), .A1(n5036) );
  inv01 U1794 ( .Y(n5028), .A(n5038) );
  nand02 U1795 ( .Y(n7495), .A0(n5039), .A1(n5040) );
  inv01 U1796 ( .Y(n5041), .A(n6970) );
  inv01 U1797 ( .Y(n5042), .A(n6974) );
  inv01 U1798 ( .Y(n5043), .A(larray[158]) );
  inv01 U1799 ( .Y(n5044), .A(larray[62]) );
  nand02 U1800 ( .Y(n5045), .A0(n5041), .A1(n5042) );
  nand02 U1801 ( .Y(n5046), .A0(n5041), .A1(n5043) );
  nand02 U1802 ( .Y(n5047), .A0(n5042), .A1(n5044) );
  nand02 U1803 ( .Y(n5048), .A0(n5043), .A1(n5044) );
  nand02 U1804 ( .Y(n5049), .A0(n5045), .A1(n5046) );
  inv01 U1805 ( .Y(n5039), .A(n5049) );
  nand02 U1806 ( .Y(n5050), .A0(n5047), .A1(n5048) );
  inv01 U1807 ( .Y(n5040), .A(n5050) );
  nand02 U1808 ( .Y(n7483), .A0(n5051), .A1(n5052) );
  inv01 U1809 ( .Y(n5053), .A(n6971) );
  inv01 U1810 ( .Y(n5054), .A(n6974) );
  inv01 U1811 ( .Y(n5055), .A(larray[168]) );
  inv01 U1812 ( .Y(n5056), .A(larray[72]) );
  nand02 U1813 ( .Y(n5057), .A0(n5053), .A1(n5054) );
  nand02 U1814 ( .Y(n5058), .A0(n5053), .A1(n5055) );
  nand02 U1815 ( .Y(n5059), .A0(n5054), .A1(n5056) );
  nand02 U1816 ( .Y(n5060), .A0(n5055), .A1(n5056) );
  nand02 U1817 ( .Y(n5061), .A0(n5057), .A1(n5058) );
  inv01 U1818 ( .Y(n5051), .A(n5061) );
  nand02 U1819 ( .Y(n5062), .A0(n5059), .A1(n5060) );
  inv01 U1820 ( .Y(n5052), .A(n5062) );
  ao22 U1821 ( .Y(n5063), .A0(larray[121]), .A1(n6974), .B0(larray[25]), .B1(
        n6970) );
  inv01 U1822 ( .Y(n5064), .A(n5063) );
  nand02 U1823 ( .Y(n7520), .A0(n5065), .A1(n5066) );
  inv01 U1824 ( .Y(n5067), .A(n6971) );
  inv01 U1825 ( .Y(n5068), .A(n6975) );
  inv01 U1826 ( .Y(n5069), .A(larray[100]) );
  inv01 U1827 ( .Y(n5070), .A(larray[4]) );
  nand02 U1828 ( .Y(n5071), .A0(n5067), .A1(n5068) );
  nand02 U1829 ( .Y(n5072), .A0(n5067), .A1(n5069) );
  nand02 U1830 ( .Y(n5073), .A0(n5068), .A1(n5070) );
  nand02 U1831 ( .Y(n5074), .A0(n5069), .A1(n5070) );
  nand02 U1832 ( .Y(n5075), .A0(n5071), .A1(n5072) );
  inv01 U1833 ( .Y(n5065), .A(n5075) );
  nand02 U1834 ( .Y(n5076), .A0(n5073), .A1(n5074) );
  inv01 U1835 ( .Y(n5066), .A(n5076) );
  nand02 U1836 ( .Y(n7533), .A0(n5077), .A1(n5078) );
  inv01 U1837 ( .Y(n5079), .A(n6971) );
  inv01 U1838 ( .Y(n5080), .A(n6975) );
  inv01 U1839 ( .Y(n5081), .A(larray[96]) );
  inv01 U1840 ( .Y(n5082), .A(larray[0]) );
  nand02 U1841 ( .Y(n5083), .A0(n5079), .A1(n5080) );
  nand02 U1842 ( .Y(n5084), .A0(n5079), .A1(n5081) );
  nand02 U1843 ( .Y(n5085), .A0(n5080), .A1(n5082) );
  nand02 U1844 ( .Y(n5086), .A0(n5081), .A1(n5082) );
  nand02 U1845 ( .Y(n5087), .A0(n5083), .A1(n5084) );
  inv01 U1846 ( .Y(n5077), .A(n5087) );
  nand02 U1847 ( .Y(n5088), .A0(n5085), .A1(n5086) );
  inv01 U1848 ( .Y(n5078), .A(n5088) );
  ao22 U1849 ( .Y(n5089), .A0(larray[135]), .A1(n6975), .B0(larray[39]), .B1(
        n6971) );
  inv01 U1850 ( .Y(n5090), .A(n5089) );
  nand02 U1851 ( .Y(n7531), .A0(n5091), .A1(n5092) );
  inv01 U1852 ( .Y(n5093), .A(n6971) );
  inv01 U1853 ( .Y(n5094), .A(n6974) );
  inv01 U1854 ( .Y(n5095), .A(larray[108]) );
  inv01 U1855 ( .Y(n5096), .A(larray[12]) );
  nand02 U1856 ( .Y(n5097), .A0(n5093), .A1(n5094) );
  nand02 U1857 ( .Y(n5098), .A0(n5093), .A1(n5095) );
  nand02 U1858 ( .Y(n5099), .A0(n5094), .A1(n5096) );
  nand02 U1859 ( .Y(n5100), .A0(n5095), .A1(n5096) );
  nand02 U1860 ( .Y(n5101), .A0(n5097), .A1(n5098) );
  inv01 U1861 ( .Y(n5091), .A(n5101) );
  nand02 U1862 ( .Y(n5102), .A0(n5099), .A1(n5100) );
  inv01 U1863 ( .Y(n5092), .A(n5102) );
  nand02 U1864 ( .Y(n7497), .A0(n5103), .A1(n5104) );
  inv01 U1865 ( .Y(n5105), .A(n6971) );
  inv01 U1866 ( .Y(n5106), .A(n6974) );
  inv01 U1867 ( .Y(n5107), .A(larray[156]) );
  inv01 U1868 ( .Y(n5108), .A(larray[60]) );
  nand02 U1869 ( .Y(n5109), .A0(n5105), .A1(n5106) );
  nand02 U1870 ( .Y(n5110), .A0(n5105), .A1(n5107) );
  nand02 U1871 ( .Y(n5111), .A0(n5106), .A1(n5108) );
  nand02 U1872 ( .Y(n5112), .A0(n5107), .A1(n5108) );
  nand02 U1873 ( .Y(n5113), .A0(n5109), .A1(n5110) );
  inv01 U1874 ( .Y(n5103), .A(n5113) );
  nand02 U1875 ( .Y(n5114), .A0(n5111), .A1(n5112) );
  inv01 U1876 ( .Y(n5104), .A(n5114) );
  nand02 U1877 ( .Y(n7480), .A0(n5115), .A1(n5116) );
  inv01 U1878 ( .Y(n5117), .A(n6971) );
  inv01 U1879 ( .Y(n5118), .A(n6974) );
  inv01 U1880 ( .Y(n5119), .A(larray[183]) );
  inv01 U1881 ( .Y(n5120), .A(larray[87]) );
  nand02 U1882 ( .Y(n5121), .A0(n5117), .A1(n5118) );
  nand02 U1883 ( .Y(n5122), .A0(n5117), .A1(n5119) );
  nand02 U1884 ( .Y(n5123), .A0(n5118), .A1(n5120) );
  nand02 U1885 ( .Y(n5124), .A0(n5119), .A1(n5120) );
  nand02 U1886 ( .Y(n5125), .A0(n5121), .A1(n5122) );
  inv01 U1887 ( .Y(n5115), .A(n5125) );
  nand02 U1888 ( .Y(n5126), .A0(n5123), .A1(n5124) );
  inv01 U1889 ( .Y(n5116), .A(n5126) );
  ao22 U1890 ( .Y(n5127), .A0(larray[146]), .A1(n6974), .B0(larray[50]), .B1(
        n6972) );
  inv01 U1891 ( .Y(n5128), .A(n5127) );
  nand02 U1892 ( .Y(n7526), .A0(n5129), .A1(n5130) );
  inv01 U1893 ( .Y(n5131), .A(n6971) );
  inv01 U1894 ( .Y(n5132), .A(n6975) );
  inv01 U1895 ( .Y(n5133), .A(larray[116]) );
  inv01 U1896 ( .Y(n5134), .A(larray[20]) );
  nand02 U1897 ( .Y(n5135), .A0(n5131), .A1(n5132) );
  nand02 U1898 ( .Y(n5136), .A0(n5131), .A1(n5133) );
  nand02 U1899 ( .Y(n5137), .A0(n5132), .A1(n5134) );
  nand02 U1900 ( .Y(n5138), .A0(n5133), .A1(n5134) );
  nand02 U1901 ( .Y(n5139), .A0(n5135), .A1(n5136) );
  inv01 U1902 ( .Y(n5129), .A(n5139) );
  nand02 U1903 ( .Y(n5140), .A0(n5137), .A1(n5138) );
  inv01 U1904 ( .Y(n5130), .A(n5140) );
  nand02 U1905 ( .Y(n7496), .A0(n5141), .A1(n5142) );
  inv01 U1906 ( .Y(n5143), .A(n6972) );
  inv01 U1907 ( .Y(n5144), .A(n6975) );
  inv01 U1908 ( .Y(n5145), .A(larray[157]) );
  inv01 U1909 ( .Y(n5146), .A(larray[61]) );
  nand02 U1910 ( .Y(n5147), .A0(n5143), .A1(n5144) );
  nand02 U1911 ( .Y(n5148), .A0(n5143), .A1(n5145) );
  nand02 U1912 ( .Y(n5149), .A0(n5144), .A1(n5146) );
  nand02 U1913 ( .Y(n5150), .A0(n5145), .A1(n5146) );
  nand02 U1914 ( .Y(n5151), .A0(n5147), .A1(n5148) );
  inv01 U1915 ( .Y(n5141), .A(n5151) );
  nand02 U1916 ( .Y(n5152), .A0(n5149), .A1(n5150) );
  inv01 U1917 ( .Y(n5142), .A(n5152) );
  nand02 U1918 ( .Y(n7522), .A0(n5153), .A1(n5154) );
  inv01 U1919 ( .Y(n5155), .A(n6972) );
  inv01 U1920 ( .Y(n5156), .A(n6975) );
  inv01 U1921 ( .Y(n5157), .A(larray[98]) );
  inv01 U1922 ( .Y(n5158), .A(larray[2]) );
  nand02 U1923 ( .Y(n5159), .A0(n5155), .A1(n5156) );
  nand02 U1924 ( .Y(n5160), .A0(n5155), .A1(n5157) );
  nand02 U1925 ( .Y(n5161), .A0(n5156), .A1(n5158) );
  nand02 U1926 ( .Y(n5162), .A0(n5157), .A1(n5158) );
  nand02 U1927 ( .Y(n5163), .A0(n5159), .A1(n5160) );
  inv01 U1928 ( .Y(n5153), .A(n5163) );
  nand02 U1929 ( .Y(n5164), .A0(n5161), .A1(n5162) );
  inv01 U1930 ( .Y(n5154), .A(n5164) );
  ao22 U1931 ( .Y(n5165), .A0(larray[151]), .A1(n6975), .B0(larray[55]), .B1(
        n6971) );
  inv01 U1932 ( .Y(n5166), .A(n5165) );
  nand02 U1933 ( .Y(n7514), .A0(n5167), .A1(n5168) );
  inv01 U1934 ( .Y(n5169), .A(n6972) );
  inv01 U1935 ( .Y(n5170), .A(n6974) );
  inv01 U1936 ( .Y(n5171), .A(larray[130]) );
  inv01 U1937 ( .Y(n5172), .A(larray[34]) );
  nand02 U1938 ( .Y(n5173), .A0(n5169), .A1(n5170) );
  nand02 U1939 ( .Y(n5174), .A0(n5169), .A1(n5171) );
  nand02 U1940 ( .Y(n5175), .A0(n5170), .A1(n5172) );
  nand02 U1941 ( .Y(n5176), .A0(n5171), .A1(n5172) );
  nand02 U1942 ( .Y(n5177), .A0(n5173), .A1(n5174) );
  inv01 U1943 ( .Y(n5167), .A(n5177) );
  nand02 U1944 ( .Y(n5178), .A0(n5175), .A1(n5176) );
  inv01 U1945 ( .Y(n5168), .A(n5178) );
  ao22 U1946 ( .Y(n5179), .A0(larray[127]), .A1(n6974), .B0(larray[31]), .B1(
        n6971) );
  inv01 U1947 ( .Y(n5180), .A(n5179) );
  nand02 U1948 ( .Y(n7523), .A0(n5181), .A1(n5182) );
  inv01 U1949 ( .Y(n5183), .A(n6971) );
  inv01 U1950 ( .Y(n5184), .A(n6974) );
  inv01 U1951 ( .Y(n5185), .A(larray[119]) );
  inv01 U1952 ( .Y(n5186), .A(larray[23]) );
  nand02 U1953 ( .Y(n5187), .A0(n5183), .A1(n5184) );
  nand02 U1954 ( .Y(n5188), .A0(n5183), .A1(n5185) );
  nand02 U1955 ( .Y(n5189), .A0(n5184), .A1(n5186) );
  nand02 U1956 ( .Y(n5190), .A0(n5185), .A1(n5186) );
  nand02 U1957 ( .Y(n5191), .A0(n5187), .A1(n5188) );
  inv01 U1958 ( .Y(n5181), .A(n5191) );
  nand02 U1959 ( .Y(n5192), .A0(n5189), .A1(n5190) );
  inv01 U1960 ( .Y(n5182), .A(n5192) );
  nand02 U1961 ( .Y(n7509), .A0(n5193), .A1(n5194) );
  inv01 U1962 ( .Y(n5195), .A(n6972) );
  inv01 U1963 ( .Y(n5196), .A(n6974) );
  inv01 U1964 ( .Y(n5197), .A(larray[136]) );
  inv01 U1965 ( .Y(n5198), .A(larray[40]) );
  nand02 U1966 ( .Y(n5199), .A0(n5195), .A1(n5196) );
  nand02 U1967 ( .Y(n5200), .A0(n5195), .A1(n5197) );
  nand02 U1968 ( .Y(n5201), .A0(n5196), .A1(n5198) );
  nand02 U1969 ( .Y(n5202), .A0(n5197), .A1(n5198) );
  nand02 U1970 ( .Y(n5203), .A0(n5199), .A1(n5200) );
  inv01 U1971 ( .Y(n5193), .A(n5203) );
  nand02 U1972 ( .Y(n5204), .A0(n5201), .A1(n5202) );
  inv01 U1973 ( .Y(n5194), .A(n5204) );
  ao22 U1974 ( .Y(n5205), .A0(larray[112]), .A1(n6974), .B0(larray[16]), .B1(
        n6972) );
  inv01 U1975 ( .Y(n5206), .A(n5205) );
  nand02 U1976 ( .Y(n7505), .A0(n5207), .A1(n5208) );
  inv01 U1977 ( .Y(n5209), .A(n6970) );
  inv01 U1978 ( .Y(n5210), .A(n6975) );
  inv01 U1979 ( .Y(n5211), .A(larray[142]) );
  inv01 U1980 ( .Y(n5212), .A(larray[46]) );
  nand02 U1981 ( .Y(n5213), .A0(n5209), .A1(n5210) );
  nand02 U1982 ( .Y(n5214), .A0(n5209), .A1(n5211) );
  nand02 U1983 ( .Y(n5215), .A0(n5210), .A1(n5212) );
  nand02 U1984 ( .Y(n5216), .A0(n5211), .A1(n5212) );
  nand02 U1985 ( .Y(n5217), .A0(n5213), .A1(n5214) );
  inv01 U1986 ( .Y(n5207), .A(n5217) );
  nand02 U1987 ( .Y(n5218), .A0(n5215), .A1(n5216) );
  inv01 U1988 ( .Y(n5208), .A(n5218) );
  nand02 U1989 ( .Y(n7532), .A0(n5219), .A1(n5220) );
  inv01 U1990 ( .Y(n5221), .A(n6970) );
  inv01 U1991 ( .Y(n5222), .A(n6975) );
  inv01 U1992 ( .Y(n5223), .A(larray[107]) );
  inv01 U1993 ( .Y(n5224), .A(larray[11]) );
  nand02 U1994 ( .Y(n5225), .A0(n5221), .A1(n5222) );
  nand02 U1995 ( .Y(n5226), .A0(n5221), .A1(n5223) );
  nand02 U1996 ( .Y(n5227), .A0(n5222), .A1(n5224) );
  nand02 U1997 ( .Y(n5228), .A0(n5223), .A1(n5224) );
  nand02 U1998 ( .Y(n5229), .A0(n5225), .A1(n5226) );
  inv01 U1999 ( .Y(n5219), .A(n5229) );
  nand02 U2000 ( .Y(n5230), .A0(n5227), .A1(n5228) );
  inv01 U2001 ( .Y(n5220), .A(n5230) );
  nand02 U2002 ( .Y(n7518), .A0(n5231), .A1(n5232) );
  inv01 U2003 ( .Y(n5233), .A(n6970) );
  inv01 U2004 ( .Y(n5234), .A(n6975) );
  inv01 U2005 ( .Y(n5235), .A(larray[102]) );
  inv01 U2006 ( .Y(n5236), .A(larray[6]) );
  nand02 U2007 ( .Y(n5237), .A0(n5233), .A1(n5234) );
  nand02 U2008 ( .Y(n5238), .A0(n5233), .A1(n5235) );
  nand02 U2009 ( .Y(n5239), .A0(n5234), .A1(n5236) );
  nand02 U2010 ( .Y(n5240), .A0(n5235), .A1(n5236) );
  nand02 U2011 ( .Y(n5241), .A0(n5237), .A1(n5238) );
  inv01 U2012 ( .Y(n5231), .A(n5241) );
  nand02 U2013 ( .Y(n5242), .A0(n5239), .A1(n5240) );
  inv01 U2014 ( .Y(n5232), .A(n5242) );
  ao22 U2015 ( .Y(n5243), .A0(larray[113]), .A1(n6975), .B0(larray[17]), .B1(
        n6970) );
  inv01 U2016 ( .Y(n5244), .A(n5243) );
  nand02 U2017 ( .Y(n7519), .A0(n5245), .A1(n5246) );
  inv01 U2018 ( .Y(n5247), .A(n6972) );
  inv01 U2019 ( .Y(n5248), .A(n6974) );
  inv01 U2020 ( .Y(n5249), .A(larray[101]) );
  inv01 U2021 ( .Y(n5250), .A(larray[5]) );
  nand02 U2022 ( .Y(n5251), .A0(n5247), .A1(n5248) );
  nand02 U2023 ( .Y(n5252), .A0(n5247), .A1(n5249) );
  nand02 U2024 ( .Y(n5253), .A0(n5248), .A1(n5250) );
  nand02 U2025 ( .Y(n5254), .A0(n5249), .A1(n5250) );
  nand02 U2026 ( .Y(n5255), .A0(n5251), .A1(n5252) );
  inv01 U2027 ( .Y(n5245), .A(n5255) );
  nand02 U2028 ( .Y(n5256), .A0(n5253), .A1(n5254) );
  inv01 U2029 ( .Y(n5246), .A(n5256) );
  ao22 U2030 ( .Y(n5257), .A0(larray[185]), .A1(n6974), .B0(larray[89]), .B1(
        n6970) );
  inv01 U2031 ( .Y(n5258), .A(n5257) );
  nand02 U2032 ( .Y(n7528), .A0(n5259), .A1(n5260) );
  inv01 U2033 ( .Y(n5261), .A(n6971) );
  inv01 U2034 ( .Y(n5262), .A(n6975) );
  inv01 U2035 ( .Y(n5263), .A(larray[111]) );
  inv01 U2036 ( .Y(n5264), .A(larray[15]) );
  nand02 U2037 ( .Y(n5265), .A0(n5261), .A1(n5262) );
  nand02 U2038 ( .Y(n5266), .A0(n5261), .A1(n5263) );
  nand02 U2039 ( .Y(n5267), .A0(n5262), .A1(n5264) );
  nand02 U2040 ( .Y(n5268), .A0(n5263), .A1(n5264) );
  nand02 U2041 ( .Y(n5269), .A0(n5265), .A1(n5266) );
  inv01 U2042 ( .Y(n5259), .A(n5269) );
  nand02 U2043 ( .Y(n5270), .A0(n5267), .A1(n5268) );
  inv01 U2044 ( .Y(n5260), .A(n5270) );
  nand02 U2045 ( .Y(n7524), .A0(n5271), .A1(n5272) );
  inv01 U2046 ( .Y(n5273), .A(n6970) );
  inv01 U2047 ( .Y(n5274), .A(n6975) );
  inv01 U2048 ( .Y(n5275), .A(larray[118]) );
  inv01 U2049 ( .Y(n5276), .A(larray[22]) );
  nand02 U2050 ( .Y(n5277), .A0(n5273), .A1(n5274) );
  nand02 U2051 ( .Y(n5278), .A0(n5273), .A1(n5275) );
  nand02 U2052 ( .Y(n5279), .A0(n5274), .A1(n5276) );
  nand02 U2053 ( .Y(n5280), .A0(n5275), .A1(n5276) );
  nand02 U2054 ( .Y(n5281), .A0(n5277), .A1(n5278) );
  inv01 U2055 ( .Y(n5271), .A(n5281) );
  nand02 U2056 ( .Y(n5282), .A0(n5279), .A1(n5280) );
  inv01 U2057 ( .Y(n5272), .A(n5282) );
  ao22 U2058 ( .Y(n5283), .A0(larray[175]), .A1(n6975), .B0(larray[79]), .B1(
        n6971) );
  inv01 U2059 ( .Y(n5284), .A(n5283) );
  nand02 U2060 ( .Y(n7499), .A0(n5285), .A1(n5286) );
  inv01 U2061 ( .Y(n5287), .A(n6972) );
  inv01 U2062 ( .Y(n5288), .A(n6974) );
  inv01 U2063 ( .Y(n5289), .A(larray[154]) );
  inv01 U2064 ( .Y(n5290), .A(larray[58]) );
  nand02 U2065 ( .Y(n5291), .A0(n5287), .A1(n5288) );
  nand02 U2066 ( .Y(n5292), .A0(n5287), .A1(n5289) );
  nand02 U2067 ( .Y(n5293), .A0(n5288), .A1(n5290) );
  nand02 U2068 ( .Y(n5294), .A0(n5289), .A1(n5290) );
  nand02 U2069 ( .Y(n5295), .A0(n5291), .A1(n5292) );
  inv01 U2070 ( .Y(n5285), .A(n5295) );
  nand02 U2071 ( .Y(n5296), .A0(n5293), .A1(n5294) );
  inv01 U2072 ( .Y(n5286), .A(n5296) );
  nand02 U2073 ( .Y(n7472), .A0(n5297), .A1(n5298) );
  inv01 U2074 ( .Y(n5299), .A(n6970) );
  inv01 U2075 ( .Y(n5300), .A(n6974) );
  inv01 U2076 ( .Y(n5301), .A(larray[174]) );
  inv01 U2077 ( .Y(n5302), .A(larray[78]) );
  nand02 U2078 ( .Y(n5303), .A0(n5299), .A1(n5300) );
  nand02 U2079 ( .Y(n5304), .A0(n5299), .A1(n5301) );
  nand02 U2080 ( .Y(n5305), .A0(n5300), .A1(n5302) );
  nand02 U2081 ( .Y(n5306), .A0(n5301), .A1(n5302) );
  nand02 U2082 ( .Y(n5307), .A0(n5303), .A1(n5304) );
  inv01 U2083 ( .Y(n5297), .A(n5307) );
  nand02 U2084 ( .Y(n5308), .A0(n5305), .A1(n5306) );
  inv01 U2085 ( .Y(n5298), .A(n5308) );
  nand02 U2086 ( .Y(n7529), .A0(n5309), .A1(n5310) );
  inv01 U2087 ( .Y(n5311), .A(n6970) );
  inv01 U2088 ( .Y(n5312), .A(n6974) );
  inv01 U2089 ( .Y(n5313), .A(larray[110]) );
  inv01 U2090 ( .Y(n5314), .A(larray[14]) );
  nand02 U2091 ( .Y(n5315), .A0(n5311), .A1(n5312) );
  nand02 U2092 ( .Y(n5316), .A0(n5311), .A1(n5313) );
  nand02 U2093 ( .Y(n5317), .A0(n5312), .A1(n5314) );
  nand02 U2094 ( .Y(n5318), .A0(n5313), .A1(n5314) );
  nand02 U2095 ( .Y(n5319), .A0(n5315), .A1(n5316) );
  inv01 U2096 ( .Y(n5309), .A(n5319) );
  nand02 U2097 ( .Y(n5320), .A0(n5317), .A1(n5318) );
  inv01 U2098 ( .Y(n5310), .A(n5320) );
  ao22 U2099 ( .Y(n5321), .A0(larray[125]), .A1(n6974), .B0(larray[29]), .B1(
        n6972) );
  inv01 U2100 ( .Y(n5322), .A(n5321) );
  nand02 U2101 ( .Y(n7500), .A0(n5323), .A1(n5324) );
  inv01 U2102 ( .Y(n5325), .A(n6971) );
  inv01 U2103 ( .Y(n5326), .A(n6975) );
  inv01 U2104 ( .Y(n5327), .A(larray[144]) );
  inv01 U2105 ( .Y(n5328), .A(larray[48]) );
  nand02 U2106 ( .Y(n5329), .A0(n5325), .A1(n5326) );
  nand02 U2107 ( .Y(n5330), .A0(n5325), .A1(n5327) );
  nand02 U2108 ( .Y(n5331), .A0(n5326), .A1(n5328) );
  nand02 U2109 ( .Y(n5332), .A0(n5327), .A1(n5328) );
  nand02 U2110 ( .Y(n5333), .A0(n5329), .A1(n5330) );
  inv01 U2111 ( .Y(n5323), .A(n5333) );
  nand02 U2112 ( .Y(n5334), .A0(n5331), .A1(n5332) );
  inv01 U2113 ( .Y(n5324), .A(n5334) );
  nand02 U2114 ( .Y(n7513), .A0(n5335), .A1(n5336) );
  inv01 U2115 ( .Y(n5337), .A(n6970) );
  inv01 U2116 ( .Y(n5338), .A(n6975) );
  inv01 U2117 ( .Y(n5339), .A(larray[131]) );
  inv01 U2118 ( .Y(n5340), .A(larray[35]) );
  nand02 U2119 ( .Y(n5341), .A0(n5337), .A1(n5338) );
  nand02 U2120 ( .Y(n5342), .A0(n5337), .A1(n5339) );
  nand02 U2121 ( .Y(n5343), .A0(n5338), .A1(n5340) );
  nand02 U2122 ( .Y(n5344), .A0(n5339), .A1(n5340) );
  nand02 U2123 ( .Y(n5345), .A0(n5341), .A1(n5342) );
  inv01 U2124 ( .Y(n5335), .A(n5345) );
  nand02 U2125 ( .Y(n5346), .A0(n5343), .A1(n5344) );
  inv01 U2126 ( .Y(n5336), .A(n5346) );
  ao22 U2127 ( .Y(n5347), .A0(larray[161]), .A1(n6975), .B0(larray[65]), .B1(
        n6970) );
  inv01 U2128 ( .Y(n5348), .A(n5347) );
  nand02 U2129 ( .Y(n7473), .A0(n5349), .A1(n5350) );
  inv01 U2130 ( .Y(n5351), .A(n6972) );
  inv01 U2131 ( .Y(n5352), .A(n6975) );
  inv01 U2132 ( .Y(n5353), .A(larray[173]) );
  inv01 U2133 ( .Y(n5354), .A(larray[77]) );
  nand02 U2134 ( .Y(n5355), .A0(n5351), .A1(n5352) );
  nand02 U2135 ( .Y(n5356), .A0(n5351), .A1(n5353) );
  nand02 U2136 ( .Y(n5357), .A0(n5352), .A1(n5354) );
  nand02 U2137 ( .Y(n5358), .A0(n5353), .A1(n5354) );
  nand02 U2138 ( .Y(n5359), .A0(n5355), .A1(n5356) );
  inv01 U2139 ( .Y(n5349), .A(n5359) );
  nand02 U2140 ( .Y(n5360), .A0(n5357), .A1(n5358) );
  inv01 U2141 ( .Y(n5350), .A(n5360) );
  ao22 U2142 ( .Y(n5361), .A0(larray[178]), .A1(n6975), .B0(larray[82]), .B1(
        n6972) );
  inv01 U2143 ( .Y(n5362), .A(n5361) );
  nand02 U2144 ( .Y(n7482), .A0(n5363), .A1(n5364) );
  inv01 U2145 ( .Y(n5365), .A(n6970) );
  inv01 U2146 ( .Y(n5366), .A(n6974) );
  inv01 U2147 ( .Y(n5367), .A(larray[179]) );
  inv01 U2148 ( .Y(n5368), .A(larray[83]) );
  nand02 U2149 ( .Y(n5369), .A0(n5365), .A1(n5366) );
  nand02 U2150 ( .Y(n5370), .A0(n5365), .A1(n5367) );
  nand02 U2151 ( .Y(n5371), .A0(n5366), .A1(n5368) );
  nand02 U2152 ( .Y(n5372), .A0(n5367), .A1(n5368) );
  nand02 U2153 ( .Y(n5373), .A0(n5369), .A1(n5370) );
  inv01 U2154 ( .Y(n5363), .A(n5373) );
  nand02 U2155 ( .Y(n5374), .A0(n5371), .A1(n5372) );
  inv01 U2156 ( .Y(n5364), .A(n5374) );
  nand02 U2157 ( .Y(n7504), .A0(n5375), .A1(n5376) );
  inv01 U2158 ( .Y(n5377), .A(n6971) );
  inv01 U2159 ( .Y(n5378), .A(n6974) );
  inv01 U2160 ( .Y(n5379), .A(larray[143]) );
  inv01 U2161 ( .Y(n5380), .A(larray[47]) );
  nand02 U2162 ( .Y(n5381), .A0(n5377), .A1(n5378) );
  nand02 U2163 ( .Y(n5382), .A0(n5377), .A1(n5379) );
  nand02 U2164 ( .Y(n5383), .A0(n5378), .A1(n5380) );
  nand02 U2165 ( .Y(n5384), .A0(n5379), .A1(n5380) );
  nand02 U2166 ( .Y(n5385), .A0(n5381), .A1(n5382) );
  inv01 U2167 ( .Y(n5375), .A(n5385) );
  nand02 U2168 ( .Y(n5386), .A0(n5383), .A1(n5384) );
  inv01 U2169 ( .Y(n5376), .A(n5386) );
  ao22 U2170 ( .Y(n5387), .A0(larray[97]), .A1(n6974), .B0(larray[1]), .B1(
        n6970) );
  inv01 U2171 ( .Y(n5388), .A(n5387) );
  nand02 U2172 ( .Y(n7470), .A0(n5389), .A1(n5390) );
  inv01 U2173 ( .Y(n5391), .A(n6970) );
  inv01 U2174 ( .Y(n5392), .A(n6975) );
  inv01 U2175 ( .Y(n5393), .A(larray[177]) );
  inv01 U2176 ( .Y(n5394), .A(larray[81]) );
  nand02 U2177 ( .Y(n5395), .A0(n5391), .A1(n5392) );
  nand02 U2178 ( .Y(n5396), .A0(n5391), .A1(n5393) );
  nand02 U2179 ( .Y(n5397), .A0(n5392), .A1(n5394) );
  nand02 U2180 ( .Y(n5398), .A0(n5393), .A1(n5394) );
  nand02 U2181 ( .Y(n5399), .A0(n5395), .A1(n5396) );
  inv01 U2182 ( .Y(n5389), .A(n5399) );
  nand02 U2183 ( .Y(n5400), .A0(n5397), .A1(n5398) );
  inv01 U2184 ( .Y(n5390), .A(n5400) );
  ao22 U2185 ( .Y(n5401), .A0(larray[137]), .A1(n6975), .B0(larray[41]), .B1(
        n6970) );
  inv01 U2186 ( .Y(n5402), .A(n5401) );
  nand02 U2187 ( .Y(n7471), .A0(n5403), .A1(n5404) );
  inv01 U2188 ( .Y(n5405), .A(n6972) );
  inv01 U2189 ( .Y(n5406), .A(n6974) );
  inv01 U2190 ( .Y(n5407), .A(larray[176]) );
  inv01 U2191 ( .Y(n5408), .A(larray[80]) );
  nand02 U2192 ( .Y(n5409), .A0(n5405), .A1(n5406) );
  nand02 U2193 ( .Y(n5410), .A0(n5405), .A1(n5407) );
  nand02 U2194 ( .Y(n5411), .A0(n5406), .A1(n5408) );
  nand02 U2195 ( .Y(n5412), .A0(n5407), .A1(n5408) );
  nand02 U2196 ( .Y(n5413), .A0(n5409), .A1(n5410) );
  inv01 U2197 ( .Y(n5403), .A(n5413) );
  nand02 U2198 ( .Y(n5414), .A0(n5411), .A1(n5412) );
  inv01 U2199 ( .Y(n5404), .A(n5414) );
  ao22 U2200 ( .Y(n5415), .A0(larray[150]), .A1(n6974), .B0(larray[54]), .B1(
        n6970) );
  inv01 U2201 ( .Y(n5416), .A(n5415) );
  nand02 U2202 ( .Y(n7484), .A0(n5417), .A1(n5418) );
  inv01 U2203 ( .Y(n5419), .A(n6970) );
  inv01 U2204 ( .Y(n5420), .A(n6975) );
  inv01 U2205 ( .Y(n5421), .A(larray[153]) );
  inv01 U2206 ( .Y(n5422), .A(larray[57]) );
  nand02 U2207 ( .Y(n5423), .A0(n5419), .A1(n5420) );
  nand02 U2208 ( .Y(n5424), .A0(n5419), .A1(n5421) );
  nand02 U2209 ( .Y(n5425), .A0(n5420), .A1(n5422) );
  nand02 U2210 ( .Y(n5426), .A0(n5421), .A1(n5422) );
  nand02 U2211 ( .Y(n5427), .A0(n5423), .A1(n5424) );
  inv01 U2212 ( .Y(n5417), .A(n5427) );
  nand02 U2213 ( .Y(n5428), .A0(n5425), .A1(n5426) );
  inv01 U2214 ( .Y(n5418), .A(n5428) );
  ao22 U2215 ( .Y(n5429), .A0(larray[126]), .A1(n6975), .B0(larray[30]), .B1(
        n6970) );
  inv01 U2216 ( .Y(n5430), .A(n5429) );
  nand02 U2217 ( .Y(n7487), .A0(n5431), .A1(n5432) );
  inv01 U2218 ( .Y(n5433), .A(n6970) );
  inv01 U2219 ( .Y(n5434), .A(n6975) );
  inv01 U2220 ( .Y(n5435), .A(larray[147]) );
  inv01 U2221 ( .Y(n5436), .A(larray[51]) );
  nand02 U2222 ( .Y(n5437), .A0(n5433), .A1(n5434) );
  nand02 U2223 ( .Y(n5438), .A0(n5433), .A1(n5435) );
  nand02 U2224 ( .Y(n5439), .A0(n5434), .A1(n5436) );
  nand02 U2225 ( .Y(n5440), .A0(n5435), .A1(n5436) );
  nand02 U2226 ( .Y(n5441), .A0(n5437), .A1(n5438) );
  inv01 U2227 ( .Y(n5431), .A(n5441) );
  nand02 U2228 ( .Y(n5442), .A0(n5439), .A1(n5440) );
  inv01 U2229 ( .Y(n5432), .A(n5442) );
  nand02 U2230 ( .Y(n7478), .A0(n5443), .A1(n5444) );
  inv01 U2231 ( .Y(n5445), .A(n6971) );
  inv01 U2232 ( .Y(n5446), .A(n6975) );
  inv01 U2233 ( .Y(n5447), .A(larray[186]) );
  inv01 U2234 ( .Y(n5448), .A(larray[90]) );
  nand02 U2235 ( .Y(n5449), .A0(n5445), .A1(n5446) );
  nand02 U2236 ( .Y(n5450), .A0(n5445), .A1(n5447) );
  nand02 U2237 ( .Y(n5451), .A0(n5446), .A1(n5448) );
  nand02 U2238 ( .Y(n5452), .A0(n5447), .A1(n5448) );
  nand02 U2239 ( .Y(n5453), .A0(n5449), .A1(n5450) );
  inv01 U2240 ( .Y(n5443), .A(n5453) );
  nand02 U2241 ( .Y(n5454), .A0(n5451), .A1(n5452) );
  inv01 U2242 ( .Y(n5444), .A(n5454) );
  ao22 U2243 ( .Y(n5455), .A0(larray[180]), .A1(n6975), .B0(larray[84]), .B1(
        n6971) );
  inv01 U2244 ( .Y(n5456), .A(n5455) );
  nand02 U2245 ( .Y(n7508), .A0(n5457), .A1(n5458) );
  inv01 U2246 ( .Y(n5459), .A(n6971) );
  inv01 U2247 ( .Y(n5460), .A(n6974) );
  inv01 U2248 ( .Y(n5461), .A(larray[138]) );
  inv01 U2249 ( .Y(n5462), .A(larray[42]) );
  nand02 U2250 ( .Y(n5463), .A0(n5459), .A1(n5460) );
  nand02 U2251 ( .Y(n5464), .A0(n5459), .A1(n5461) );
  nand02 U2252 ( .Y(n5465), .A0(n5460), .A1(n5462) );
  nand02 U2253 ( .Y(n5466), .A0(n5461), .A1(n5462) );
  nand02 U2254 ( .Y(n5467), .A0(n5463), .A1(n5464) );
  inv01 U2255 ( .Y(n5457), .A(n5467) );
  nand02 U2256 ( .Y(n5468), .A0(n5465), .A1(n5466) );
  inv01 U2257 ( .Y(n5458), .A(n5468) );
  nand02 U2258 ( .Y(n7501), .A0(n5469), .A1(n5470) );
  inv01 U2259 ( .Y(n5471), .A(n6970) );
  inv01 U2260 ( .Y(n5472), .A(n6974) );
  inv01 U2261 ( .Y(n5473), .A(larray[129]) );
  inv01 U2262 ( .Y(n5474), .A(larray[33]) );
  nand02 U2263 ( .Y(n5475), .A0(n5471), .A1(n5472) );
  nand02 U2264 ( .Y(n5476), .A0(n5471), .A1(n5473) );
  nand02 U2265 ( .Y(n5477), .A0(n5472), .A1(n5474) );
  nand02 U2266 ( .Y(n5478), .A0(n5473), .A1(n5474) );
  nand02 U2267 ( .Y(n5479), .A0(n5475), .A1(n5476) );
  inv01 U2268 ( .Y(n5469), .A(n5479) );
  nand02 U2269 ( .Y(n5480), .A0(n5477), .A1(n5478) );
  inv01 U2270 ( .Y(n5470), .A(n5480) );
  nand02 U2271 ( .Y(n7510), .A0(n5481), .A1(n5482) );
  inv01 U2272 ( .Y(n5483), .A(n6970) );
  inv01 U2273 ( .Y(n5484), .A(n6974) );
  inv01 U2274 ( .Y(n5485), .A(larray[134]) );
  inv01 U2275 ( .Y(n5486), .A(larray[38]) );
  nand02 U2276 ( .Y(n5487), .A0(n5483), .A1(n5484) );
  nand02 U2277 ( .Y(n5488), .A0(n5483), .A1(n5485) );
  nand02 U2278 ( .Y(n5489), .A0(n5484), .A1(n5486) );
  nand02 U2279 ( .Y(n5490), .A0(n5485), .A1(n5486) );
  nand02 U2280 ( .Y(n5491), .A0(n5487), .A1(n5488) );
  inv01 U2281 ( .Y(n5481), .A(n5491) );
  nand02 U2282 ( .Y(n5492), .A0(n5489), .A1(n5490) );
  inv01 U2283 ( .Y(n5482), .A(n5492) );
  ao22 U2284 ( .Y(n5493), .A0(larray[106]), .A1(n6974), .B0(larray[10]), .B1(
        n6972) );
  inv01 U2285 ( .Y(n5494), .A(n5493) );
  nand02 U2286 ( .Y(n7506), .A0(n5495), .A1(n5496) );
  inv01 U2287 ( .Y(n5497), .A(n6972) );
  inv01 U2288 ( .Y(n5498), .A(n6974) );
  inv01 U2289 ( .Y(n5499), .A(larray[141]) );
  inv01 U2290 ( .Y(n5500), .A(larray[45]) );
  nand02 U2291 ( .Y(n5501), .A0(n5497), .A1(n5498) );
  nand02 U2292 ( .Y(n5502), .A0(n5497), .A1(n5499) );
  nand02 U2293 ( .Y(n5503), .A0(n5498), .A1(n5500) );
  nand02 U2294 ( .Y(n5504), .A0(n5499), .A1(n5500) );
  nand02 U2295 ( .Y(n5505), .A0(n5501), .A1(n5502) );
  inv01 U2296 ( .Y(n5495), .A(n5505) );
  nand02 U2297 ( .Y(n5506), .A0(n5503), .A1(n5504) );
  inv01 U2298 ( .Y(n5496), .A(n5506) );
  ao22 U2299 ( .Y(n5507), .A0(larray[172]), .A1(n6974), .B0(larray[76]), .B1(
        n6971) );
  inv01 U2300 ( .Y(n5508), .A(n5507) );
  nand02 U2301 ( .Y(n7498), .A0(n5509), .A1(n5510) );
  inv01 U2302 ( .Y(n5511), .A(n6970) );
  inv01 U2303 ( .Y(n5512), .A(n6975) );
  inv01 U2304 ( .Y(n5513), .A(larray[155]) );
  inv01 U2305 ( .Y(n5514), .A(larray[59]) );
  nand02 U2306 ( .Y(n5515), .A0(n5511), .A1(n5512) );
  nand02 U2307 ( .Y(n5516), .A0(n5511), .A1(n5513) );
  nand02 U2308 ( .Y(n5517), .A0(n5512), .A1(n5514) );
  nand02 U2309 ( .Y(n5518), .A0(n5513), .A1(n5514) );
  nand02 U2310 ( .Y(n5519), .A0(n5515), .A1(n5516) );
  inv01 U2311 ( .Y(n5509), .A(n5519) );
  nand02 U2312 ( .Y(n5520), .A0(n5517), .A1(n5518) );
  inv01 U2313 ( .Y(n5510), .A(n5520) );
  nand02 U2314 ( .Y(n7530), .A0(n5521), .A1(n5522) );
  inv01 U2315 ( .Y(n5523), .A(n6972) );
  inv01 U2316 ( .Y(n5524), .A(n6975) );
  inv01 U2317 ( .Y(n5525), .A(larray[109]) );
  inv01 U2318 ( .Y(n5526), .A(larray[13]) );
  nand02 U2319 ( .Y(n5527), .A0(n5523), .A1(n5524) );
  nand02 U2320 ( .Y(n5528), .A0(n5523), .A1(n5525) );
  nand02 U2321 ( .Y(n5529), .A0(n5524), .A1(n5526) );
  nand02 U2322 ( .Y(n5530), .A0(n5525), .A1(n5526) );
  nand02 U2323 ( .Y(n5531), .A0(n5527), .A1(n5528) );
  inv01 U2324 ( .Y(n5521), .A(n5531) );
  nand02 U2325 ( .Y(n5532), .A0(n5529), .A1(n5530) );
  inv01 U2326 ( .Y(n5522), .A(n5532) );
  ao22 U2327 ( .Y(n5533), .A0(larray[122]), .A1(n6975), .B0(larray[26]), .B1(
        n6972) );
  inv01 U2328 ( .Y(n5534), .A(n5533) );
  nand02 U2329 ( .Y(n7507), .A0(n5535), .A1(n5536) );
  inv01 U2330 ( .Y(n5537), .A(n6971) );
  inv01 U2331 ( .Y(n5538), .A(n6975) );
  inv01 U2332 ( .Y(n5539), .A(larray[140]) );
  inv01 U2333 ( .Y(n5540), .A(larray[44]) );
  nand02 U2334 ( .Y(n5541), .A0(n5537), .A1(n5538) );
  nand02 U2335 ( .Y(n5542), .A0(n5537), .A1(n5539) );
  nand02 U2336 ( .Y(n5543), .A0(n5538), .A1(n5540) );
  nand02 U2337 ( .Y(n5544), .A0(n5539), .A1(n5540) );
  nand02 U2338 ( .Y(n5545), .A0(n5541), .A1(n5542) );
  inv01 U2339 ( .Y(n5535), .A(n5545) );
  nand02 U2340 ( .Y(n5546), .A0(n5543), .A1(n5544) );
  inv01 U2341 ( .Y(n5536), .A(n5546) );
  ao22 U2342 ( .Y(n5547), .A0(larray[149]), .A1(n6975), .B0(larray[53]), .B1(
        n6972) );
  inv01 U2343 ( .Y(n5548), .A(n5547) );
  nand02 U2344 ( .Y(n7486), .A0(n5549), .A1(n5550) );
  inv01 U2345 ( .Y(n5551), .A(n6971) );
  inv01 U2346 ( .Y(n5552), .A(n6974) );
  inv01 U2347 ( .Y(n5553), .A(larray[148]) );
  inv01 U2348 ( .Y(n5554), .A(larray[52]) );
  nand02 U2349 ( .Y(n5555), .A0(n5551), .A1(n5552) );
  nand02 U2350 ( .Y(n5556), .A0(n5551), .A1(n5553) );
  nand02 U2351 ( .Y(n5557), .A0(n5552), .A1(n5554) );
  nand02 U2352 ( .Y(n5558), .A0(n5553), .A1(n5554) );
  nand02 U2353 ( .Y(n5559), .A0(n5555), .A1(n5556) );
  inv01 U2354 ( .Y(n5549), .A(n5559) );
  nand02 U2355 ( .Y(n5560), .A0(n5557), .A1(n5558) );
  inv01 U2356 ( .Y(n5550), .A(n5560) );
  nand02 U2357 ( .Y(n7476), .A0(n5561), .A1(n5562) );
  inv01 U2358 ( .Y(n5563), .A(n6970) );
  inv01 U2359 ( .Y(n5564), .A(n6974) );
  inv01 U2360 ( .Y(n5565), .A(larray[190]) );
  inv01 U2361 ( .Y(n5566), .A(larray[94]) );
  nand02 U2362 ( .Y(n5567), .A0(n5563), .A1(n5564) );
  nand02 U2363 ( .Y(n5568), .A0(n5563), .A1(n5565) );
  nand02 U2364 ( .Y(n5569), .A0(n5564), .A1(n5566) );
  nand02 U2365 ( .Y(n5570), .A0(n5565), .A1(n5566) );
  nand02 U2366 ( .Y(n5571), .A0(n5567), .A1(n5568) );
  inv01 U2367 ( .Y(n5561), .A(n5571) );
  nand02 U2368 ( .Y(n5572), .A0(n5569), .A1(n5570) );
  inv01 U2369 ( .Y(n5562), .A(n5572) );
  nand02 U2370 ( .Y(n7488), .A0(n5573), .A1(n5574) );
  inv01 U2371 ( .Y(n5575), .A(n6971) );
  inv01 U2372 ( .Y(n5576), .A(n6974) );
  inv01 U2373 ( .Y(n5577), .A(larray[167]) );
  inv01 U2374 ( .Y(n5578), .A(larray[71]) );
  nand02 U2375 ( .Y(n5579), .A0(n5575), .A1(n5576) );
  nand02 U2376 ( .Y(n5580), .A0(n5575), .A1(n5577) );
  nand02 U2377 ( .Y(n5581), .A0(n5576), .A1(n5578) );
  nand02 U2378 ( .Y(n5582), .A0(n5577), .A1(n5578) );
  nand02 U2379 ( .Y(n5583), .A0(n5579), .A1(n5580) );
  inv01 U2380 ( .Y(n5573), .A(n5583) );
  nand02 U2381 ( .Y(n5584), .A0(n5581), .A1(n5582) );
  inv01 U2382 ( .Y(n5574), .A(n5584) );
  ao22 U2383 ( .Y(n5585), .A0(larray[114]), .A1(n6974), .B0(larray[18]), .B1(
        n6971) );
  inv01 U2384 ( .Y(n5586), .A(n5585) );
  ao22 U2385 ( .Y(n5587), .A0(larray[105]), .A1(n6974), .B0(larray[9]), .B1(
        n6970) );
  inv01 U2386 ( .Y(n5588), .A(n5587) );
  nand02 U2387 ( .Y(n7475), .A0(n5589), .A1(n5590) );
  inv01 U2388 ( .Y(n5591), .A(n6972) );
  inv01 U2389 ( .Y(n5592), .A(n6974) );
  inv01 U2390 ( .Y(n5593), .A(larray[170]) );
  inv01 U2391 ( .Y(n5594), .A(larray[74]) );
  nand02 U2392 ( .Y(n5595), .A0(n5591), .A1(n5592) );
  nand02 U2393 ( .Y(n5596), .A0(n5591), .A1(n5593) );
  nand02 U2394 ( .Y(n5597), .A0(n5592), .A1(n5594) );
  nand02 U2395 ( .Y(n5598), .A0(n5593), .A1(n5594) );
  nand02 U2396 ( .Y(n5599), .A0(n5595), .A1(n5596) );
  inv01 U2397 ( .Y(n5589), .A(n5599) );
  nand02 U2398 ( .Y(n5600), .A0(n5597), .A1(n5598) );
  inv01 U2399 ( .Y(n5590), .A(n5600) );
  nand02 U2400 ( .Y(n7512), .A0(n5601), .A1(n5602) );
  inv01 U2401 ( .Y(n5603), .A(n6971) );
  inv01 U2402 ( .Y(n5604), .A(n6974) );
  inv01 U2403 ( .Y(n5605), .A(larray[132]) );
  inv01 U2404 ( .Y(n5606), .A(larray[36]) );
  nand02 U2405 ( .Y(n5607), .A0(n5603), .A1(n5604) );
  nand02 U2406 ( .Y(n5608), .A0(n5603), .A1(n5605) );
  nand02 U2407 ( .Y(n5609), .A0(n5604), .A1(n5606) );
  nand02 U2408 ( .Y(n5610), .A0(n5605), .A1(n5606) );
  nand02 U2409 ( .Y(n5611), .A0(n5607), .A1(n5608) );
  inv01 U2410 ( .Y(n5601), .A(n5611) );
  nand02 U2411 ( .Y(n5612), .A0(n5609), .A1(n5610) );
  inv01 U2412 ( .Y(n5602), .A(n5612) );
  ao22 U2413 ( .Y(n5613), .A0(larray[188]), .A1(n6974), .B0(larray[92]), .B1(
        n6971) );
  inv01 U2414 ( .Y(n5614), .A(n5613) );
  or02 U2415 ( .Y(n5615), .A0(n6986), .A1(n7233) );
  inv01 U2416 ( .Y(n5616), .A(n5615) );
  or02 U2417 ( .Y(n5617), .A0(n6986), .A1(n7260) );
  inv01 U2418 ( .Y(n5618), .A(n5617) );
  or02 U2419 ( .Y(n5619), .A0(n6986), .A1(n7230) );
  inv01 U2420 ( .Y(n5620), .A(n5619) );
  or02 U2421 ( .Y(n5621), .A0(n6987), .A1(n7292) );
  inv01 U2422 ( .Y(n5622), .A(n5621) );
  or02 U2423 ( .Y(n5623), .A0(n6987), .A1(n7259) );
  inv01 U2424 ( .Y(n5624), .A(n5623) );
  or02 U2425 ( .Y(n5625), .A0(n6986), .A1(n7365) );
  inv01 U2426 ( .Y(n5626), .A(n5625) );
  or02 U2427 ( .Y(n5627), .A0(n6986), .A1(n7296) );
  inv01 U2428 ( .Y(n5628), .A(n5627) );
  or02 U2429 ( .Y(n5629), .A0(n6986), .A1(n7293) );
  inv01 U2430 ( .Y(n5630), .A(n5629) );
  or02 U2431 ( .Y(n5631), .A0(n6986), .A1(n7326) );
  inv01 U2432 ( .Y(n5632), .A(n5631) );
  or02 U2433 ( .Y(n5633), .A0(n6986), .A1(n7359) );
  inv01 U2434 ( .Y(n5634), .A(n5633) );
  or02 U2435 ( .Y(n5635), .A0(n6987), .A1(n7226) );
  inv01 U2436 ( .Y(n5636), .A(n5635) );
  or02 U2437 ( .Y(n5637), .A0(n6987), .A1(n7229) );
  inv01 U2438 ( .Y(n5638), .A(n5637) );
  or02 U2439 ( .Y(n5639), .A0(n6987), .A1(n7358) );
  inv01 U2440 ( .Y(n5640), .A(n5639) );
  or02 U2441 ( .Y(n5641), .A0(n6987), .A1(n7262) );
  inv01 U2442 ( .Y(n5642), .A(n5641) );
  or02 U2443 ( .Y(n5643), .A0(n6986), .A1(n7263) );
  inv01 U2444 ( .Y(n5644), .A(n5643) );
  or02 U2445 ( .Y(n5645), .A0(n6986), .A1(n7227) );
  inv01 U2446 ( .Y(n5646), .A(n5645) );
  or02 U2447 ( .Y(n5647), .A0(n6986), .A1(n7356) );
  inv01 U2448 ( .Y(n5648), .A(n5647) );
  or02 U2449 ( .Y(n5649), .A0(n6986), .A1(n7362) );
  inv01 U2450 ( .Y(n5650), .A(n5649) );
  or02 U2451 ( .Y(n5651), .A0(n6987), .A1(n7355) );
  inv01 U2452 ( .Y(n5652), .A(n5651) );
  or02 U2453 ( .Y(n5653), .A0(n6987), .A1(n7361) );
  inv01 U2454 ( .Y(n5654), .A(n5653) );
  or02 U2455 ( .Y(n5655), .A0(n6987), .A1(n7289) );
  inv01 U2456 ( .Y(n5656), .A(n5655) );
  or02 U2457 ( .Y(n5657), .A0(n6987), .A1(n7223) );
  inv01 U2458 ( .Y(n5658), .A(n5657) );
  or02 U2459 ( .Y(n5659), .A0(n6986), .A1(n7329) );
  inv01 U2460 ( .Y(n5660), .A(n5659) );
  or02 U2461 ( .Y(n5661), .A0(n6986), .A1(n7299) );
  inv01 U2462 ( .Y(n5662), .A(n5661) );
  or02 U2463 ( .Y(n5663), .A0(n6986), .A1(n7290) );
  inv01 U2464 ( .Y(n5664), .A(n5663) );
  or02 U2465 ( .Y(n5665), .A0(n6986), .A1(n7224) );
  inv01 U2466 ( .Y(n5666), .A(n5665) );
  or02 U2467 ( .Y(n5667), .A0(n6984), .A1(n7034) );
  inv01 U2468 ( .Y(n5668), .A(n5667) );
  or02 U2469 ( .Y(n5669), .A0(n6984), .A1(n7097) );
  inv01 U2470 ( .Y(n5670), .A(n5669) );
  or02 U2471 ( .Y(n5671), .A0(n6987), .A1(n7298) );
  inv01 U2472 ( .Y(n5672), .A(n5671) );
  or02 U2473 ( .Y(n5673), .A0(n6987), .A1(n7325) );
  inv01 U2474 ( .Y(n5674), .A(n5673) );
  or02 U2475 ( .Y(n5675), .A0(n6987), .A1(n7232) );
  inv01 U2476 ( .Y(n5676), .A(n5675) );
  or02 U2477 ( .Y(n5677), .A0(n6987), .A1(n7364) );
  inv01 U2478 ( .Y(n5678), .A(n5677) );
  or02 U2479 ( .Y(n5679), .A0(n6987), .A1(n7295) );
  inv01 U2480 ( .Y(n5680), .A(n5679) );
  or02 U2481 ( .Y(n5681), .A0(n6987), .A1(n7328) );
  inv01 U2482 ( .Y(n5682), .A(n5681) );
  or02 U2483 ( .Y(n5683), .A0(n6984), .A1(n7121) );
  inv01 U2484 ( .Y(n5684), .A(n5683) );
  or02 U2485 ( .Y(n5685), .A0(n6984), .A1(n7079) );
  inv01 U2486 ( .Y(n5686), .A(n5685) );
  or02 U2487 ( .Y(n5687), .A0(n6984), .A1(n7037) );
  inv01 U2488 ( .Y(n5688), .A(n5687) );
  or02 U2489 ( .Y(n5689), .A0(n6984), .A1(n7115) );
  inv01 U2490 ( .Y(n5690), .A(n5689) );
  or02 U2491 ( .Y(n5691), .A0(n6984), .A1(n7031) );
  inv01 U2492 ( .Y(n5692), .A(n5691) );
  or02 U2493 ( .Y(n5693), .A0(n6984), .A1(n7028) );
  inv01 U2494 ( .Y(n5694), .A(n5693) );
  or02 U2495 ( .Y(n5695), .A0(n6984), .A1(n7094) );
  inv01 U2496 ( .Y(n5696), .A(n5695) );
  or02 U2497 ( .Y(n5697), .A0(n6984), .A1(n7112) );
  inv01 U2498 ( .Y(n5698), .A(n5697) );
  or02 U2499 ( .Y(n5699), .A0(n6984), .A1(n7055) );
  inv01 U2500 ( .Y(n5700), .A(n5699) );
  or02 U2501 ( .Y(n5701), .A0(n6984), .A1(n7118) );
  inv01 U2502 ( .Y(n5702), .A(n5701) );
  or02 U2503 ( .Y(n5703), .A0(n6984), .A1(n7070) );
  inv01 U2504 ( .Y(n5704), .A(n5703) );
  or02 U2505 ( .Y(n5705), .A0(n6984), .A1(n7052) );
  inv01 U2506 ( .Y(n5706), .A(n5705) );
  or02 U2507 ( .Y(n5707), .A0(n6984), .A1(n7076) );
  inv01 U2508 ( .Y(n5708), .A(n5707) );
  or02 U2509 ( .Y(n5709), .A0(n6984), .A1(n7073) );
  inv01 U2510 ( .Y(n5710), .A(n5709) );
  or02 U2511 ( .Y(n5711), .A0(n6982), .A1(n7075) );
  inv01 U2512 ( .Y(n5712), .A(n5711) );
  or02 U2513 ( .Y(n5713), .A0(n6982), .A1(n7033) );
  inv01 U2514 ( .Y(n5714), .A(n5713) );
  or02 U2515 ( .Y(n5715), .A0(n6982), .A1(n7114) );
  inv01 U2516 ( .Y(n5716), .A(n5715) );
  or02 U2517 ( .Y(n5717), .A0(n6982), .A1(n7099) );
  inv01 U2518 ( .Y(n5718), .A(n5717) );
  or02 U2519 ( .Y(n5719), .A0(n6982), .A1(n7081) );
  inv01 U2520 ( .Y(n5720), .A(n5719) );
  or02 U2521 ( .Y(n5721), .A0(n6982), .A1(n7054) );
  inv01 U2522 ( .Y(n5722), .A(n5721) );
  or02 U2523 ( .Y(n5723), .A0(n6982), .A1(n7078) );
  inv01 U2524 ( .Y(n5724), .A(n5723) );
  or02 U2525 ( .Y(n5725), .A0(n6982), .A1(n7057) );
  inv01 U2526 ( .Y(n5726), .A(n5725) );
  or02 U2527 ( .Y(n5727), .A0(n6982), .A1(n7072) );
  inv01 U2528 ( .Y(n5728), .A(n5727) );
  or02 U2529 ( .Y(n5729), .A0(n6982), .A1(n7039) );
  inv01 U2530 ( .Y(n5730), .A(n5729) );
  or02 U2531 ( .Y(n5731), .A0(n6982), .A1(n7120) );
  inv01 U2532 ( .Y(n5732), .A(n5731) );
  or02 U2533 ( .Y(n5733), .A0(n6982), .A1(n7036) );
  inv01 U2534 ( .Y(n5734), .A(n5733) );
  or02 U2535 ( .Y(n5735), .A0(n6982), .A1(n7117) );
  inv01 U2536 ( .Y(n5736), .A(n5735) );
  or02 U2537 ( .Y(n5737), .A0(n6982), .A1(n7030) );
  inv01 U2538 ( .Y(n5738), .A(n5737) );
  or02 U2539 ( .Y(n5739), .A0(n6982), .A1(n7096) );
  inv01 U2540 ( .Y(n5740), .A(n5739) );
  or02 U2541 ( .Y(n5741), .A0(n6982), .A1(n7123) );
  inv01 U2542 ( .Y(n5742), .A(n5741) );
  or02 U2543 ( .Y(n5743), .A0(n6988), .A1(n7294) );
  inv01 U2544 ( .Y(n5744), .A(n5743) );
  or02 U2545 ( .Y(n5745), .A0(n6988), .A1(n7291) );
  inv01 U2546 ( .Y(n5746), .A(n5745) );
  or02 U2547 ( .Y(n5747), .A0(n6988), .A1(n7231) );
  inv01 U2548 ( .Y(n5748), .A(n5747) );
  or02 U2549 ( .Y(n5749), .A0(n6988), .A1(n7327) );
  inv01 U2550 ( .Y(n5750), .A(n5749) );
  or02 U2551 ( .Y(n5751), .A0(n6983), .A1(n7032) );
  inv01 U2552 ( .Y(n5752), .A(n5751) );
  or02 U2553 ( .Y(n5753), .A0(n6983), .A1(n7056) );
  inv01 U2554 ( .Y(n5754), .A(n5753) );
  or02 U2555 ( .Y(n5755), .A0(n6983), .A1(n7053) );
  inv01 U2556 ( .Y(n5756), .A(n5755) );
  or02 U2557 ( .Y(n5757), .A0(n6988), .A1(n7324) );
  inv01 U2558 ( .Y(n5758), .A(n5757) );
  or02 U2559 ( .Y(n5759), .A0(n6988), .A1(n7357) );
  inv01 U2560 ( .Y(n5760), .A(n5759) );
  or02 U2561 ( .Y(n5761), .A0(n6988), .A1(n7228) );
  inv01 U2562 ( .Y(n5762), .A(n5761) );
  or02 U2563 ( .Y(n5763), .A0(n6988), .A1(n7363) );
  inv01 U2564 ( .Y(n5764), .A(n5763) );
  or02 U2565 ( .Y(n5765), .A0(n6983), .A1(n7077) );
  inv01 U2566 ( .Y(n5766), .A(n5765) );
  or02 U2567 ( .Y(n5767), .A0(n6983), .A1(n7080) );
  inv01 U2568 ( .Y(n5768), .A(n5767) );
  or02 U2569 ( .Y(n5769), .A0(n6983), .A1(n7035) );
  inv01 U2570 ( .Y(n5770), .A(n5769) );
  or02 U2571 ( .Y(n5771), .A0(n6988), .A1(n7360) );
  inv01 U2572 ( .Y(n5772), .A(n5771) );
  or02 U2573 ( .Y(n5773), .A0(n6988), .A1(n7288) );
  inv01 U2574 ( .Y(n5774), .A(n5773) );
  or02 U2575 ( .Y(n5775), .A0(n6988), .A1(n7354) );
  inv01 U2576 ( .Y(n5776), .A(n5775) );
  or02 U2577 ( .Y(n5777), .A0(n6988), .A1(n7258) );
  inv01 U2578 ( .Y(n5778), .A(n5777) );
  or02 U2579 ( .Y(n5779), .A0(n6983), .A1(n7113) );
  inv01 U2580 ( .Y(n5780), .A(n5779) );
  or02 U2581 ( .Y(n5781), .A0(n6983), .A1(n7074) );
  inv01 U2582 ( .Y(n5782), .A(n5781) );
  or02 U2583 ( .Y(n5783), .A0(n6983), .A1(n7122) );
  inv01 U2584 ( .Y(n5784), .A(n5783) );
  or02 U2585 ( .Y(n5785), .A0(n6988), .A1(n7222) );
  inv01 U2586 ( .Y(n5786), .A(n5785) );
  or02 U2587 ( .Y(n5787), .A0(n6988), .A1(n7225) );
  inv01 U2588 ( .Y(n5788), .A(n5787) );
  or02 U2589 ( .Y(n5789), .A0(n6988), .A1(n7261) );
  inv01 U2590 ( .Y(n5790), .A(n5789) );
  or02 U2591 ( .Y(n5791), .A0(n6988), .A1(n7297) );
  inv01 U2592 ( .Y(n5792), .A(n5791) );
  or02 U2593 ( .Y(n5793), .A0(n6983), .A1(n7098) );
  inv01 U2594 ( .Y(n5794), .A(n5793) );
  or02 U2595 ( .Y(n5795), .A0(n6983), .A1(n7095) );
  inv01 U2596 ( .Y(n5796), .A(n5795) );
  or02 U2597 ( .Y(n5797), .A0(n6983), .A1(n7119) );
  inv01 U2598 ( .Y(n5798), .A(n5797) );
  or02 U2599 ( .Y(n5799), .A0(n6983), .A1(n7071) );
  inv01 U2600 ( .Y(n5800), .A(n5799) );
  or02 U2601 ( .Y(n5801), .A0(n6983), .A1(n7029) );
  inv01 U2602 ( .Y(n5802), .A(n5801) );
  or02 U2603 ( .Y(n5803), .A0(n6983), .A1(n7038) );
  inv01 U2604 ( .Y(n5804), .A(n5803) );
  or02 U2605 ( .Y(n5805), .A0(n6983), .A1(n7116) );
  inv01 U2606 ( .Y(n5806), .A(n5805) );
  or02 U2607 ( .Y(n5807), .A0(s_state83), .A1(n4782) );
  inv01 U2608 ( .Y(n5808), .A(n5807) );
  or02 U2609 ( .Y(n5809), .A0(n6990), .A1(n7170) );
  inv01 U2610 ( .Y(n5810), .A(n5809) );
  or02 U2611 ( .Y(n5811), .A0(n6991), .A1(n7136) );
  inv01 U2612 ( .Y(n5812), .A(n5811) );
  or02 U2613 ( .Y(n5813), .A0(n6991), .A1(n7171) );
  inv01 U2614 ( .Y(n5814), .A(n5813) );
  or02 U2615 ( .Y(n5815), .A0(n6991), .A1(n7135) );
  inv01 U2616 ( .Y(n5816), .A(n5815) );
  or02 U2617 ( .Y(n5817), .A0(n6992), .A1(n7126) );
  inv01 U2618 ( .Y(n5818), .A(n5817) );
  or02 U2619 ( .Y(n5819), .A0(n6992), .A1(n7216) );
  inv01 U2620 ( .Y(n5820), .A(n5819) );
  or02 U2621 ( .Y(n5821), .A0(n6992), .A1(n7178) );
  inv01 U2622 ( .Y(n5822), .A(n5821) );
  or02 U2623 ( .Y(n5823), .A0(n6992), .A1(n7220) );
  inv01 U2624 ( .Y(n5824), .A(n5823) );
  or02 U2625 ( .Y(n5825), .A0(n6990), .A1(n7215) );
  inv01 U2626 ( .Y(n5826), .A(n5825) );
  or02 U2627 ( .Y(n5827), .A0(n6990), .A1(n7150) );
  inv01 U2628 ( .Y(n5828), .A(n5827) );
  or02 U2629 ( .Y(n5829), .A0(n6990), .A1(n7151) );
  inv01 U2630 ( .Y(n5830), .A(n5829) );
  or02 U2631 ( .Y(n5831), .A0(n6990), .A1(n7192) );
  inv01 U2632 ( .Y(n5832), .A(n5831) );
  or02 U2633 ( .Y(n5833), .A0(n6950), .A1(n7461) );
  inv01 U2634 ( .Y(n5834), .A(n5833) );
  or02 U2635 ( .Y(n5835), .A0(n6991), .A1(n7213) );
  inv01 U2636 ( .Y(n5836), .A(n5835) );
  or02 U2637 ( .Y(n5837), .A0(n6991), .A1(n7191) );
  inv01 U2638 ( .Y(n5838), .A(n5837) );
  or02 U2639 ( .Y(n5839), .A0(n6991), .A1(n7169) );
  inv01 U2640 ( .Y(n5840), .A(n5839) );
  or02 U2641 ( .Y(n5841), .A0(n6949), .A1(n7375) );
  inv01 U2642 ( .Y(n5842), .A(n5841) );
  or02 U2643 ( .Y(n5843), .A0(n6991), .A1(n7167) );
  inv01 U2644 ( .Y(n5844), .A(n5843) );
  or02 U2645 ( .Y(n5845), .A0(n6990), .A1(n7125) );
  inv01 U2646 ( .Y(n5846), .A(n5845) );
  or02 U2647 ( .Y(n5847), .A0(n6990), .A1(n7149) );
  inv01 U2648 ( .Y(n5848), .A(n5847) );
  or02 U2649 ( .Y(n5849), .A0(n6992), .A1(n7133) );
  inv01 U2650 ( .Y(n5850), .A(n5849) );
  or02 U2651 ( .Y(n5851), .A0(n6992), .A1(n7211) );
  inv01 U2652 ( .Y(n5852), .A(n5851) );
  or02 U2653 ( .Y(n5853), .A0(n6992), .A1(n7214) );
  inv01 U2654 ( .Y(n5854), .A(n5853) );
  or02 U2655 ( .Y(n5855), .A0(n6992), .A1(n7130) );
  inv01 U2656 ( .Y(n5856), .A(n5855) );
  or02 U2657 ( .Y(n5857), .A0(n6990), .A1(n7168) );
  inv01 U2658 ( .Y(n5858), .A(n5857) );
  or02 U2659 ( .Y(n5859), .A0(n6991), .A1(n7194) );
  inv01 U2660 ( .Y(n5860), .A(n5859) );
  or02 U2661 ( .Y(n5861), .A0(n6991), .A1(n7196) );
  inv01 U2662 ( .Y(n5862), .A(n5861) );
  or02 U2663 ( .Y(n5863), .A0(n6990), .A1(n7129) );
  inv01 U2664 ( .Y(n5864), .A(n5863) );
  or02 U2665 ( .Y(n5865), .A0(n6950), .A1(n7455) );
  inv01 U2666 ( .Y(n5866), .A(n5865) );
  or02 U2667 ( .Y(n5867), .A0(n6950), .A1(n7414) );
  inv01 U2668 ( .Y(n5868), .A(n5867) );
  or02 U2669 ( .Y(n5869), .A0(n6950), .A1(n7418) );
  inv01 U2670 ( .Y(n5870), .A(n5869) );
  or02 U2671 ( .Y(n5871), .A0(n6949), .A1(n7368) );
  inv01 U2672 ( .Y(n5872), .A(n5871) );
  or02 U2673 ( .Y(n5873), .A0(n6949), .A1(n7392) );
  inv01 U2674 ( .Y(n5874), .A(n5873) );
  or02 U2675 ( .Y(n5875), .A0(n6949), .A1(n7378) );
  inv01 U2676 ( .Y(n5876), .A(n5875) );
  or02 U2677 ( .Y(n5877), .A0(n6992), .A1(n7174) );
  inv01 U2678 ( .Y(n5878), .A(n5877) );
  or02 U2679 ( .Y(n5879), .A0(n6992), .A1(n7210) );
  inv01 U2680 ( .Y(n5880), .A(n5879) );
  or02 U2681 ( .Y(n5881), .A0(n6992), .A1(n7134) );
  inv01 U2682 ( .Y(n5882), .A(n5881) );
  or02 U2683 ( .Y(n5883), .A0(n6990), .A1(n7195) );
  inv01 U2684 ( .Y(n5884), .A(n5883) );
  or02 U2685 ( .Y(n5885), .A0(n6990), .A1(n7209) );
  inv01 U2686 ( .Y(n5886), .A(n5885) );
  or02 U2687 ( .Y(n5887), .A0(n6990), .A1(n7132) );
  inv01 U2688 ( .Y(n5888), .A(n5887) );
  or02 U2689 ( .Y(n5889), .A0(n6991), .A1(n7175) );
  inv01 U2690 ( .Y(n5890), .A(n5889) );
  or02 U2691 ( .Y(n5891), .A0(n6991), .A1(n7219) );
  inv01 U2692 ( .Y(n5892), .A(n5891) );
  or02 U2693 ( .Y(n5893), .A0(n6991), .A1(n7173) );
  inv01 U2694 ( .Y(n5894), .A(n5893) );
  or02 U2695 ( .Y(n5895), .A0(n6991), .A1(n7177) );
  inv01 U2696 ( .Y(n5896), .A(n5895) );
  or02 U2697 ( .Y(n5897), .A0(n6950), .A1(n7409) );
  inv01 U2698 ( .Y(n5898), .A(n5897) );
  or02 U2699 ( .Y(n5899), .A0(n6950), .A1(n7456) );
  inv01 U2700 ( .Y(n5900), .A(n5899) );
  or02 U2701 ( .Y(n5901), .A0(n6950), .A1(n7451) );
  inv01 U2702 ( .Y(n5902), .A(n5901) );
  or02 U2703 ( .Y(n5903), .A0(n6950), .A1(n7420) );
  inv01 U2704 ( .Y(n5904), .A(n5903) );
  or02 U2705 ( .Y(n5905), .A0(n6949), .A1(n7412) );
  inv01 U2706 ( .Y(n5906), .A(n5905) );
  or02 U2707 ( .Y(n5907), .A0(n6949), .A1(n7417) );
  inv01 U2708 ( .Y(n5908), .A(n5907) );
  or02 U2709 ( .Y(n5909), .A0(n6949), .A1(n7415) );
  inv01 U2710 ( .Y(n5910), .A(n5909) );
  or02 U2711 ( .Y(n5911), .A0(n6949), .A1(n7419) );
  inv01 U2712 ( .Y(n5912), .A(n5911) );
  or02 U2713 ( .Y(n5913), .A0(n6992), .A1(n7212) );
  inv01 U2714 ( .Y(n5914), .A(n5913) );
  or02 U2715 ( .Y(n5915), .A0(n6992), .A1(n7193) );
  inv01 U2716 ( .Y(n5916), .A(n5915) );
  or02 U2717 ( .Y(n5917), .A0(n6992), .A1(n7176) );
  inv01 U2718 ( .Y(n5918), .A(n5917) );
  or02 U2719 ( .Y(n5919), .A0(n6992), .A1(n7153) );
  inv01 U2720 ( .Y(n5920), .A(n5919) );
  or02 U2721 ( .Y(n5921), .A0(n6990), .A1(n7218) );
  inv01 U2722 ( .Y(n5922), .A(n5921) );
  or02 U2723 ( .Y(n5923), .A0(n6990), .A1(n7152) );
  inv01 U2724 ( .Y(n5924), .A(n5923) );
  or02 U2725 ( .Y(n5925), .A0(n6990), .A1(n7172) );
  inv01 U2726 ( .Y(n5926), .A(n5925) );
  or02 U2727 ( .Y(n5927), .A0(n6990), .A1(n7127) );
  inv01 U2728 ( .Y(n5928), .A(n5927) );
  or02 U2729 ( .Y(n5929), .A0(n6992), .A1(n7217) );
  inv01 U2730 ( .Y(n5930), .A(n5929) );
  or02 U2731 ( .Y(n5931), .A0(n6991), .A1(n7154) );
  inv01 U2732 ( .Y(n5932), .A(n5931) );
  or02 U2733 ( .Y(n5933), .A0(n6991), .A1(n7131) );
  inv01 U2734 ( .Y(n5934), .A(n5933) );
  or02 U2735 ( .Y(n5935), .A0(n6991), .A1(n7128) );
  inv01 U2736 ( .Y(n5936), .A(n5935) );
  or02 U2737 ( .Y(n5937), .A0(n6950), .A1(n7462) );
  inv01 U2738 ( .Y(n5938), .A(n5937) );
  or02 U2739 ( .Y(n5939), .A0(n6950), .A1(n7395) );
  inv01 U2740 ( .Y(n5940), .A(n5939) );
  or02 U2741 ( .Y(n5941), .A0(n6950), .A1(n7452) );
  inv01 U2742 ( .Y(n5942), .A(n5941) );
  or02 U2743 ( .Y(n5943), .A0(n6950), .A1(n7372) );
  inv01 U2744 ( .Y(n5944), .A(n5943) );
  or02 U2745 ( .Y(n5945), .A0(n6949), .A1(n7410) );
  inv01 U2746 ( .Y(n5946), .A(n5945) );
  or02 U2747 ( .Y(n5947), .A0(n6949), .A1(n7396) );
  inv01 U2748 ( .Y(n5948), .A(n5947) );
  or02 U2749 ( .Y(n5949), .A0(n6949), .A1(n7374) );
  inv01 U2750 ( .Y(n5950), .A(n5949) );
  or02 U2751 ( .Y(n5951), .A0(n6949), .A1(n7367) );
  inv01 U2752 ( .Y(n5952), .A(n5951) );
  or02 U2753 ( .Y(n5953), .A0(n6950), .A1(n7393) );
  inv01 U2754 ( .Y(n5954), .A(n5953) );
  or02 U2755 ( .Y(n5955), .A0(n6950), .A1(n7435) );
  inv01 U2756 ( .Y(n5956), .A(n5955) );
  or02 U2757 ( .Y(n5957), .A0(n6950), .A1(n7370) );
  inv01 U2758 ( .Y(n5958), .A(n5957) );
  or02 U2759 ( .Y(n5959), .A0(n6950), .A1(n7394) );
  inv01 U2760 ( .Y(n5960), .A(n5959) );
  or02 U2761 ( .Y(n5961), .A0(n6949), .A1(n7458) );
  inv01 U2762 ( .Y(n5962), .A(n5961) );
  or02 U2763 ( .Y(n5963), .A0(n6949), .A1(n7377) );
  inv01 U2764 ( .Y(n5964), .A(n5963) );
  or02 U2765 ( .Y(n5965), .A0(n6949), .A1(n7459) );
  inv01 U2766 ( .Y(n5966), .A(n5965) );
  or02 U2767 ( .Y(n5967), .A0(n6948), .A1(n7373) );
  inv01 U2768 ( .Y(n5968), .A(n5967) );
  or02 U2769 ( .Y(n5969), .A0(n6948), .A1(n7376) );
  inv01 U2770 ( .Y(n5970), .A(n5969) );
  or02 U2771 ( .Y(n5971), .A0(n6948), .A1(n7413) );
  inv01 U2772 ( .Y(n5972), .A(n5971) );
  or02 U2773 ( .Y(n5973), .A0(n6948), .A1(n7371) );
  inv01 U2774 ( .Y(n5974), .A(n5973) );
  or02 U2775 ( .Y(n5975), .A0(n6948), .A1(n7391) );
  inv01 U2776 ( .Y(n5976), .A(n5975) );
  or02 U2777 ( .Y(n5977), .A0(n6948), .A1(n7453) );
  inv01 U2778 ( .Y(n5978), .A(n5977) );
  or02 U2779 ( .Y(n5979), .A0(n6948), .A1(n7457) );
  inv01 U2780 ( .Y(n5980), .A(n5979) );
  or02 U2781 ( .Y(n5981), .A0(n6948), .A1(n7416) );
  inv01 U2782 ( .Y(n5982), .A(n5981) );
  or02 U2783 ( .Y(n5983), .A0(n6948), .A1(n7369) );
  inv01 U2784 ( .Y(n5984), .A(n5983) );
  or02 U2785 ( .Y(n5985), .A0(n6948), .A1(n7438) );
  inv01 U2786 ( .Y(n5986), .A(n5985) );
  or02 U2787 ( .Y(n5987), .A0(n6948), .A1(n7434) );
  inv01 U2788 ( .Y(n5988), .A(n5987) );
  or02 U2789 ( .Y(n5989), .A0(n6948), .A1(n7437) );
  inv01 U2790 ( .Y(n5990), .A(n5989) );
  or02 U2791 ( .Y(n5991), .A0(n6948), .A1(n7454) );
  inv01 U2792 ( .Y(n5992), .A(n5991) );
  or02 U2793 ( .Y(n5993), .A0(n6948), .A1(n7411) );
  inv01 U2794 ( .Y(n5994), .A(n5993) );
  or02 U2795 ( .Y(n5995), .A0(n6948), .A1(n7460) );
  inv01 U2796 ( .Y(n5996), .A(n5995) );
  or02 U2797 ( .Y(n5997), .A0(n6948), .A1(n7436) );
  inv01 U2798 ( .Y(n5998), .A(n5997) );
  or02 U2799 ( .Y(n5999), .A0(n6948), .A1(n7433) );
  inv01 U2800 ( .Y(n6000), .A(n5999) );
  nand02 U2801 ( .Y(n4744), .A0(n6001), .A1(n6002) );
  inv01 U2802 ( .Y(n6003), .A(n6997) );
  inv01 U2803 ( .Y(n6004), .A(n4214) );
  inv01 U2804 ( .Y(n6005), .A(n6951) );
  nand02 U2805 ( .Y(n6001), .A0(n6951), .A1(n6003) );
  nand02 U2806 ( .Y(n6002), .A0(n6004), .A1(n6005) );
  nand02 U2807 ( .Y(n4696), .A0(n6006), .A1(n6007) );
  inv01 U2808 ( .Y(n6008), .A(n6997) );
  inv01 U2809 ( .Y(n6009), .A(n4262) );
  inv01 U2810 ( .Y(n6010), .A(n6954) );
  nand02 U2811 ( .Y(n6006), .A0(n6954), .A1(n6008) );
  nand02 U2812 ( .Y(n6007), .A0(n6009), .A1(n6010) );
  buf02 U2813 ( .Y(n6011), .A(n4720) );
  inv01 U2814 ( .Y(n4768), .A(n6012) );
  inv01 U2815 ( .Y(n6013), .A(n6953) );
  nor02 U2816 ( .Y(n6014), .A0(n6997), .A1(n6013) );
  nor02 U2817 ( .Y(n6015), .A0(n6953), .A1(n4190) );
  nor02 U2818 ( .Y(n6012), .A0(n6014), .A1(n6015) );
  inv02 U2819 ( .Y(n6997), .A(n____return2214_0_) );
  buf02 U2820 ( .Y(n6016), .A(n4693) );
  nand02 U2821 ( .Y(n4746), .A0(n6017), .A1(n6018) );
  inv01 U2822 ( .Y(n6019), .A(n7020) );
  inv01 U2823 ( .Y(n6020), .A(n4204) );
  inv01 U2824 ( .Y(n6021), .A(n6953) );
  nand02 U2825 ( .Y(n6017), .A0(n6953), .A1(n6019) );
  nand02 U2826 ( .Y(n6018), .A0(n6020), .A1(n6021) );
  buf02 U2827 ( .Y(n6022), .A(n4722) );
  buf02 U2828 ( .Y(n6023), .A(n4692) );
  buf02 U2829 ( .Y(n6024), .A(n4707) );
  buf02 U2830 ( .Y(n6025), .A(n4677) );
  nand02 U2831 ( .Y(n4767), .A0(n6026), .A1(n6027) );
  inv01 U2832 ( .Y(n6028), .A(n6999) );
  inv01 U2833 ( .Y(n6029), .A(n4201) );
  inv01 U2834 ( .Y(n6030), .A(n6953) );
  nand02 U2835 ( .Y(n6026), .A0(n6953), .A1(n6028) );
  nand02 U2836 ( .Y(n6027), .A0(n6029), .A1(n6030) );
  buf02 U2837 ( .Y(n6031), .A(n4719) );
  buf02 U2838 ( .Y(n6032), .A(n4705) );
  buf02 U2839 ( .Y(n6033), .A(n4702) );
  buf02 U2840 ( .Y(n6034), .A(n4738) );
  buf02 U2841 ( .Y(n6035), .A(n4755) );
  buf02 U2842 ( .Y(n6036), .A(n4691) );
  buf02 U2843 ( .Y(n6037), .A(n4699) );
  buf02 U2844 ( .Y(n6038), .A(n4700) );
  buf02 U2845 ( .Y(n6039), .A(n4703) );
  buf02 U2846 ( .Y(n6040), .A(n4676) );
  buf02 U2847 ( .Y(n6041), .A(n4731) );
  buf02 U2848 ( .Y(n6042), .A(n4752) );
  buf02 U2849 ( .Y(n6043), .A(n4749) );
  buf02 U2850 ( .Y(n6044), .A(n4730) );
  buf02 U2851 ( .Y(n6045), .A(n4766) );
  nand02 U2852 ( .Y(n4708), .A0(n6046), .A1(n6047) );
  inv01 U2853 ( .Y(n6048), .A(n7010) );
  inv01 U2854 ( .Y(n6049), .A(n4241) );
  inv01 U2855 ( .Y(n6050), .A(n6952) );
  nand02 U2856 ( .Y(n6046), .A0(n6952), .A1(n6048) );
  nand02 U2857 ( .Y(n6047), .A0(n6049), .A1(n6050) );
  buf02 U2858 ( .Y(n6051), .A(n4684) );
  buf02 U2859 ( .Y(n6052), .A(n4727) );
  buf02 U2860 ( .Y(n6053), .A(n4740) );
  buf02 U2861 ( .Y(n6054), .A(n4736) );
  buf02 U2862 ( .Y(n6055), .A(n4757) );
  buf02 U2863 ( .Y(n6056), .A(n4747) );
  buf02 U2864 ( .Y(n6057), .A(n4763) );
  buf02 U2865 ( .Y(n6058), .A(n4713) );
  buf02 U2866 ( .Y(n6059), .A(n4735) );
  buf02 U2867 ( .Y(n6060), .A(n4737) );
  buf02 U2868 ( .Y(n6061), .A(n4734) );
  buf02 U2869 ( .Y(n6062), .A(n4681) );
  buf02 U2870 ( .Y(n6063), .A(n4706) );
  buf02 U2871 ( .Y(n6064), .A(n4675) );
  buf02 U2872 ( .Y(n6065), .A(n4712) );
  buf02 U2873 ( .Y(n6066), .A(n4711) );
  buf02 U2874 ( .Y(n6067), .A(n4751) );
  buf02 U2875 ( .Y(n6068), .A(n4716) );
  buf02 U2876 ( .Y(n6069), .A(n4688) );
  buf02 U2877 ( .Y(n6070), .A(n4748) );
  buf02 U2878 ( .Y(n6071), .A(n4742) );
  buf02 U2879 ( .Y(n6072), .A(n4750) );
  buf02 U2880 ( .Y(n6073), .A(n4709) );
  buf02 U2881 ( .Y(n6074), .A(n4759) );
  buf02 U2882 ( .Y(n6075), .A(n4690) );
  buf02 U2883 ( .Y(n6076), .A(n4678) );
  buf02 U2884 ( .Y(n6077), .A(n4714) );
  buf02 U2885 ( .Y(n6078), .A(n4729) );
  buf02 U2886 ( .Y(n6079), .A(n4756) );
  buf02 U2887 ( .Y(n6080), .A(n4754) );
  buf02 U2888 ( .Y(n6081), .A(n4726) );
  buf02 U2889 ( .Y(n6082), .A(n4686) );
  buf02 U2890 ( .Y(n6083), .A(n4764) );
  nand02 U2891 ( .Y(n4717), .A0(n6084), .A1(n6085) );
  inv01 U2892 ( .Y(n6086), .A(n7001) );
  inv01 U2893 ( .Y(n6087), .A(n4255) );
  inv01 U2894 ( .Y(n6088), .A(n6952) );
  nand02 U2895 ( .Y(n6084), .A0(n6952), .A1(n6086) );
  nand02 U2896 ( .Y(n6085), .A0(n6087), .A1(n6088) );
  buf02 U2897 ( .Y(n6089), .A(n4710) );
  buf02 U2898 ( .Y(n6090), .A(n4765) );
  buf02 U2899 ( .Y(n6091), .A(n4687) );
  buf02 U2900 ( .Y(n6092), .A(n4715) );
  buf02 U2901 ( .Y(n6093), .A(n4679) );
  buf02 U2902 ( .Y(n6094), .A(n4741) );
  buf02 U2903 ( .Y(n6095), .A(n4743) );
  buf02 U2904 ( .Y(n6096), .A(n4701) );
  buf02 U2905 ( .Y(n6097), .A(n4723) );
  buf02 U2906 ( .Y(n6098), .A(n4704) );
  buf02 U2907 ( .Y(n6099), .A(n4760) );
  buf02 U2908 ( .Y(n6100), .A(n4733) );
  buf02 U2909 ( .Y(n6101), .A(n4694) );
  buf02 U2910 ( .Y(n6102), .A(n4725) );
  buf02 U2911 ( .Y(n6103), .A(n4762) );
  buf02 U2912 ( .Y(n6104), .A(n4680) );
  buf02 U2913 ( .Y(n6105), .A(n4682) );
  buf02 U2914 ( .Y(n6106), .A(n4724) );
  buf02 U2915 ( .Y(n6107), .A(n4761) );
  buf02 U2916 ( .Y(n6108), .A(n4683) );
  buf02 U2917 ( .Y(n6109), .A(n4695) );
  buf02 U2918 ( .Y(n6110), .A(n4718) );
  buf02 U2919 ( .Y(n6111), .A(n4753) );
  buf02 U2920 ( .Y(n6112), .A(n4685) );
  buf02 U2921 ( .Y(n6113), .A(n4739) );
  buf02 U2922 ( .Y(n6114), .A(n4689) );
  buf02 U2923 ( .Y(n6115), .A(n4728) );
  buf02 U2924 ( .Y(n6116), .A(n4732) );
  buf02 U2925 ( .Y(n6117), .A(n4758) );
  nand02 U2926 ( .Y(n4745), .A0(n6118), .A1(n6119) );
  inv01 U2927 ( .Y(n6120), .A(n7021) );
  inv01 U2928 ( .Y(n6121), .A(n4205) );
  inv01 U2929 ( .Y(n6122), .A(n6953) );
  nand02 U2930 ( .Y(n6118), .A0(n6953), .A1(n6120) );
  nand02 U2931 ( .Y(n6119), .A0(n6121), .A1(n6122) );
  nand02 U2932 ( .Y(n4697), .A0(n6123), .A1(n6124) );
  inv01 U2933 ( .Y(n6125), .A(n7021) );
  inv01 U2934 ( .Y(n6126), .A(n4253) );
  inv01 U2935 ( .Y(n6127), .A(n6952) );
  nand02 U2936 ( .Y(n6123), .A0(n6952), .A1(n6125) );
  nand02 U2937 ( .Y(n6124), .A0(n6126), .A1(n6127) );
  buf02 U2938 ( .Y(n6128), .A(n4673) );
  nand02 U2939 ( .Y(n4674), .A0(n6129), .A1(n6130) );
  inv01 U2940 ( .Y(n6131), .A(n7020) );
  inv01 U2941 ( .Y(n6132), .A(n4276) );
  inv01 U2942 ( .Y(n6133), .A(n6954) );
  nand02 U2943 ( .Y(n6129), .A0(n6954), .A1(n6131) );
  nand02 U2944 ( .Y(n6130), .A0(n6132), .A1(n6133) );
  buf02 U2945 ( .Y(n6134), .A(n4698) );
  buf02 U2946 ( .Y(n6135), .A(n4721) );
  buf02 U2947 ( .Y(n6136), .A(n4371) );
  buf02 U2948 ( .Y(n6137), .A(n4329) );
  buf02 U2949 ( .Y(n6138), .A(n4353) );
  buf02 U2950 ( .Y(n6139), .A(n4425) );
  buf02 U2951 ( .Y(n6140), .A(n4467) );
  buf02 U2952 ( .Y(n6141), .A(n4407) );
  buf02 U2953 ( .Y(n6142), .A(n4449) );
  buf02 U2954 ( .Y(n6143), .A(n4311) );
  buf02 U2955 ( .Y(n6144), .A(n4319) );
  buf02 U2956 ( .Y(n6145), .A(n4439) );
  nand02 U2957 ( .Y(n4301), .A0(n6146), .A1(n6147) );
  inv01 U2958 ( .Y(n6148), .A(n7353) );
  inv01 U2959 ( .Y(n6149), .A(n7450) );
  inv01 U2960 ( .Y(n6150), .A(n6949) );
  nand02 U2961 ( .Y(n6146), .A0(n6949), .A1(n6148) );
  nand02 U2962 ( .Y(n6147), .A0(n6149), .A1(n6150) );
  buf02 U2963 ( .Y(n6151), .A(n4397) );
  nand02 U2964 ( .Y(n4361), .A0(n6152), .A1(n6153) );
  inv01 U2965 ( .Y(n6154), .A(n7257) );
  inv01 U2966 ( .Y(n6155), .A(n7390) );
  inv01 U2967 ( .Y(n6156), .A(n6949) );
  nand02 U2968 ( .Y(n6152), .A0(n6949), .A1(n6154) );
  nand02 U2969 ( .Y(n6153), .A0(n6155), .A1(n6156) );
  buf02 U2970 ( .Y(n6157), .A(n4457) );
  buf02 U2971 ( .Y(n6158), .A(n4415) );
  buf02 U2972 ( .Y(n6159), .A(n4343) );
  nand02 U2973 ( .Y(n4328), .A0(n6160), .A1(n6161) );
  inv01 U2974 ( .Y(n6162), .A(n7305) );
  inv01 U2975 ( .Y(n6163), .A(n7423) );
  inv01 U2976 ( .Y(n6164), .A(n6948) );
  nand02 U2977 ( .Y(n6160), .A0(n6948), .A1(n6162) );
  nand02 U2978 ( .Y(n6161), .A0(n6163), .A1(n6164) );
  buf02 U2979 ( .Y(n6165), .A(n4424) );
  buf02 U2980 ( .Y(n6166), .A(n4369) );
  buf02 U2981 ( .Y(n6167), .A(n4370) );
  buf02 U2982 ( .Y(n6168), .A(n4465) );
  nand02 U2983 ( .Y(n4404), .A0(n6169), .A1(n6170) );
  inv01 U2984 ( .Y(n6171), .A(n7339) );
  inv01 U2985 ( .Y(n6172), .A(n7338) );
  inv01 U2986 ( .Y(n6173), .A(n6987) );
  nand02 U2987 ( .Y(n6169), .A0(n6987), .A1(n6171) );
  nand02 U2988 ( .Y(n6170), .A0(n6172), .A1(n6173) );
  buf02 U2989 ( .Y(n6174), .A(n4308) );
  buf02 U2990 ( .Y(n6175), .A(n4310) );
  buf02 U2991 ( .Y(n6176), .A(n4406) );
  nand02 U2992 ( .Y(n4448), .A0(n6177), .A1(n6178) );
  inv01 U2993 ( .Y(n6179), .A(n7269) );
  inv01 U2994 ( .Y(n6180), .A(n7268) );
  inv01 U2995 ( .Y(n6181), .A(n6986) );
  nand02 U2996 ( .Y(n6177), .A0(n6986), .A1(n6179) );
  nand02 U2997 ( .Y(n6178), .A0(n6180), .A1(n6181) );
  buf02 U2998 ( .Y(n6182), .A(n4352) );
  buf02 U2999 ( .Y(n6183), .A(n4466) );
  buf02 U3000 ( .Y(n6184), .A(n4345) );
  buf02 U3001 ( .Y(n6185), .A(n4346) );
  buf02 U3002 ( .Y(n6186), .A(n4323) );
  buf02 U3003 ( .Y(n6187), .A(n4447) );
  nand02 U3004 ( .Y(n4401), .A0(n6188), .A1(n6189) );
  inv01 U3005 ( .Y(n6190), .A(n7345) );
  inv01 U3006 ( .Y(n6191), .A(n7344) );
  inv01 U3007 ( .Y(n6192), .A(n6987) );
  nand02 U3008 ( .Y(n6188), .A0(n6987), .A1(n6190) );
  nand02 U3009 ( .Y(n6189), .A0(n6191), .A1(n6192) );
  buf02 U3010 ( .Y(n6193), .A(n4398) );
  buf02 U3011 ( .Y(n6194), .A(n4326) );
  buf02 U3012 ( .Y(n6195), .A(n4305) );
  buf02 U3013 ( .Y(n6196), .A(n4309) );
  buf02 U3014 ( .Y(n6197), .A(n4304) );
  buf02 U3015 ( .Y(n6198), .A(n4327) );
  buf02 U3016 ( .Y(n6199), .A(n4417) );
  buf02 U3017 ( .Y(n6200), .A(n4303) );
  buf02 U3018 ( .Y(n6201), .A(n4344) );
  buf02 U3019 ( .Y(n6202), .A(n4460) );
  buf02 U3020 ( .Y(n6203), .A(n4462) );
  buf02 U3021 ( .Y(n6204), .A(n4420) );
  buf02 U3022 ( .Y(n6205), .A(n4320) );
  buf02 U3023 ( .Y(n6206), .A(n4459) );
  buf02 U3024 ( .Y(n6207), .A(n4351) );
  buf02 U3025 ( .Y(n6208), .A(n4441) );
  buf02 U3026 ( .Y(n6209), .A(n4362) );
  nand02 U3027 ( .Y(n4463), .A0(n6210), .A1(n6211) );
  inv01 U3028 ( .Y(n6212), .A(n7245) );
  inv01 U3029 ( .Y(n6213), .A(n7244) );
  inv01 U3030 ( .Y(n6214), .A(n6986) );
  nand02 U3031 ( .Y(n6210), .A0(n6986), .A1(n6212) );
  nand02 U3032 ( .Y(n6211), .A0(n6213), .A1(n6214) );
  buf02 U3033 ( .Y(n6215), .A(n4367) );
  buf02 U3034 ( .Y(n6216), .A(n4402) );
  nand02 U3035 ( .Y(n4421), .A0(n6217), .A1(n6218) );
  inv01 U3036 ( .Y(n6219), .A(n7311) );
  inv01 U3037 ( .Y(n6220), .A(n7310) );
  inv01 U3038 ( .Y(n6221), .A(n6986) );
  nand02 U3039 ( .Y(n6217), .A0(n6986), .A1(n6219) );
  nand02 U3040 ( .Y(n6218), .A0(n6220), .A1(n6221) );
  buf02 U3041 ( .Y(n6222), .A(n4325) );
  buf02 U3042 ( .Y(n6223), .A(n4418) );
  buf02 U3043 ( .Y(n6224), .A(n4348) );
  buf02 U3044 ( .Y(n6225), .A(n4364) );
  buf02 U3045 ( .Y(n6226), .A(n4322) );
  buf02 U3046 ( .Y(n6227), .A(n4307) );
  buf02 U3047 ( .Y(n6228), .A(n4405) );
  buf02 U3048 ( .Y(n6229), .A(n4423) );
  buf02 U3049 ( .Y(n6230), .A(n4349) );
  buf02 U3050 ( .Y(n6231), .A(n4324) );
  buf02 U3051 ( .Y(n6232), .A(n4302) );
  buf02 U3052 ( .Y(n6233), .A(n4445) );
  buf02 U3053 ( .Y(n6234), .A(n4366) );
  buf02 U3054 ( .Y(n6235), .A(n4458) );
  buf02 U3055 ( .Y(n6236), .A(n4363) );
  buf02 U3056 ( .Y(n6237), .A(n4442) );
  buf02 U3057 ( .Y(n6238), .A(n4440) );
  buf02 U3058 ( .Y(n6239), .A(n4365) );
  nand02 U3059 ( .Y(n4350), .A0(n6240), .A1(n6241) );
  inv01 U3060 ( .Y(n6242), .A(n7273) );
  inv01 U3061 ( .Y(n6243), .A(n7401) );
  inv01 U3062 ( .Y(n6244), .A(n6950) );
  nand02 U3063 ( .Y(n6240), .A0(n6950), .A1(n6242) );
  nand02 U3064 ( .Y(n6241), .A0(n6243), .A1(n6244) );
  buf02 U3065 ( .Y(n6245), .A(n4347) );
  buf02 U3066 ( .Y(n6246), .A(n4446) );
  buf02 U3067 ( .Y(n6247), .A(n4321) );
  buf02 U3068 ( .Y(n6248), .A(n4461) );
  buf02 U3069 ( .Y(n6249), .A(n4464) );
  buf02 U3070 ( .Y(n6250), .A(n4399) );
  buf02 U3071 ( .Y(n6251), .A(n4403) );
  buf02 U3072 ( .Y(n6252), .A(n4416) );
  buf02 U3073 ( .Y(n6253), .A(n4444) );
  buf02 U3074 ( .Y(n6254), .A(n4422) );
  buf02 U3075 ( .Y(n6255), .A(n4443) );
  buf02 U3076 ( .Y(n6256), .A(n4368) );
  buf02 U3077 ( .Y(n6257), .A(n4419) );
  buf02 U3078 ( .Y(n6258), .A(n4400) );
  buf02 U3079 ( .Y(n6259), .A(n4306) );
  nand02 U3080 ( .Y(n4330), .A0(n6260), .A1(n6261) );
  inv01 U3081 ( .Y(n6262), .A(n7301) );
  inv01 U3082 ( .Y(n6263), .A(n7421) );
  inv01 U3083 ( .Y(n6264), .A(n6948) );
  nand02 U3084 ( .Y(n6260), .A0(n6948), .A1(n6262) );
  nand02 U3085 ( .Y(n6261), .A0(n6263), .A1(n6264) );
  buf02 U3086 ( .Y(n6265), .A(n4372) );
  buf02 U3087 ( .Y(n6266), .A(n4354) );
  buf02 U3088 ( .Y(n6267), .A(n4426) );
  nand02 U3089 ( .Y(n4408), .A0(n6268), .A1(n6269) );
  inv01 U3090 ( .Y(n6270), .A(n7331) );
  inv01 U3091 ( .Y(n6271), .A(n7330) );
  inv01 U3092 ( .Y(n6272), .A(n6988) );
  nand02 U3093 ( .Y(n6268), .A0(n6988), .A1(n6270) );
  nand02 U3094 ( .Y(n6269), .A0(n6271), .A1(n6272) );
  buf02 U3095 ( .Y(n6273), .A(n4450) );
  buf02 U3096 ( .Y(n6274), .A(n4312) );
  buf02 U3097 ( .Y(n6275), .A(n4468) );
  inv12 U3098 ( .Y(n6992), .A(n6989) );
  inv12 U3099 ( .Y(n6991), .A(n6989) );
  inv12 U3100 ( .Y(n6990), .A(n6989) );
  xor2 U3101 ( .Y(n6276), .A0(s_signb_i), .A1(n3535) );
  inv01 U3102 ( .Y(sign_o), .A(n6276) );
  or02 U3103 ( .Y(n6278), .A0(n6958), .A1(n7025) );
  inv01 U3104 ( .Y(n6279), .A(n6278) );
  or02 U3105 ( .Y(n6280), .A0(n6965), .A1(n7025) );
  inv01 U3106 ( .Y(n6281), .A(n6280) );
  ao22 U3107 ( .Y(n6282), .A0(n7468), .A1(n6946), .B0(n7469), .B1(n7221) );
  inv01 U3108 ( .Y(n6283), .A(n6282) );
  ao22 U3109 ( .Y(n6284), .A0(n7466), .A1(n6940), .B0(n7467), .B1(n7366) );
  inv01 U3110 ( .Y(n6285), .A(n6284) );
  inv04 U3111 ( .Y(n6957), .A(n7024) );
  or03 U3112 ( .Y(n6286), .A0(n6942), .A1(n6936), .A2(n6946) );
  inv01 U3113 ( .Y(n6287), .A(n6286) );
  inv01 U3114 ( .Y(n7027), .A(n6288) );
  inv01 U3115 ( .Y(n6289), .A(n6944) );
  inv01 U3116 ( .Y(n6290), .A(n6936) );
  inv01 U3117 ( .Y(n6291), .A(n6940) );
  nand02 U3118 ( .Y(n6288), .A0(n6291), .A1(n6292) );
  nand02 U3119 ( .Y(n6293), .A0(n6289), .A1(n6290) );
  inv01 U3120 ( .Y(n6292), .A(n6293) );
  buf02 U3121 ( .Y(n6944), .A(count_0_) );
  or03 U3122 ( .Y(n6294), .A0(n6946), .A1(n6936), .A2(n7366) );
  inv01 U3123 ( .Y(n6295), .A(n6294) );
  inv01 U3124 ( .Y(n6985), .A(n6296) );
  inv01 U3125 ( .Y(n6297), .A(n7366) );
  inv01 U3126 ( .Y(n6298), .A(n6936) );
  inv01 U3127 ( .Y(n6299), .A(n6943) );
  nand02 U3128 ( .Y(n6296), .A0(n6299), .A1(n6300) );
  nand02 U3129 ( .Y(n6301), .A0(n6297), .A1(n6298) );
  inv01 U3130 ( .Y(n6300), .A(n6301) );
  buf02 U3131 ( .Y(n6943), .A(count_0_) );
  or02 U3132 ( .Y(n6302), .A0(n6995), .A1(s_state83) );
  inv02 U3133 ( .Y(n6303), .A(n6302) );
  or02 U3134 ( .Y(n6304), .A0(n6995), .A1(n6982) );
  inv02 U3135 ( .Y(n6305), .A(n6304) );
  or02 U3136 ( .Y(n6306), .A0(n6938), .A1(n6946) );
  inv02 U3137 ( .Y(n6307), .A(n6306) );
  inv02 U3138 ( .Y(member2137_3__9_), .A(n6308) );
  nor02 U3139 ( .Y(n6309), .A0(n6958), .A1(n7348) );
  nor02 U3140 ( .Y(n6310), .A0(n6965), .A1(n7448) );
  inv01 U3141 ( .Y(n6311), .A(n7470) );
  nor02 U3142 ( .Y(n6308), .A0(n6311), .A1(n6312) );
  nor02 U3143 ( .Y(n6313), .A0(n6309), .A1(n6310) );
  inv01 U3144 ( .Y(n6312), .A(n6313) );
  inv02 U3145 ( .Y(member2137_3__10_), .A(n6314) );
  nor02 U3146 ( .Y(n6315), .A0(n6962), .A1(n7350) );
  nor02 U3147 ( .Y(n6316), .A0(n6967), .A1(n7449) );
  inv01 U3148 ( .Y(n6317), .A(n5362) );
  nor02 U3149 ( .Y(n6314), .A0(n6317), .A1(n6318) );
  nor02 U3150 ( .Y(n6319), .A0(n6315), .A1(n6316) );
  inv01 U3151 ( .Y(n6318), .A(n6319) );
  inv02 U3152 ( .Y(member2137_3__23_), .A(n6320) );
  nor02 U3153 ( .Y(n6321), .A0(n6960), .A1(n7365) );
  nor02 U3154 ( .Y(n6322), .A0(n6966), .A1(n7462) );
  inv01 U3155 ( .Y(n6323), .A(n4808) );
  nor02 U3156 ( .Y(n6320), .A0(n6323), .A1(n6324) );
  nor02 U3157 ( .Y(n6325), .A0(n6321), .A1(n6322) );
  inv01 U3158 ( .Y(n6324), .A(n6325) );
  inv02 U3159 ( .Y(member2137_3__1_), .A(n6326) );
  nor02 U3160 ( .Y(n6327), .A0(n6958), .A1(n7332) );
  nor02 U3161 ( .Y(n6328), .A0(n6965), .A1(n7440) );
  inv01 U3162 ( .Y(n6329), .A(n4846) );
  nor02 U3163 ( .Y(n6326), .A0(n6329), .A1(n6330) );
  nor02 U3164 ( .Y(n6331), .A0(n6327), .A1(n6328) );
  inv01 U3165 ( .Y(n6330), .A(n6331) );
  inv02 U3166 ( .Y(member2137_3__16_), .A(n6332) );
  nor02 U3167 ( .Y(n6333), .A0(n6962), .A1(n7358) );
  nor02 U3168 ( .Y(n6334), .A0(n6967), .A1(n7455) );
  inv01 U3169 ( .Y(n6335), .A(n7479) );
  nor02 U3170 ( .Y(n6332), .A0(n6335), .A1(n6336) );
  nor02 U3171 ( .Y(n6337), .A0(n6333), .A1(n6334) );
  inv01 U3172 ( .Y(n6336), .A(n6337) );
  inv02 U3173 ( .Y(member2137_3__18_), .A(n6338) );
  nor02 U3174 ( .Y(n6339), .A0(n6960), .A1(n7360) );
  nor02 U3175 ( .Y(n6340), .A0(n6966), .A1(n7457) );
  inv01 U3176 ( .Y(n6341), .A(n7478) );
  nor02 U3177 ( .Y(n6338), .A0(n6341), .A1(n6342) );
  nor02 U3178 ( .Y(n6343), .A0(n6339), .A1(n6340) );
  inv01 U3179 ( .Y(n6342), .A(n6343) );
  inv02 U3180 ( .Y(member2137_3__12_), .A(n6344) );
  nor02 U3181 ( .Y(n6345), .A0(n6960), .A1(n7354) );
  nor02 U3182 ( .Y(n6346), .A0(n6966), .A1(n7451) );
  inv01 U3183 ( .Y(n6347), .A(n5456) );
  nor02 U3184 ( .Y(n6344), .A0(n6347), .A1(n6348) );
  nor02 U3185 ( .Y(n6349), .A0(n6345), .A1(n6346) );
  inv01 U3186 ( .Y(n6348), .A(n6349) );
  inv02 U3187 ( .Y(member2137_3__21_), .A(n6350) );
  nor02 U3188 ( .Y(n6351), .A0(n6962), .A1(n7363) );
  nor02 U3189 ( .Y(n6352), .A0(n6967), .A1(n7460) );
  inv01 U3190 ( .Y(n6353), .A(n4886) );
  nor02 U3191 ( .Y(n6350), .A0(n6353), .A1(n6354) );
  nor02 U3192 ( .Y(n6355), .A0(n6351), .A1(n6352) );
  inv01 U3193 ( .Y(n6354), .A(n6355) );
  inv02 U3194 ( .Y(member2137_3__5_), .A(n6356) );
  nor02 U3195 ( .Y(n6357), .A0(n6962), .A1(n7340) );
  nor02 U3196 ( .Y(n6358), .A0(n6967), .A1(n7444) );
  inv01 U3197 ( .Y(n6359), .A(n7473) );
  nor02 U3198 ( .Y(n6356), .A0(n6359), .A1(n6360) );
  nor02 U3199 ( .Y(n6361), .A0(n6357), .A1(n6358) );
  inv01 U3200 ( .Y(n6360), .A(n6361) );
  inv02 U3201 ( .Y(member2137_3__7_), .A(n6362) );
  nor02 U3202 ( .Y(n6363), .A0(n6960), .A1(n7344) );
  nor02 U3203 ( .Y(n6364), .A0(n6966), .A1(n7446) );
  inv01 U3204 ( .Y(n6365), .A(n5284) );
  nor02 U3205 ( .Y(n6362), .A0(n6365), .A1(n6366) );
  nor02 U3206 ( .Y(n6367), .A0(n6363), .A1(n6364) );
  inv01 U3207 ( .Y(n6366), .A(n6367) );
  inv02 U3208 ( .Y(member2137_3__14_), .A(n6368) );
  nor02 U3209 ( .Y(n6369), .A0(n6958), .A1(n7356) );
  nor02 U3210 ( .Y(n6370), .A0(n6965), .A1(n7453) );
  inv01 U3211 ( .Y(n6371), .A(n5026) );
  nor02 U3212 ( .Y(n6368), .A0(n6371), .A1(n6372) );
  nor02 U3213 ( .Y(n6373), .A0(n6369), .A1(n6370) );
  inv01 U3214 ( .Y(n6372), .A(n6373) );
  inv02 U3215 ( .Y(member2137_3__3_), .A(n6374) );
  nor02 U3216 ( .Y(n6375), .A0(n6958), .A1(n7336) );
  nor02 U3217 ( .Y(n6376), .A0(n6965), .A1(n7442) );
  inv01 U3218 ( .Y(n6377), .A(n7474) );
  nor02 U3219 ( .Y(n6374), .A0(n6377), .A1(n6378) );
  nor02 U3220 ( .Y(n6379), .A0(n6375), .A1(n6376) );
  inv01 U3221 ( .Y(n6378), .A(n6379) );
  inv02 U3222 ( .Y(member2137_3__15_), .A(n6380) );
  nor02 U3223 ( .Y(n6381), .A0(n6960), .A1(n7357) );
  nor02 U3224 ( .Y(n6382), .A0(n6966), .A1(n7454) );
  inv01 U3225 ( .Y(n6383), .A(n7480) );
  nor02 U3226 ( .Y(n6380), .A0(n6383), .A1(n6384) );
  nor02 U3227 ( .Y(n6385), .A0(n6381), .A1(n6382) );
  inv01 U3228 ( .Y(n6384), .A(n6385) );
  inv02 U3229 ( .Y(member2137_3__17_), .A(n6386) );
  nor02 U3230 ( .Y(n6387), .A0(n6958), .A1(n7359) );
  nor02 U3231 ( .Y(n6388), .A0(n6965), .A1(n7456) );
  inv01 U3232 ( .Y(n6389), .A(n5258) );
  nor02 U3233 ( .Y(n6386), .A0(n6389), .A1(n6390) );
  nor02 U3234 ( .Y(n6391), .A0(n6387), .A1(n6388) );
  inv01 U3235 ( .Y(n6390), .A(n6391) );
  inv02 U3236 ( .Y(member2137_3__2_), .A(n6392) );
  nor02 U3237 ( .Y(n6393), .A0(n6962), .A1(n7334) );
  nor02 U3238 ( .Y(n6394), .A0(n6967), .A1(n7441) );
  inv01 U3239 ( .Y(n6395), .A(n7475) );
  nor02 U3240 ( .Y(n6392), .A0(n6395), .A1(n6396) );
  nor02 U3241 ( .Y(n6397), .A0(n6393), .A1(n6394) );
  inv01 U3242 ( .Y(n6396), .A(n6397) );
  inv02 U3243 ( .Y(member1883_1__22_), .A(n6398) );
  nor02 U3244 ( .Y(n6399), .A0(n6958), .A1(n7292) );
  nor02 U3245 ( .Y(n6400), .A0(n6965), .A1(n7413) );
  inv01 U3246 ( .Y(n6401), .A(n7505) );
  nor02 U3247 ( .Y(n6398), .A0(n6401), .A1(n6402) );
  nor02 U3248 ( .Y(n6403), .A0(n6399), .A1(n6400) );
  inv01 U3249 ( .Y(n6402), .A(n6403) );
  inv02 U3250 ( .Y(member2137_3__22_), .A(n6404) );
  nor02 U3251 ( .Y(n6405), .A0(n6958), .A1(n7364) );
  nor02 U3252 ( .Y(n6406), .A0(n6965), .A1(n7461) );
  inv01 U3253 ( .Y(n6407), .A(n7476) );
  nor02 U3254 ( .Y(n6404), .A0(n6407), .A1(n6408) );
  nor02 U3255 ( .Y(n6409), .A0(n6405), .A1(n6406) );
  inv01 U3256 ( .Y(n6408), .A(n6409) );
  inv02 U3257 ( .Y(member2137_3__4_), .A(n6410) );
  nor02 U3258 ( .Y(n6411), .A0(n6960), .A1(n7338) );
  nor02 U3259 ( .Y(n6412), .A0(n6966), .A1(n7443) );
  inv01 U3260 ( .Y(n6413), .A(n5508) );
  nor02 U3261 ( .Y(n6410), .A0(n6413), .A1(n6414) );
  nor02 U3262 ( .Y(n6415), .A0(n6411), .A1(n6412) );
  inv01 U3263 ( .Y(n6414), .A(n6415) );
  inv02 U3264 ( .Y(member2137_3__20_), .A(n6416) );
  nor02 U3265 ( .Y(n6417), .A0(n6960), .A1(n7362) );
  nor02 U3266 ( .Y(n6418), .A0(n6966), .A1(n7459) );
  inv01 U3267 ( .Y(n6419), .A(n5614) );
  nor02 U3268 ( .Y(n6416), .A0(n6419), .A1(n6420) );
  nor02 U3269 ( .Y(n6421), .A0(n6417), .A1(n6418) );
  inv01 U3270 ( .Y(n6420), .A(n6421) );
  inv02 U3271 ( .Y(member1883_1__23_), .A(n6422) );
  nor02 U3272 ( .Y(n6423), .A0(n6960), .A1(n7293) );
  nor02 U3273 ( .Y(n6424), .A0(n6966), .A1(n7414) );
  inv01 U3274 ( .Y(n6425), .A(n7504) );
  nor02 U3275 ( .Y(n6422), .A0(n6425), .A1(n6426) );
  nor02 U3276 ( .Y(n6427), .A0(n6423), .A1(n6424) );
  inv01 U3277 ( .Y(n6426), .A(n6427) );
  inv02 U3278 ( .Y(member2137_3__13_), .A(n6428) );
  nor02 U3279 ( .Y(n6429), .A0(n6962), .A1(n7355) );
  nor02 U3280 ( .Y(n6430), .A0(n6967), .A1(n7452) );
  inv01 U3281 ( .Y(n6431), .A(n7481) );
  nor02 U3282 ( .Y(n6428), .A0(n6431), .A1(n6432) );
  nor02 U3283 ( .Y(n6433), .A0(n6429), .A1(n6430) );
  inv01 U3284 ( .Y(n6432), .A(n6433) );
  inv02 U3285 ( .Y(member2137_3__8_), .A(n6434) );
  nor02 U3286 ( .Y(n6435), .A0(n6962), .A1(n7346) );
  nor02 U3287 ( .Y(n6436), .A0(n6967), .A1(n7447) );
  inv01 U3288 ( .Y(n6437), .A(n7471) );
  nor02 U3289 ( .Y(n6434), .A0(n6437), .A1(n6438) );
  nor02 U3290 ( .Y(n6439), .A0(n6435), .A1(n6436) );
  inv01 U3291 ( .Y(n6438), .A(n6439) );
  inv02 U3292 ( .Y(member2137_3__19_), .A(n6440) );
  nor02 U3293 ( .Y(n6441), .A0(n6962), .A1(n7361) );
  nor02 U3294 ( .Y(n6442), .A0(n6967), .A1(n7458) );
  inv01 U3295 ( .Y(n6443), .A(n7477) );
  nor02 U3296 ( .Y(n6440), .A0(n6443), .A1(n6444) );
  nor02 U3297 ( .Y(n6445), .A0(n6441), .A1(n6442) );
  inv01 U3298 ( .Y(n6444), .A(n6445) );
  inv02 U3299 ( .Y(member1883_1__21_), .A(n6446) );
  nor02 U3300 ( .Y(n6447), .A0(n6962), .A1(n7291) );
  nor02 U3301 ( .Y(n6448), .A0(n6967), .A1(n7412) );
  inv01 U3302 ( .Y(n6449), .A(n7506) );
  nor02 U3303 ( .Y(n6446), .A0(n6449), .A1(n6450) );
  nor02 U3304 ( .Y(n6451), .A0(n6447), .A1(n6448) );
  inv01 U3305 ( .Y(n6450), .A(n6451) );
  inv02 U3306 ( .Y(member2137_3__6_), .A(n6452) );
  nor02 U3307 ( .Y(n6453), .A0(n6958), .A1(n7342) );
  nor02 U3308 ( .Y(n6454), .A0(n6965), .A1(n7445) );
  inv01 U3309 ( .Y(n6455), .A(n7472) );
  nor02 U3310 ( .Y(n6452), .A0(n6455), .A1(n6456) );
  nor02 U3311 ( .Y(n6457), .A0(n6453), .A1(n6454) );
  inv01 U3312 ( .Y(n6456), .A(n6457) );
  inv02 U3313 ( .Y(member2137_3__11_), .A(n6458) );
  nor02 U3314 ( .Y(n6459), .A0(n6958), .A1(n7352) );
  nor02 U3315 ( .Y(n6460), .A0(n6965), .A1(n7450) );
  inv01 U3316 ( .Y(n6461), .A(n7482) );
  nor02 U3317 ( .Y(n6458), .A0(n6461), .A1(n6462) );
  nor02 U3318 ( .Y(n6463), .A0(n6459), .A1(n6460) );
  inv01 U3319 ( .Y(n6462), .A(n6463) );
  inv02 U3320 ( .Y(member1883_1__20_), .A(n6464) );
  nor02 U3321 ( .Y(n6465), .A0(n6960), .A1(n7290) );
  nor02 U3322 ( .Y(n6466), .A0(n6966), .A1(n7411) );
  inv01 U3323 ( .Y(n6467), .A(n7507) );
  nor02 U3324 ( .Y(n6464), .A0(n6467), .A1(n6468) );
  nor02 U3325 ( .Y(n6469), .A0(n6465), .A1(n6466) );
  inv01 U3326 ( .Y(n6468), .A(n6469) );
  inv02 U3327 ( .Y(member1883_1__18_), .A(n6470) );
  nor02 U3328 ( .Y(n6471), .A0(n6960), .A1(n7288) );
  nor02 U3329 ( .Y(n6472), .A0(n6966), .A1(n7409) );
  inv01 U3330 ( .Y(n6473), .A(n7508) );
  nor02 U3331 ( .Y(n6470), .A0(n6473), .A1(n6474) );
  nor02 U3332 ( .Y(n6475), .A0(n6471), .A1(n6472) );
  inv01 U3333 ( .Y(n6474), .A(n6475) );
  inv02 U3334 ( .Y(member1883_1__19_), .A(n6476) );
  nor02 U3335 ( .Y(n6477), .A0(n6962), .A1(n7289) );
  nor02 U3336 ( .Y(n6478), .A0(n6967), .A1(n7410) );
  inv01 U3337 ( .Y(n6479), .A(n4950) );
  nor02 U3338 ( .Y(n6476), .A0(n6479), .A1(n6480) );
  nor02 U3339 ( .Y(n6481), .A0(n6477), .A1(n6478) );
  inv01 U3340 ( .Y(n6480), .A(n6481) );
  inv02 U3341 ( .Y(member1883_1__16_), .A(n6482) );
  nor02 U3342 ( .Y(n6483), .A0(n6962), .A1(n7284) );
  nor02 U3343 ( .Y(n6484), .A0(n6967), .A1(n7407) );
  inv01 U3344 ( .Y(n6485), .A(n7509) );
  nor02 U3345 ( .Y(n6482), .A0(n6485), .A1(n6486) );
  nor02 U3346 ( .Y(n6487), .A0(n6483), .A1(n6484) );
  inv01 U3347 ( .Y(n6486), .A(n6487) );
  inv02 U3348 ( .Y(member1883_1__17_), .A(n6488) );
  nor02 U3349 ( .Y(n6489), .A0(n6958), .A1(n7286) );
  nor02 U3350 ( .Y(n6490), .A0(n6965), .A1(n7408) );
  inv01 U3351 ( .Y(n6491), .A(n5402) );
  nor02 U3352 ( .Y(n6488), .A0(n6491), .A1(n6492) );
  nor02 U3353 ( .Y(n6493), .A0(n6489), .A1(n6490) );
  inv01 U3354 ( .Y(n6492), .A(n6493) );
  inv02 U3355 ( .Y(member1883_1__14_), .A(n6494) );
  nor02 U3356 ( .Y(n6495), .A0(n6958), .A1(n7280) );
  nor02 U3357 ( .Y(n6496), .A0(n6965), .A1(n7405) );
  inv01 U3358 ( .Y(n6497), .A(n7510) );
  nor02 U3359 ( .Y(n6494), .A0(n6497), .A1(n6498) );
  nor02 U3360 ( .Y(n6499), .A0(n6495), .A1(n6496) );
  inv01 U3361 ( .Y(n6498), .A(n6499) );
  inv02 U3362 ( .Y(member1883_1__15_), .A(n6500) );
  nor02 U3363 ( .Y(n6501), .A0(n6960), .A1(n7282) );
  nor02 U3364 ( .Y(n6502), .A0(n6966), .A1(n7406) );
  inv01 U3365 ( .Y(n6503), .A(n5090) );
  nor02 U3366 ( .Y(n6500), .A0(n6503), .A1(n6504) );
  nor02 U3367 ( .Y(n6505), .A0(n6501), .A1(n6502) );
  inv01 U3368 ( .Y(n6504), .A(n6505) );
  inv02 U3369 ( .Y(member1883_1__12_), .A(n6506) );
  nor02 U3370 ( .Y(n6507), .A0(n6960), .A1(n7276) );
  nor02 U3371 ( .Y(n6508), .A0(n6966), .A1(n7403) );
  inv01 U3372 ( .Y(n6509), .A(n7512) );
  nor02 U3373 ( .Y(n6506), .A0(n6509), .A1(n6510) );
  nor02 U3374 ( .Y(n6511), .A0(n6507), .A1(n6508) );
  inv01 U3375 ( .Y(n6510), .A(n6511) );
  inv02 U3376 ( .Y(member1883_1__13_), .A(n6512) );
  nor02 U3377 ( .Y(n6513), .A0(n6962), .A1(n7278) );
  nor02 U3378 ( .Y(n6514), .A0(n6967), .A1(n7404) );
  inv01 U3379 ( .Y(n6515), .A(n7511) );
  nor02 U3380 ( .Y(n6512), .A0(n6515), .A1(n6516) );
  nor02 U3381 ( .Y(n6517), .A0(n6513), .A1(n6514) );
  inv01 U3382 ( .Y(n6516), .A(n6517) );
  inv02 U3383 ( .Y(member1883_1__10_), .A(n6518) );
  nor02 U3384 ( .Y(n6519), .A0(n6962), .A1(n7272) );
  nor02 U3385 ( .Y(n6520), .A0(n6967), .A1(n7401) );
  inv01 U3386 ( .Y(n6521), .A(n7514) );
  nor02 U3387 ( .Y(n6518), .A0(n6521), .A1(n6522) );
  nor02 U3388 ( .Y(n6523), .A0(n6519), .A1(n6520) );
  inv01 U3389 ( .Y(n6522), .A(n6523) );
  inv02 U3390 ( .Y(member1883_1__11_), .A(n6524) );
  nor02 U3391 ( .Y(n6525), .A0(n6958), .A1(n7274) );
  nor02 U3392 ( .Y(n6526), .A0(n6965), .A1(n7402) );
  inv01 U3393 ( .Y(n6527), .A(n7513) );
  nor02 U3394 ( .Y(n6524), .A0(n6527), .A1(n6528) );
  nor02 U3395 ( .Y(n6529), .A0(n6525), .A1(n6526) );
  inv01 U3396 ( .Y(n6528), .A(n6529) );
  inv02 U3397 ( .Y(member1883_1__9_), .A(n6530) );
  nor02 U3398 ( .Y(n6531), .A0(n6958), .A1(n7270) );
  nor02 U3399 ( .Y(n6532), .A0(n6965), .A1(n7400) );
  inv01 U3400 ( .Y(n6533), .A(n7501) );
  nor02 U3401 ( .Y(n6530), .A0(n6533), .A1(n6534) );
  nor02 U3402 ( .Y(n6535), .A0(n6531), .A1(n6532) );
  inv01 U3403 ( .Y(n6534), .A(n6535) );
  inv02 U3404 ( .Y(member1883_1__8_), .A(n6536) );
  nor02 U3405 ( .Y(n6537), .A0(n6962), .A1(n7268) );
  nor02 U3406 ( .Y(n6538), .A0(n6967), .A1(n7399) );
  inv01 U3407 ( .Y(n6539), .A(n7502) );
  nor02 U3408 ( .Y(n6536), .A0(n6539), .A1(n6540) );
  nor02 U3409 ( .Y(n6541), .A0(n6537), .A1(n6538) );
  inv01 U3410 ( .Y(n6540), .A(n6541) );
  inv02 U3411 ( .Y(member1883_1__7_), .A(n6542) );
  nor02 U3412 ( .Y(n6543), .A0(n6960), .A1(n7266) );
  nor02 U3413 ( .Y(n6544), .A0(n6966), .A1(n7398) );
  inv01 U3414 ( .Y(n6545), .A(n5180) );
  nor02 U3415 ( .Y(n6542), .A0(n6545), .A1(n6546) );
  nor02 U3416 ( .Y(n6547), .A0(n6543), .A1(n6544) );
  inv01 U3417 ( .Y(n6546), .A(n6547) );
  inv02 U3418 ( .Y(member1883_1__6_), .A(n6548) );
  nor02 U3419 ( .Y(n6549), .A0(n6958), .A1(n7264) );
  nor02 U3420 ( .Y(n6550), .A0(n6965), .A1(n7397) );
  inv01 U3421 ( .Y(n6551), .A(n5430) );
  nor02 U3422 ( .Y(n6548), .A0(n6551), .A1(n6552) );
  nor02 U3423 ( .Y(n6553), .A0(n6549), .A1(n6550) );
  inv01 U3424 ( .Y(n6552), .A(n6553) );
  inv02 U3425 ( .Y(member1883_1__5_), .A(n6554) );
  nor02 U3426 ( .Y(n6555), .A0(n6962), .A1(n7263) );
  nor02 U3427 ( .Y(n6556), .A0(n6967), .A1(n7396) );
  inv01 U3428 ( .Y(n6557), .A(n5322) );
  nor02 U3429 ( .Y(n6554), .A0(n6557), .A1(n6558) );
  nor02 U3430 ( .Y(n6559), .A0(n6555), .A1(n6556) );
  inv01 U3431 ( .Y(n6558), .A(n6559) );
  inv02 U3432 ( .Y(member1883_1__4_), .A(n6560) );
  nor02 U3433 ( .Y(n6561), .A0(n6960), .A1(n7262) );
  nor02 U3434 ( .Y(n6562), .A0(n6966), .A1(n7395) );
  inv01 U3435 ( .Y(n6563), .A(n7503) );
  nor02 U3436 ( .Y(n6560), .A0(n6563), .A1(n6564) );
  nor02 U3437 ( .Y(n6565), .A0(n6561), .A1(n6562) );
  inv01 U3438 ( .Y(n6564), .A(n6565) );
  inv02 U3439 ( .Y(member1883_1__3_), .A(n6566) );
  nor02 U3440 ( .Y(n6567), .A0(n6958), .A1(n7261) );
  nor02 U3441 ( .Y(n6568), .A0(n6965), .A1(n7394) );
  inv01 U3442 ( .Y(n6569), .A(n4988) );
  nor02 U3443 ( .Y(n6566), .A0(n6569), .A1(n6570) );
  nor02 U3444 ( .Y(n6571), .A0(n6567), .A1(n6568) );
  inv01 U3445 ( .Y(n6570), .A(n6571) );
  inv02 U3446 ( .Y(member1883_1__2_), .A(n6572) );
  nor02 U3447 ( .Y(n6573), .A0(n6962), .A1(n7260) );
  nor02 U3448 ( .Y(n6574), .A0(n6967), .A1(n7393) );
  inv01 U3449 ( .Y(n6575), .A(n5534) );
  nor02 U3450 ( .Y(n6572), .A0(n6575), .A1(n6576) );
  nor02 U3451 ( .Y(n6577), .A0(n6573), .A1(n6574) );
  inv01 U3452 ( .Y(n6576), .A(n6577) );
  inv02 U3453 ( .Y(member1883_1__1_), .A(n6578) );
  nor02 U3454 ( .Y(n6579), .A0(n6958), .A1(n7259) );
  nor02 U3455 ( .Y(n6580), .A0(n6965), .A1(n7392) );
  inv01 U3456 ( .Y(n6581), .A(n5064) );
  nor02 U3457 ( .Y(n6578), .A0(n6581), .A1(n6582) );
  nor02 U3458 ( .Y(n6583), .A0(n6579), .A1(n6580) );
  inv01 U3459 ( .Y(n6582), .A(n6583) );
  inv02 U3460 ( .Y(member2010_2__11_), .A(n6584) );
  nor02 U3461 ( .Y(n6585), .A0(n6958), .A1(n7310) );
  nor02 U3462 ( .Y(n6586), .A0(n6965), .A1(n7426) );
  inv01 U3463 ( .Y(n6587), .A(n7498) );
  nor02 U3464 ( .Y(n6584), .A0(n6587), .A1(n6588) );
  nor02 U3465 ( .Y(n6589), .A0(n6585), .A1(n6586) );
  inv01 U3466 ( .Y(n6588), .A(n6589) );
  inv02 U3467 ( .Y(member2010_2__12_), .A(n6590) );
  nor02 U3468 ( .Y(n6591), .A0(n6960), .A1(n7312) );
  nor02 U3469 ( .Y(n6592), .A0(n6966), .A1(n7427) );
  inv01 U3470 ( .Y(n6593), .A(n7497) );
  nor02 U3471 ( .Y(n6590), .A0(n6593), .A1(n6594) );
  nor02 U3472 ( .Y(n6595), .A0(n6591), .A1(n6592) );
  inv01 U3473 ( .Y(n6594), .A(n6595) );
  inv02 U3474 ( .Y(member1796_0__16_), .A(n6596) );
  nor02 U3475 ( .Y(n6597), .A0(n6962), .A1(n7242) );
  nor02 U3476 ( .Y(n6598), .A0(n6967), .A1(n7383) );
  inv01 U3477 ( .Y(n6599), .A(n5206) );
  nor02 U3478 ( .Y(n6596), .A0(n6599), .A1(n6600) );
  nor02 U3479 ( .Y(n6601), .A0(n6597), .A1(n6598) );
  inv01 U3480 ( .Y(n6600), .A(n6601) );
  inv02 U3481 ( .Y(member2010_2__4_), .A(n6602) );
  nor02 U3482 ( .Y(n6603), .A0(n6960), .A1(n7298) );
  nor02 U3483 ( .Y(n6604), .A0(n6966), .A1(n7419) );
  inv01 U3484 ( .Y(n6605), .A(n7486) );
  nor02 U3485 ( .Y(n6602), .A0(n6605), .A1(n6606) );
  nor02 U3486 ( .Y(n6607), .A0(n6603), .A1(n6604) );
  inv01 U3487 ( .Y(n6606), .A(n6607) );
  inv02 U3488 ( .Y(member2010_2__6_), .A(n6608) );
  nor02 U3489 ( .Y(n6609), .A0(n6958), .A1(n7300) );
  nor02 U3490 ( .Y(n6610), .A0(n6965), .A1(n7421) );
  inv01 U3491 ( .Y(n6611), .A(n5416) );
  nor02 U3492 ( .Y(n6608), .A0(n6611), .A1(n6612) );
  nor02 U3493 ( .Y(n6613), .A0(n6609), .A1(n6610) );
  inv01 U3494 ( .Y(n6612), .A(n6613) );
  inv02 U3495 ( .Y(member2010_2__23_), .A(n6614) );
  nor02 U3496 ( .Y(n6615), .A0(n6960), .A1(n7329) );
  nor02 U3497 ( .Y(n6616), .A0(n6966), .A1(n7438) );
  inv01 U3498 ( .Y(n6617), .A(n7488) );
  nor02 U3499 ( .Y(n6614), .A0(n6617), .A1(n6618) );
  nor02 U3500 ( .Y(n6619), .A0(n6615), .A1(n6616) );
  inv01 U3501 ( .Y(n6618), .A(n6619) );
  inv02 U3502 ( .Y(member1796_0__23_), .A(n6620) );
  nor02 U3503 ( .Y(n6621), .A0(n6960), .A1(n7256) );
  nor02 U3504 ( .Y(n6622), .A0(n6966), .A1(n7390) );
  inv01 U3505 ( .Y(n6623), .A(n7523) );
  nor02 U3506 ( .Y(n6620), .A0(n6623), .A1(n6624) );
  nor02 U3507 ( .Y(n6625), .A0(n6621), .A1(n6622) );
  inv01 U3508 ( .Y(n6624), .A(n6625) );
  inv02 U3509 ( .Y(member1796_0__6_), .A(n6626) );
  nor02 U3510 ( .Y(n6627), .A0(n6958), .A1(n7228) );
  nor02 U3511 ( .Y(n6628), .A0(n6965), .A1(n7373) );
  inv01 U3512 ( .Y(n6629), .A(n7518) );
  nor02 U3513 ( .Y(n6626), .A0(n6629), .A1(n6630) );
  nor02 U3514 ( .Y(n6631), .A0(n6627), .A1(n6628) );
  inv01 U3515 ( .Y(n6630), .A(n6631) );
  inv02 U3516 ( .Y(member1796_0__11_), .A(n6632) );
  nor02 U3517 ( .Y(n6633), .A0(n6958), .A1(n7233) );
  nor02 U3518 ( .Y(n6634), .A0(n6965), .A1(n7378) );
  inv01 U3519 ( .Y(n6635), .A(n7532) );
  nor02 U3520 ( .Y(n6632), .A0(n6635), .A1(n6636) );
  nor02 U3521 ( .Y(n6637), .A0(n6633), .A1(n6634) );
  inv01 U3522 ( .Y(n6636), .A(n6637) );
  inv02 U3523 ( .Y(member1796_0__3_), .A(n6638) );
  nor02 U3524 ( .Y(n6639), .A0(n6958), .A1(n7225) );
  nor02 U3525 ( .Y(n6640), .A0(n6965), .A1(n7370) );
  inv01 U3526 ( .Y(n6641), .A(n7521) );
  nor02 U3527 ( .Y(n6638), .A0(n6641), .A1(n6642) );
  nor02 U3528 ( .Y(n6643), .A0(n6639), .A1(n6640) );
  inv01 U3529 ( .Y(n6642), .A(n6643) );
  inv02 U3530 ( .Y(member1796_0__21_), .A(n6644) );
  nor02 U3531 ( .Y(n6645), .A0(n6962), .A1(n7252) );
  nor02 U3532 ( .Y(n6646), .A0(n6967), .A1(n7388) );
  inv01 U3533 ( .Y(n6647), .A(n7525) );
  nor02 U3534 ( .Y(n6644), .A0(n6647), .A1(n6648) );
  nor02 U3535 ( .Y(n6649), .A0(n6645), .A1(n6646) );
  inv01 U3536 ( .Y(n6648), .A(n6649) );
  inv02 U3537 ( .Y(member2010_2__2_), .A(n6650) );
  nor02 U3538 ( .Y(n6651), .A0(n6962), .A1(n7296) );
  nor02 U3539 ( .Y(n6652), .A0(n6967), .A1(n7417) );
  inv01 U3540 ( .Y(n6653), .A(n5128) );
  nor02 U3541 ( .Y(n6650), .A0(n6653), .A1(n6654) );
  nor02 U3542 ( .Y(n6655), .A0(n6651), .A1(n6652) );
  inv01 U3543 ( .Y(n6654), .A(n6655) );
  inv02 U3544 ( .Y(member2010_2__19_), .A(n6656) );
  nor02 U3545 ( .Y(n6657), .A0(n6962), .A1(n7325) );
  nor02 U3546 ( .Y(n6658), .A0(n6967), .A1(n7434) );
  inv01 U3547 ( .Y(n6659), .A(n7493) );
  nor02 U3548 ( .Y(n6656), .A0(n6659), .A1(n6660) );
  nor02 U3549 ( .Y(n6661), .A0(n6657), .A1(n6658) );
  inv01 U3550 ( .Y(n6660), .A(n6661) );
  inv02 U3551 ( .Y(member1796_0__15_), .A(n6662) );
  nor02 U3552 ( .Y(n6663), .A0(n6960), .A1(n7240) );
  nor02 U3553 ( .Y(n6664), .A0(n6966), .A1(n7382) );
  inv01 U3554 ( .Y(n6665), .A(n7528) );
  nor02 U3555 ( .Y(n6662), .A0(n6665), .A1(n6666) );
  nor02 U3556 ( .Y(n6667), .A0(n6663), .A1(n6664) );
  inv01 U3557 ( .Y(n6666), .A(n6667) );
  inv02 U3558 ( .Y(member2010_2__20_), .A(n6668) );
  nor02 U3559 ( .Y(n6669), .A0(n6960), .A1(n7326) );
  nor02 U3560 ( .Y(n6670), .A0(n6966), .A1(n7435) );
  inv01 U3561 ( .Y(n6671), .A(n7491) );
  nor02 U3562 ( .Y(n6668), .A0(n6671), .A1(n6672) );
  nor02 U3563 ( .Y(n6673), .A0(n6669), .A1(n6670) );
  inv01 U3564 ( .Y(n6672), .A(n6673) );
  inv02 U3565 ( .Y(member1796_0__7_), .A(n6674) );
  nor02 U3566 ( .Y(n6675), .A0(n6960), .A1(n7229) );
  nor02 U3567 ( .Y(n6676), .A0(n6966), .A1(n7374) );
  inv01 U3568 ( .Y(n6677), .A(n7517) );
  nor02 U3569 ( .Y(n6674), .A0(n6677), .A1(n6678) );
  nor02 U3570 ( .Y(n6679), .A0(n6675), .A1(n6676) );
  inv01 U3571 ( .Y(n6678), .A(n6679) );
  inv02 U3572 ( .Y(member2010_2__1_), .A(n6680) );
  nor02 U3573 ( .Y(n6681), .A0(n6958), .A1(n7295) );
  nor02 U3574 ( .Y(n6682), .A0(n6965), .A1(n7416) );
  inv01 U3575 ( .Y(n6683), .A(n7492) );
  nor02 U3576 ( .Y(n6680), .A0(n6683), .A1(n6684) );
  nor02 U3577 ( .Y(n6685), .A0(n6681), .A1(n6682) );
  inv01 U3578 ( .Y(n6684), .A(n6685) );
  inv02 U3579 ( .Y(member2010_2__9_), .A(n6686) );
  nor02 U3580 ( .Y(n6687), .A0(n6958), .A1(n7306) );
  nor02 U3581 ( .Y(n6688), .A0(n6965), .A1(n7424) );
  inv01 U3582 ( .Y(n6689), .A(n7484) );
  nor02 U3583 ( .Y(n6686), .A0(n6689), .A1(n6690) );
  nor02 U3584 ( .Y(n6691), .A0(n6687), .A1(n6688) );
  inv01 U3585 ( .Y(n6690), .A(n6691) );
  inv02 U3586 ( .Y(member1796_0__1_), .A(n6692) );
  nor02 U3587 ( .Y(n6693), .A0(n6958), .A1(n7223) );
  nor02 U3588 ( .Y(n6694), .A0(n6965), .A1(n7368) );
  inv01 U3589 ( .Y(n6695), .A(n5388) );
  nor02 U3590 ( .Y(n6692), .A0(n6695), .A1(n6696) );
  nor02 U3591 ( .Y(n6697), .A0(n6693), .A1(n6694) );
  inv01 U3592 ( .Y(n6696), .A(n6697) );
  inv02 U3593 ( .Y(member1796_0__10_), .A(n6698) );
  nor02 U3594 ( .Y(n6699), .A0(n6962), .A1(n7232) );
  nor02 U3595 ( .Y(n6700), .A0(n6967), .A1(n7377) );
  inv01 U3596 ( .Y(n6701), .A(n5494) );
  nor02 U3597 ( .Y(n6698), .A0(n6701), .A1(n6702) );
  nor02 U3598 ( .Y(n6703), .A0(n6699), .A1(n6700) );
  inv01 U3599 ( .Y(n6702), .A(n6703) );
  inv02 U3600 ( .Y(member1796_0__5_), .A(n6704) );
  nor02 U3601 ( .Y(n6705), .A0(n6962), .A1(n7227) );
  nor02 U3602 ( .Y(n6706), .A0(n6967), .A1(n7372) );
  inv01 U3603 ( .Y(n6707), .A(n7519) );
  nor02 U3604 ( .Y(n6704), .A0(n6707), .A1(n6708) );
  nor02 U3605 ( .Y(n6709), .A0(n6705), .A1(n6706) );
  inv01 U3606 ( .Y(n6708), .A(n6709) );
  inv02 U3607 ( .Y(member2010_2__21_), .A(n6710) );
  nor02 U3608 ( .Y(n6711), .A0(n6962), .A1(n7327) );
  nor02 U3609 ( .Y(n6712), .A0(n6967), .A1(n7436) );
  inv01 U3610 ( .Y(n6713), .A(n7490) );
  nor02 U3611 ( .Y(n6710), .A0(n6713), .A1(n6714) );
  nor02 U3612 ( .Y(n6715), .A0(n6711), .A1(n6712) );
  inv01 U3613 ( .Y(n6714), .A(n6715) );
  inv02 U3614 ( .Y(member2010_2__7_), .A(n6716) );
  nor02 U3615 ( .Y(n6717), .A0(n6960), .A1(n7302) );
  nor02 U3616 ( .Y(n6718), .A0(n6966), .A1(n7422) );
  inv01 U3617 ( .Y(n6719), .A(n5166) );
  nor02 U3618 ( .Y(n6716), .A0(n6719), .A1(n6720) );
  nor02 U3619 ( .Y(n6721), .A0(n6717), .A1(n6718) );
  inv01 U3620 ( .Y(n6720), .A(n6721) );
  inv02 U3621 ( .Y(member2010_2__15_), .A(n6722) );
  nor02 U3622 ( .Y(n6723), .A0(n6960), .A1(n7318) );
  nor02 U3623 ( .Y(n6724), .A0(n6966), .A1(n7430) );
  inv01 U3624 ( .Y(n6725), .A(n7494) );
  nor02 U3625 ( .Y(n6722), .A0(n6725), .A1(n6726) );
  nor02 U3626 ( .Y(n6727), .A0(n6723), .A1(n6724) );
  inv01 U3627 ( .Y(n6726), .A(n6727) );
  inv02 U3628 ( .Y(member2010_2__3_), .A(n6728) );
  nor02 U3629 ( .Y(n6729), .A0(n6958), .A1(n7297) );
  nor02 U3630 ( .Y(n6730), .A0(n6965), .A1(n7418) );
  inv01 U3631 ( .Y(n6731), .A(n7487) );
  nor02 U3632 ( .Y(n6728), .A0(n6731), .A1(n6732) );
  nor02 U3633 ( .Y(n6733), .A0(n6729), .A1(n6730) );
  inv01 U3634 ( .Y(n6732), .A(n6733) );
  inv02 U3635 ( .Y(member2010_2__14_), .A(n6734) );
  nor02 U3636 ( .Y(n6735), .A0(n6958), .A1(n7316) );
  nor02 U3637 ( .Y(n6736), .A0(n6965), .A1(n7429) );
  inv01 U3638 ( .Y(n6737), .A(n7495) );
  nor02 U3639 ( .Y(n6734), .A0(n6737), .A1(n6738) );
  nor02 U3640 ( .Y(n6739), .A0(n6735), .A1(n6736) );
  inv01 U3641 ( .Y(n6738), .A(n6739) );
  inv02 U3642 ( .Y(member1796_0__22_), .A(n6740) );
  nor02 U3643 ( .Y(n6741), .A0(n6958), .A1(n7254) );
  nor02 U3644 ( .Y(n6742), .A0(n6965), .A1(n7389) );
  inv01 U3645 ( .Y(n6743), .A(n7524) );
  nor02 U3646 ( .Y(n6740), .A0(n6743), .A1(n6744) );
  nor02 U3647 ( .Y(n6745), .A0(n6741), .A1(n6742) );
  inv01 U3648 ( .Y(n6744), .A(n6745) );
  inv02 U3649 ( .Y(member1796_0__13_), .A(n6746) );
  nor02 U3650 ( .Y(n6747), .A0(n6962), .A1(n7236) );
  nor02 U3651 ( .Y(n6748), .A0(n6967), .A1(n7380) );
  inv01 U3652 ( .Y(n6749), .A(n7530) );
  nor02 U3653 ( .Y(n6746), .A0(n6749), .A1(n6750) );
  nor02 U3654 ( .Y(n6751), .A0(n6747), .A1(n6748) );
  inv01 U3655 ( .Y(n6750), .A(n6751) );
  inv02 U3656 ( .Y(member2010_2__16_), .A(n6752) );
  nor02 U3657 ( .Y(n6753), .A0(n6962), .A1(n7320) );
  nor02 U3658 ( .Y(n6754), .A0(n6967), .A1(n7431) );
  inv01 U3659 ( .Y(n6755), .A(n4872) );
  nor02 U3660 ( .Y(n6752), .A0(n6755), .A1(n6756) );
  nor02 U3661 ( .Y(n6757), .A0(n6753), .A1(n6754) );
  inv01 U3662 ( .Y(n6756), .A(n6757) );
  inv02 U3663 ( .Y(member2010_2__13_), .A(n6758) );
  nor02 U3664 ( .Y(n6759), .A0(n6962), .A1(n7314) );
  nor02 U3665 ( .Y(n6760), .A0(n6967), .A1(n7428) );
  inv01 U3666 ( .Y(n6761), .A(n7496) );
  nor02 U3667 ( .Y(n6758), .A0(n6761), .A1(n6762) );
  nor02 U3668 ( .Y(n6763), .A0(n6759), .A1(n6760) );
  inv01 U3669 ( .Y(n6762), .A(n6763) );
  inv02 U3670 ( .Y(member1796_0__20_), .A(n6764) );
  nor02 U3671 ( .Y(n6765), .A0(n6960), .A1(n7250) );
  nor02 U3672 ( .Y(n6766), .A0(n6966), .A1(n7387) );
  inv01 U3673 ( .Y(n6767), .A(n7526) );
  nor02 U3674 ( .Y(n6764), .A0(n6767), .A1(n6768) );
  nor02 U3675 ( .Y(n6769), .A0(n6765), .A1(n6766) );
  inv01 U3676 ( .Y(n6768), .A(n6769) );
  inv02 U3677 ( .Y(member1796_0__18_), .A(n6770) );
  nor02 U3678 ( .Y(n6771), .A0(n6960), .A1(n7246) );
  nor02 U3679 ( .Y(n6772), .A0(n6966), .A1(n7385) );
  inv01 U3680 ( .Y(n6773), .A(n5586) );
  nor02 U3681 ( .Y(n6770), .A0(n6773), .A1(n6774) );
  nor02 U3682 ( .Y(n6775), .A0(n6771), .A1(n6772) );
  inv01 U3683 ( .Y(n6774), .A(n6775) );
  inv02 U3684 ( .Y(member1796_0__12_), .A(n6776) );
  nor02 U3685 ( .Y(n6777), .A0(n6960), .A1(n7234) );
  nor02 U3686 ( .Y(n6778), .A0(n6966), .A1(n7379) );
  inv01 U3687 ( .Y(n6779), .A(n7531) );
  nor02 U3688 ( .Y(n6776), .A0(n6779), .A1(n6780) );
  nor02 U3689 ( .Y(n6781), .A0(n6777), .A1(n6778) );
  inv01 U3690 ( .Y(n6780), .A(n6781) );
  inv02 U3691 ( .Y(member1796_0__4_), .A(n6782) );
  nor02 U3692 ( .Y(n6783), .A0(n6960), .A1(n7226) );
  nor02 U3693 ( .Y(n6784), .A0(n6966), .A1(n7371) );
  inv01 U3694 ( .Y(n6785), .A(n7520) );
  nor02 U3695 ( .Y(n6782), .A0(n6785), .A1(n6786) );
  nor02 U3696 ( .Y(n6787), .A0(n6783), .A1(n6784) );
  inv01 U3697 ( .Y(n6786), .A(n6787) );
  inv02 U3698 ( .Y(member2010_2__18_), .A(n6788) );
  nor02 U3699 ( .Y(n6789), .A0(n6960), .A1(n7324) );
  nor02 U3700 ( .Y(n6790), .A0(n6966), .A1(n7433) );
  inv01 U3701 ( .Y(n6791), .A(n4912) );
  nor02 U3702 ( .Y(n6788), .A0(n6791), .A1(n6792) );
  nor02 U3703 ( .Y(n6793), .A0(n6789), .A1(n6790) );
  inv01 U3704 ( .Y(n6792), .A(n6793) );
  inv02 U3705 ( .Y(member2010_2__10_), .A(n6794) );
  nor02 U3706 ( .Y(n6795), .A0(n6962), .A1(n7308) );
  nor02 U3707 ( .Y(n6796), .A0(n6967), .A1(n7425) );
  inv01 U3708 ( .Y(n6797), .A(n7499) );
  nor02 U3709 ( .Y(n6794), .A0(n6797), .A1(n6798) );
  nor02 U3710 ( .Y(n6799), .A0(n6795), .A1(n6796) );
  inv01 U3711 ( .Y(n6798), .A(n6799) );
  inv02 U3712 ( .Y(member2010_2__8_), .A(n6800) );
  nor02 U3713 ( .Y(n6801), .A0(n6962), .A1(n7304) );
  nor02 U3714 ( .Y(n6802), .A0(n6967), .A1(n7423) );
  inv01 U3715 ( .Y(n6803), .A(n7485) );
  nor02 U3716 ( .Y(n6800), .A0(n6803), .A1(n6804) );
  nor02 U3717 ( .Y(n6805), .A0(n6801), .A1(n6802) );
  inv01 U3718 ( .Y(n6804), .A(n6805) );
  inv02 U3719 ( .Y(member1796_0__8_), .A(n6806) );
  nor02 U3720 ( .Y(n6807), .A0(n6962), .A1(n7230) );
  nor02 U3721 ( .Y(n6808), .A0(n6967), .A1(n7375) );
  inv01 U3722 ( .Y(n6809), .A(n7516) );
  nor02 U3723 ( .Y(n6806), .A0(n6809), .A1(n6810) );
  nor02 U3724 ( .Y(n6811), .A0(n6807), .A1(n6808) );
  inv01 U3725 ( .Y(n6810), .A(n6811) );
  inv02 U3726 ( .Y(member2010_2__22_), .A(n6812) );
  nor02 U3727 ( .Y(n6813), .A0(n6958), .A1(n7328) );
  nor02 U3728 ( .Y(n6814), .A0(n6965), .A1(n7437) );
  inv01 U3729 ( .Y(n6815), .A(n7489) );
  nor02 U3730 ( .Y(n6812), .A0(n6815), .A1(n6816) );
  nor02 U3731 ( .Y(n6817), .A0(n6813), .A1(n6814) );
  inv01 U3732 ( .Y(n6816), .A(n6817) );
  inv02 U3733 ( .Y(member1796_0__14_), .A(n6818) );
  nor02 U3734 ( .Y(n6819), .A0(n6958), .A1(n7238) );
  nor02 U3735 ( .Y(n6820), .A0(n6965), .A1(n7381) );
  inv01 U3736 ( .Y(n6821), .A(n7529) );
  nor02 U3737 ( .Y(n6818), .A0(n6821), .A1(n6822) );
  nor02 U3738 ( .Y(n6823), .A0(n6819), .A1(n6820) );
  inv01 U3739 ( .Y(n6822), .A(n6823) );
  inv02 U3740 ( .Y(member1796_0__2_), .A(n6824) );
  nor02 U3741 ( .Y(n6825), .A0(n6962), .A1(n7224) );
  nor02 U3742 ( .Y(n6826), .A0(n6967), .A1(n7369) );
  inv01 U3743 ( .Y(n6827), .A(n7522) );
  nor02 U3744 ( .Y(n6824), .A0(n6827), .A1(n6828) );
  nor02 U3745 ( .Y(n6829), .A0(n6825), .A1(n6826) );
  inv01 U3746 ( .Y(n6828), .A(n6829) );
  inv02 U3747 ( .Y(member1796_0__19_), .A(n6830) );
  nor02 U3748 ( .Y(n6831), .A0(n6962), .A1(n7248) );
  nor02 U3749 ( .Y(n6832), .A0(n6967), .A1(n7386) );
  inv01 U3750 ( .Y(n6833), .A(n7527) );
  nor02 U3751 ( .Y(n6830), .A0(n6833), .A1(n6834) );
  nor02 U3752 ( .Y(n6835), .A0(n6831), .A1(n6832) );
  inv01 U3753 ( .Y(n6834), .A(n6835) );
  inv02 U3754 ( .Y(member2010_2__5_), .A(n6836) );
  nor02 U3755 ( .Y(n6837), .A0(n6962), .A1(n7299) );
  nor02 U3756 ( .Y(n6838), .A0(n6967), .A1(n7420) );
  inv01 U3757 ( .Y(n6839), .A(n5548) );
  nor02 U3758 ( .Y(n6836), .A0(n6839), .A1(n6840) );
  nor02 U3759 ( .Y(n6841), .A0(n6837), .A1(n6838) );
  inv01 U3760 ( .Y(n6840), .A(n6841) );
  inv02 U3761 ( .Y(member2010_2__17_), .A(n6842) );
  nor02 U3762 ( .Y(n6843), .A0(n6958), .A1(n7322) );
  nor02 U3763 ( .Y(n6844), .A0(n6965), .A1(n7432) );
  inv01 U3764 ( .Y(n6845), .A(n5348) );
  nor02 U3765 ( .Y(n6842), .A0(n6845), .A1(n6846) );
  nor02 U3766 ( .Y(n6847), .A0(n6843), .A1(n6844) );
  inv01 U3767 ( .Y(n6846), .A(n6847) );
  inv02 U3768 ( .Y(member1796_0__9_), .A(n6848) );
  nor02 U3769 ( .Y(n6849), .A0(n6958), .A1(n7231) );
  nor02 U3770 ( .Y(n6850), .A0(n6965), .A1(n7376) );
  inv01 U3771 ( .Y(n6851), .A(n5588) );
  nor02 U3772 ( .Y(n6848), .A0(n6851), .A1(n6852) );
  nor02 U3773 ( .Y(n6853), .A0(n6849), .A1(n6850) );
  inv01 U3774 ( .Y(n6852), .A(n6853) );
  inv02 U3775 ( .Y(member1796_0__17_), .A(n6854) );
  nor02 U3776 ( .Y(n6855), .A0(n6958), .A1(n7244) );
  nor02 U3777 ( .Y(n6856), .A0(n6965), .A1(n7384) );
  inv01 U3778 ( .Y(n6857), .A(n5244) );
  nor02 U3779 ( .Y(n6854), .A0(n6857), .A1(n6858) );
  nor02 U3780 ( .Y(n6859), .A0(n6855), .A1(n6856) );
  inv01 U3781 ( .Y(n6858), .A(n6859) );
  inv02 U3782 ( .Y(member1883_1__0_), .A(n6860) );
  nor02 U3783 ( .Y(n6861), .A0(n6960), .A1(n7258) );
  nor02 U3784 ( .Y(n6862), .A0(n6966), .A1(n7391) );
  inv01 U3785 ( .Y(n6863), .A(n7515) );
  nor02 U3786 ( .Y(n6860), .A0(n6863), .A1(n6864) );
  nor02 U3787 ( .Y(n6865), .A0(n6861), .A1(n6862) );
  inv01 U3788 ( .Y(n6864), .A(n6865) );
  inv02 U3789 ( .Y(member2010_2__0_), .A(n6866) );
  nor02 U3790 ( .Y(n6867), .A0(n6960), .A1(n7294) );
  nor02 U3791 ( .Y(n6868), .A0(n6966), .A1(n7415) );
  inv01 U3792 ( .Y(n6869), .A(n7500) );
  nor02 U3793 ( .Y(n6866), .A0(n6869), .A1(n6870) );
  nor02 U3794 ( .Y(n6871), .A0(n6867), .A1(n6868) );
  inv01 U3795 ( .Y(n6870), .A(n6871) );
  inv02 U3796 ( .Y(member1796_0__0_), .A(n6872) );
  nor02 U3797 ( .Y(n6873), .A0(n6960), .A1(n7222) );
  nor02 U3798 ( .Y(n6874), .A0(n6966), .A1(n7367) );
  inv01 U3799 ( .Y(n6875), .A(n7533) );
  nor02 U3800 ( .Y(n6872), .A0(n6875), .A1(n6876) );
  nor02 U3801 ( .Y(n6877), .A0(n6873), .A1(n6874) );
  inv01 U3802 ( .Y(n6876), .A(n6877) );
  inv02 U3803 ( .Y(member2137_3__0_), .A(n6878) );
  nor02 U3804 ( .Y(n6879), .A0(n6960), .A1(n7330) );
  nor02 U3805 ( .Y(n6880), .A0(n6966), .A1(n7439) );
  inv01 U3806 ( .Y(n6881), .A(n7483) );
  nor02 U3807 ( .Y(n6878), .A0(n6881), .A1(n6882) );
  nor02 U3808 ( .Y(n6883), .A0(n6879), .A1(n6880) );
  inv01 U3809 ( .Y(n6882), .A(n6883) );
  inv02 U3810 ( .Y(n7124), .A(n6884) );
  inv01 U3811 ( .Y(n6885), .A(n7221) );
  inv01 U3812 ( .Y(n6886), .A(n6936) );
  inv01 U3813 ( .Y(n6887), .A(n6942) );
  nand02 U3814 ( .Y(n6884), .A0(n6887), .A1(n6888) );
  nand02 U3815 ( .Y(n6889), .A0(n6885), .A1(n6886) );
  inv01 U3816 ( .Y(n6888), .A(n6889) );
  buf04 U3817 ( .Y(n6942), .A(count_1_) );
  inv04 U3818 ( .Y(n6936), .A(n6935) );
  buf02 U3819 ( .Y(n6890), .A(n6996) );
  buf02 U3820 ( .Y(n6892), .A(n6996) );
  buf02 U3821 ( .Y(n6891), .A(n6996) );
  buf02 U3822 ( .Y(n6893), .A(member996_4__4_) );
  buf02 U3823 ( .Y(n6894), .A(member996_4__2_) );
  buf02 U3824 ( .Y(n6895), .A(member360_1__1_) );
  buf02 U3825 ( .Y(n6896), .A(member360_1__3_) );
  buf02 U3826 ( .Y(n6897), .A(member638_2__3_) );
  buf02 U3827 ( .Y(n6898), .A(member996_4__1_) );
  ao22 U3828 ( .Y(n6899), .A0(n3540), .A1(n6943), .B0(n3552), .B1(n7221) );
  inv02 U3829 ( .Y(n6900), .A(n6899) );
  ao22 U3830 ( .Y(n6901), .A0(n3537), .A1(n6943), .B0(n3549), .B1(n7221) );
  inv02 U3831 ( .Y(n6902), .A(n6901) );
  ao22 U3832 ( .Y(n6903), .A0(n3544), .A1(n6943), .B0(n3556), .B1(n7221) );
  inv02 U3833 ( .Y(n6904), .A(n6903) );
  ao22 U3834 ( .Y(n6905), .A0(n3542), .A1(n6943), .B0(n3554), .B1(n7221) );
  inv02 U3835 ( .Y(n6906), .A(n6905) );
  ao22 U3836 ( .Y(n6907), .A0(n3547), .A1(n6945), .B0(n3559), .B1(n7221) );
  inv02 U3837 ( .Y(n6908), .A(n6907) );
  ao22 U3838 ( .Y(n6909), .A0(n3565), .A1(n6941), .B0(n3577), .B1(n7366) );
  inv02 U3839 ( .Y(n6910), .A(n6909) );
  ao22 U3840 ( .Y(n6911), .A0(n3567), .A1(n6941), .B0(n3579), .B1(n7366) );
  inv02 U3841 ( .Y(n6912), .A(n6911) );
  ao22 U3842 ( .Y(n6913), .A0(n3538), .A1(n6943), .B0(n3550), .B1(n7221) );
  inv02 U3843 ( .Y(n6914), .A(n6913) );
  ao22 U3844 ( .Y(n6915), .A0(n3536), .A1(n6945), .B0(n3548), .B1(n7221) );
  inv02 U3845 ( .Y(n6916), .A(n6915) );
  ao22 U3846 ( .Y(n6917), .A0(n3546), .A1(n6945), .B0(n3558), .B1(n7221) );
  inv02 U3847 ( .Y(n6918), .A(n6917) );
  ao22 U3848 ( .Y(n6919), .A0(n3541), .A1(n6945), .B0(n3553), .B1(n7221) );
  inv02 U3849 ( .Y(n6920), .A(n6919) );
  ao22 U3850 ( .Y(n6921), .A0(n3539), .A1(n6945), .B0(n3551), .B1(n7221) );
  inv02 U3851 ( .Y(n6922), .A(n6921) );
  ao22 U3852 ( .Y(n6923), .A0(n3560), .A1(n6942), .B0(n3572), .B1(n7366) );
  inv02 U3853 ( .Y(n6924), .A(n6923) );
  ao22 U3854 ( .Y(n6925), .A0(n3570), .A1(n6942), .B0(n3582), .B1(n7366) );
  inv02 U3855 ( .Y(n6926), .A(n6925) );
  ao22 U3856 ( .Y(n6927), .A0(n3568), .A1(n6942), .B0(n3580), .B1(n7366) );
  inv02 U3857 ( .Y(n6928), .A(n6927) );
  ao22 U3858 ( .Y(n6929), .A0(n3566), .A1(n6942), .B0(n3578), .B1(n7366) );
  inv02 U3859 ( .Y(n6930), .A(n6929) );
  ao22 U3860 ( .Y(n6931), .A0(n3571), .A1(n6942), .B0(n3583), .B1(n7366) );
  inv02 U3861 ( .Y(n6932), .A(n6931) );
  ao22 U3862 ( .Y(n6933), .A0(n3563), .A1(n6942), .B0(n3575), .B1(n7366) );
  inv02 U3863 ( .Y(n6934), .A(n6933) );
  inv02 U3864 ( .Y(n7012), .A(n____return2214_14_) );
  inv02 U3865 ( .Y(n7017), .A(n____return2214_19_) );
  inv02 U3866 ( .Y(n7015), .A(n____return2214_17_) );
  inv02 U3867 ( .Y(n7013), .A(n____return2214_15_) );
  inv02 U3868 ( .Y(n7002), .A(n____return2214_4_) );
  inv02 U3869 ( .Y(n7018), .A(n____return2214_20_) );
  inv02 U3870 ( .Y(n7003), .A(n____return2214_5_) );
  inv02 U3871 ( .Y(n7005), .A(n____return2214_7_) );
  inv02 U3872 ( .Y(n7011), .A(n____return2214_13_) );
  inv02 U3873 ( .Y(n7020), .A(n____return2214_22_) );
  inv02 U3874 ( .Y(n6999), .A(n____return2214_1_) );
  inv02 U3875 ( .Y(n7016), .A(n____return2214_18_) );
  inv02 U3876 ( .Y(n7009), .A(n____return2214_11_) );
  inv02 U3877 ( .Y(n7006), .A(n____return2214_8_) );
  inv02 U3878 ( .Y(n7004), .A(n____return2214_6_) );
  inv02 U3879 ( .Y(n7010), .A(n____return2214_12_) );
  inv02 U3880 ( .Y(n7021), .A(n____return2214_23_) );
  inv02 U3881 ( .Y(n7014), .A(n____return2214_16_) );
  inv02 U3882 ( .Y(n7019), .A(n____return2214_21_) );
  inv02 U3883 ( .Y(n7001), .A(n____return2214_3_) );
  inv02 U3884 ( .Y(n7000), .A(n____return2214_2_) );
  inv02 U3885 ( .Y(n7007), .A(n____return2214_9_) );
  inv08 U3886 ( .Y(n6995), .A(s_state) );
  inv02 U3887 ( .Y(n7008), .A(n____return2214_10_) );
  inv08 U3888 ( .Y(n6935), .A(count_2_) );
  aoi22 U3889 ( .Y(n6937), .A0(n7366), .A1(n6946), .B0(n6940), .B1(n7221) );
  buf02 U3890 ( .Y(n6938), .A(n7534) );
  buf02 U3891 ( .Y(n6939), .A(n6937) );
  buf08 U3892 ( .Y(n6941), .A(count_1_) );
  buf16 U3893 ( .Y(n6946), .A(count_0_) );
  buf08 U3894 ( .Y(n6945), .A(count_0_) );
  buf08 U3895 ( .Y(n6947), .A(n6976) );
  inv12 U3896 ( .Y(n6948), .A(n6947) );
  inv12 U3897 ( .Y(n6950), .A(n6947) );
  inv12 U3898 ( .Y(n6949), .A(n6947) );
  buf16 U3899 ( .Y(n6951), .A(n7023) );
  buf16 U3900 ( .Y(n6952), .A(n6279) );
  buf16 U3901 ( .Y(n6953), .A(n6998) );
  buf16 U3902 ( .Y(n6954), .A(n6281) );
  nand02 U3903 ( .Y(n6955), .A0(n6938), .A1(n6945) );
  nand02 U3904 ( .Y(n6956), .A0(n6939), .A1(n6943) );
  inv16 U3905 ( .Y(n6958), .A(n6957) );
  inv04 U3906 ( .Y(n6959), .A(n6955) );
  inv16 U3907 ( .Y(n6960), .A(n6959) );
  inv04 U3908 ( .Y(n6961), .A(n6956) );
  inv16 U3909 ( .Y(n6962), .A(n6961) );
  nand02 U3910 ( .Y(n6963), .A0(n6938), .A1(n7221) );
  nand02 U3911 ( .Y(n6964), .A0(n6938), .A1(n7221) );
  buf16 U3912 ( .Y(n6965), .A(n7026) );
  buf16 U3913 ( .Y(n6966), .A(n6963) );
  buf16 U3914 ( .Y(n6967), .A(n6964) );
  nor02 U3915 ( .Y(n6968), .A0(n7221), .A1(n6939) );
  nor02 U3916 ( .Y(n6969), .A0(n7221), .A1(n6938) );
  buf12 U3917 ( .Y(n6970), .A(n7022) );
  buf12 U3918 ( .Y(n6971), .A(n6968) );
  buf12 U3919 ( .Y(n6972), .A(n6969) );
  inv08 U3920 ( .Y(n6973), .A(n6307) );
  inv16 U3921 ( .Y(n6974), .A(n6973) );
  inv16 U3922 ( .Y(n6975), .A(n6973) );
  inv01 U3923 ( .Y(n6977), .A(n7221) );
  inv01 U3924 ( .Y(n6978), .A(n6936) );
  inv01 U3925 ( .Y(n6979), .A(n7366) );
  nand02 U3926 ( .Y(n6976), .A0(n6979), .A1(n6980) );
  nand02 U3927 ( .Y(n6981), .A0(n6977), .A1(n6978) );
  inv01 U3928 ( .Y(n6980), .A(n6981) );
  buf16 U3929 ( .Y(n6982), .A(n7027) );
  buf16 U3930 ( .Y(n6983), .A(n6287) );
  buf16 U3931 ( .Y(n6984), .A(n6983) );
  buf16 U3932 ( .Y(n6986), .A(n6988) );
  buf16 U3933 ( .Y(n6987), .A(n6985) );
  buf16 U3934 ( .Y(n6988), .A(n6295) );
  inv08 U3935 ( .Y(n6989), .A(n7124) );
  inv08 U3936 ( .Y(n7366), .A(n6941) );
  inv08 U3937 ( .Y(n7221), .A(n6944) );
  ao21 U3961 ( .Y(n4770), .A0(n6303), .A1(n6993), .B0(n4772) );
  inv01 U3962 ( .Y(n6993), .A(n6892) );
  ao21 U3963 ( .Y(n4769), .A0(s_state), .A1(n6890), .B0(s_state83) );
  mux21 U3964 ( .Y(n4766), .A0(n4206), .A1(n7000), .S0(n6953) );
  mux21 U3965 ( .Y(n4765), .A0(n4207), .A1(n7001), .S0(n6953) );
  mux21 U3966 ( .Y(n4764), .A0(n4208), .A1(n7002), .S0(n6953) );
  mux21 U3967 ( .Y(n4763), .A0(n4209), .A1(n7003), .S0(n6953) );
  mux21 U3968 ( .Y(n4762), .A0(n4210), .A1(n7004), .S0(n6953) );
  mux21 U3969 ( .Y(n4761), .A0(n4211), .A1(n7005), .S0(n6953) );
  mux21 U3970 ( .Y(n4760), .A0(n4212), .A1(n7006), .S0(n6953) );
  mux21 U3971 ( .Y(n4759), .A0(n4213), .A1(n7007), .S0(n6953) );
  mux21 U3972 ( .Y(n4758), .A0(n4191), .A1(n7008), .S0(n6953) );
  mux21 U3973 ( .Y(n4757), .A0(n4192), .A1(n7009), .S0(n6953) );
  mux21 U3974 ( .Y(n4756), .A0(n4193), .A1(n7010), .S0(n6953) );
  mux21 U3975 ( .Y(n4755), .A0(n4194), .A1(n7011), .S0(n6953) );
  mux21 U3976 ( .Y(n4754), .A0(n4195), .A1(n7012), .S0(n6953) );
  mux21 U3977 ( .Y(n4753), .A0(n4196), .A1(n7013), .S0(n6953) );
  mux21 U3978 ( .Y(n4752), .A0(n4197), .A1(n7014), .S0(n6953) );
  mux21 U3979 ( .Y(n4751), .A0(n4198), .A1(n7015), .S0(n6953) );
  mux21 U3980 ( .Y(n4750), .A0(n4199), .A1(n7016), .S0(n6953) );
  mux21 U3981 ( .Y(n4749), .A0(n4200), .A1(n7017), .S0(n6953) );
  mux21 U3982 ( .Y(n4748), .A0(n4202), .A1(n7018), .S0(n6953) );
  mux21 U3983 ( .Y(n4747), .A0(n4203), .A1(n7019), .S0(n6953) );
  and02 U3984 ( .Y(n6998), .A0(n6970), .A1(n6305) );
  mux21 U3985 ( .Y(n4743), .A0(n4225), .A1(n6999), .S0(n6951) );
  mux21 U3986 ( .Y(n4742), .A0(n4230), .A1(n7000), .S0(n6951) );
  mux21 U3987 ( .Y(n4741), .A0(n4231), .A1(n7001), .S0(n6951) );
  mux21 U3988 ( .Y(n4740), .A0(n4232), .A1(n7002), .S0(n6951) );
  mux21 U3989 ( .Y(n4739), .A0(n4233), .A1(n7003), .S0(n6951) );
  mux21 U3990 ( .Y(n4738), .A0(n4234), .A1(n7004), .S0(n6951) );
  mux21 U3991 ( .Y(n4737), .A0(n4235), .A1(n7005), .S0(n6951) );
  mux21 U3992 ( .Y(n4736), .A0(n4236), .A1(n7006), .S0(n6951) );
  mux21 U3993 ( .Y(n4735), .A0(n4237), .A1(n7007), .S0(n6951) );
  mux21 U3994 ( .Y(n4734), .A0(n4215), .A1(n7008), .S0(n6951) );
  mux21 U3995 ( .Y(n4733), .A0(n4216), .A1(n7009), .S0(n6951) );
  mux21 U3996 ( .Y(n4732), .A0(n4217), .A1(n7010), .S0(n6951) );
  mux21 U3997 ( .Y(n4731), .A0(n4218), .A1(n7011), .S0(n6951) );
  mux21 U3998 ( .Y(n4730), .A0(n4219), .A1(n7012), .S0(n6951) );
  mux21 U3999 ( .Y(n4729), .A0(n4220), .A1(n7013), .S0(n6951) );
  mux21 U4000 ( .Y(n4728), .A0(n4221), .A1(n7014), .S0(n6951) );
  mux21 U4001 ( .Y(n4727), .A0(n4222), .A1(n7015), .S0(n6951) );
  mux21 U4002 ( .Y(n4726), .A0(n4223), .A1(n7016), .S0(n6951) );
  mux21 U4003 ( .Y(n4725), .A0(n4224), .A1(n7017), .S0(n6951) );
  mux21 U4004 ( .Y(n4724), .A0(n4226), .A1(n7018), .S0(n6951) );
  mux21 U4005 ( .Y(n4723), .A0(n4227), .A1(n7019), .S0(n6951) );
  mux21 U4006 ( .Y(n4722), .A0(n4228), .A1(n7020), .S0(n6951) );
  mux21 U4007 ( .Y(n4721), .A0(n4229), .A1(n7021), .S0(n6951) );
  and02 U4008 ( .Y(n7023), .A0(n6974), .A1(n6305) );
  mux21 U4009 ( .Y(n4720), .A0(n4238), .A1(n6997), .S0(n6952) );
  mux21 U4010 ( .Y(n4719), .A0(n4249), .A1(n6999), .S0(n6952) );
  mux21 U4011 ( .Y(n4718), .A0(n4254), .A1(n7000), .S0(n6952) );
  mux21 U4012 ( .Y(n4716), .A0(n4256), .A1(n7002), .S0(n6952) );
  mux21 U4013 ( .Y(n4715), .A0(n4257), .A1(n7003), .S0(n6952) );
  mux21 U4014 ( .Y(n4714), .A0(n4258), .A1(n7004), .S0(n6952) );
  mux21 U4015 ( .Y(n4713), .A0(n4259), .A1(n7005), .S0(n6952) );
  mux21 U4016 ( .Y(n4712), .A0(n4260), .A1(n7006), .S0(n6952) );
  mux21 U4017 ( .Y(n4711), .A0(n4261), .A1(n7007), .S0(n6952) );
  mux21 U4018 ( .Y(n4710), .A0(n4239), .A1(n7008), .S0(n6952) );
  mux21 U4019 ( .Y(n4709), .A0(n4240), .A1(n7009), .S0(n6952) );
  mux21 U4020 ( .Y(n4707), .A0(n4242), .A1(n7011), .S0(n6952) );
  mux21 U4021 ( .Y(n4706), .A0(n4243), .A1(n7012), .S0(n6952) );
  mux21 U4022 ( .Y(n4705), .A0(n4244), .A1(n7013), .S0(n6952) );
  mux21 U4023 ( .Y(n4704), .A0(n4245), .A1(n7014), .S0(n6952) );
  mux21 U4024 ( .Y(n4703), .A0(n4246), .A1(n7015), .S0(n6952) );
  mux21 U4025 ( .Y(n4702), .A0(n4247), .A1(n7016), .S0(n6952) );
  mux21 U4026 ( .Y(n4701), .A0(n4248), .A1(n7017), .S0(n6952) );
  mux21 U4027 ( .Y(n4700), .A0(n4250), .A1(n7018), .S0(n6952) );
  mux21 U4028 ( .Y(n4699), .A0(n4251), .A1(n7019), .S0(n6952) );
  mux21 U4029 ( .Y(n4698), .A0(n4252), .A1(n7020), .S0(n6952) );
  mux21 U4030 ( .Y(n4695), .A0(n4273), .A1(n6999), .S0(n6954) );
  mux21 U4031 ( .Y(n4694), .A0(n4278), .A1(n7000), .S0(n6954) );
  mux21 U4032 ( .Y(n4693), .A0(n4279), .A1(n7001), .S0(n6954) );
  mux21 U4033 ( .Y(n4692), .A0(n4280), .A1(n7002), .S0(n6954) );
  mux21 U4034 ( .Y(n4691), .A0(n4281), .A1(n7003), .S0(n6954) );
  mux21 U4035 ( .Y(n4690), .A0(n4282), .A1(n7004), .S0(n6954) );
  mux21 U4036 ( .Y(n4689), .A0(n4283), .A1(n7005), .S0(n6954) );
  mux21 U4037 ( .Y(n4688), .A0(n4284), .A1(n7006), .S0(n6954) );
  mux21 U4038 ( .Y(n4687), .A0(n4285), .A1(n7007), .S0(n6954) );
  mux21 U4039 ( .Y(n4686), .A0(n4263), .A1(n7008), .S0(n6954) );
  mux21 U4040 ( .Y(n4685), .A0(n4264), .A1(n7009), .S0(n6954) );
  mux21 U4041 ( .Y(n4684), .A0(n4265), .A1(n7010), .S0(n6954) );
  mux21 U4042 ( .Y(n4683), .A0(n4266), .A1(n7011), .S0(n6954) );
  mux21 U4043 ( .Y(n4682), .A0(n4267), .A1(n7012), .S0(n6954) );
  mux21 U4044 ( .Y(n4681), .A0(n4268), .A1(n7013), .S0(n6954) );
  mux21 U4045 ( .Y(n4680), .A0(n4269), .A1(n7014), .S0(n6954) );
  mux21 U4046 ( .Y(n4679), .A0(n4270), .A1(n7015), .S0(n6954) );
  mux21 U4047 ( .Y(n4678), .A0(n4271), .A1(n7016), .S0(n6954) );
  mux21 U4048 ( .Y(n4677), .A0(n4272), .A1(n7017), .S0(n6954) );
  mux21 U4049 ( .Y(n4676), .A0(n4274), .A1(n7018), .S0(n6954) );
  mux21 U4050 ( .Y(n4675), .A0(n4275), .A1(n7019), .S0(n6954) );
  mux21 U4051 ( .Y(n4673), .A0(n4277), .A1(n7021), .S0(n6954) );
  inv01 U4052 ( .Y(n7025), .A(n6305) );
  inv01 U4053 ( .Y(n7028), .A(larray[0]) );
  inv01 U4054 ( .Y(n7029), .A(larray[1]) );
  inv01 U4055 ( .Y(n7030), .A(larray[2]) );
  inv01 U4056 ( .Y(n7031), .A(larray[3]) );
  inv01 U4057 ( .Y(n7032), .A(larray[4]) );
  inv01 U4058 ( .Y(n7033), .A(larray[5]) );
  inv01 U4059 ( .Y(n7034), .A(larray[6]) );
  inv01 U4060 ( .Y(n7035), .A(larray[7]) );
  inv01 U4061 ( .Y(n7036), .A(larray[8]) );
  inv01 U4062 ( .Y(n7037), .A(larray[9]) );
  inv01 U4063 ( .Y(n7038), .A(larray[10]) );
  inv01 U4064 ( .Y(n7039), .A(larray[11]) );
  inv01 U4065 ( .Y(n4660), .A(n7040) );
  mux21 U4066 ( .Y(n7040), .A0(larray[12]), .A1(n____return437_0_), .S0(n6982)
         );
  inv01 U4067 ( .Y(n4659), .A(n7041) );
  mux21 U4068 ( .Y(n7041), .A0(larray[13]), .A1(n____return437_1_), .S0(n6984)
         );
  inv01 U4069 ( .Y(n4658), .A(n7042) );
  mux21 U4070 ( .Y(n7042), .A0(larray[14]), .A1(n____return437_2_), .S0(n6983)
         );
  inv01 U4071 ( .Y(n4657), .A(n7043) );
  mux21 U4072 ( .Y(n7043), .A0(larray[15]), .A1(n____return437_3_), .S0(n6982)
         );
  inv01 U4073 ( .Y(n4656), .A(n7044) );
  mux21 U4074 ( .Y(n7044), .A0(larray[16]), .A1(n____return437_4_), .S0(n6984)
         );
  inv01 U4075 ( .Y(n4655), .A(n7045) );
  mux21 U4076 ( .Y(n7045), .A0(larray[17]), .A1(n____return437_5_), .S0(n6983)
         );
  inv01 U4077 ( .Y(n4654), .A(n7046) );
  mux21 U4078 ( .Y(n7046), .A0(larray[18]), .A1(n____return437_6_), .S0(n6982)
         );
  inv01 U4079 ( .Y(n4653), .A(n7047) );
  mux21 U4080 ( .Y(n7047), .A0(larray[19]), .A1(n____return437_7_), .S0(n6984)
         );
  inv01 U4081 ( .Y(n4652), .A(n7048) );
  mux21 U4082 ( .Y(n7048), .A0(larray[20]), .A1(n____return437_8_), .S0(n6983)
         );
  inv01 U4083 ( .Y(n4651), .A(n7049) );
  mux21 U4084 ( .Y(n7049), .A0(larray[21]), .A1(n____return437_9_), .S0(n6982)
         );
  inv01 U4085 ( .Y(n4650), .A(n7050) );
  mux21 U4086 ( .Y(n7050), .A0(larray[22]), .A1(n____return437_10_), .S0(n6984) );
  inv01 U4087 ( .Y(n4649), .A(n7051) );
  mux21 U4088 ( .Y(n7051), .A0(larray[23]), .A1(n____return437_11_), .S0(n6983) );
  inv01 U4089 ( .Y(n7052), .A(larray[24]) );
  inv01 U4090 ( .Y(n7053), .A(larray[25]) );
  inv01 U4091 ( .Y(n7054), .A(larray[26]) );
  inv01 U4092 ( .Y(n7055), .A(larray[27]) );
  inv01 U4093 ( .Y(n7056), .A(larray[28]) );
  inv01 U4094 ( .Y(n7057), .A(larray[29]) );
  inv01 U4095 ( .Y(n4642), .A(n7058) );
  mux21 U4096 ( .Y(n7058), .A0(larray[30]), .A1(n____return792_0_), .S0(n6982)
         );
  inv01 U4097 ( .Y(n4641), .A(n7059) );
  mux21 U4098 ( .Y(n7059), .A0(larray[31]), .A1(n____return792_1_), .S0(n6984)
         );
  inv01 U4099 ( .Y(n4640), .A(n7060) );
  mux21 U4100 ( .Y(n7060), .A0(larray[32]), .A1(n____return792_2_), .S0(n6983)
         );
  inv01 U4101 ( .Y(n4639), .A(n7061) );
  mux21 U4102 ( .Y(n7061), .A0(larray[33]), .A1(n____return792_3_), .S0(n6982)
         );
  inv01 U4103 ( .Y(n4638), .A(n7062) );
  mux21 U4104 ( .Y(n7062), .A0(larray[34]), .A1(n____return792_4_), .S0(n6984)
         );
  inv01 U4105 ( .Y(n4637), .A(n7063) );
  mux21 U4106 ( .Y(n7063), .A0(larray[35]), .A1(n____return792_5_), .S0(n6983)
         );
  inv01 U4107 ( .Y(n4636), .A(n7064) );
  mux21 U4108 ( .Y(n7064), .A0(larray[36]), .A1(n____return792_6_), .S0(n6982)
         );
  inv01 U4109 ( .Y(n4635), .A(n7065) );
  mux21 U4110 ( .Y(n7065), .A0(larray[37]), .A1(n____return792_7_), .S0(n6984)
         );
  inv01 U4111 ( .Y(n4634), .A(n7066) );
  mux21 U4112 ( .Y(n7066), .A0(larray[38]), .A1(n____return792_8_), .S0(n6983)
         );
  inv01 U4113 ( .Y(n4633), .A(n7067) );
  mux21 U4114 ( .Y(n7067), .A0(larray[39]), .A1(n____return792_9_), .S0(n6982)
         );
  inv01 U4115 ( .Y(n4632), .A(n7068) );
  mux21 U4116 ( .Y(n7068), .A0(larray[40]), .A1(n____return792_10_), .S0(n6984) );
  inv01 U4117 ( .Y(n4631), .A(n7069) );
  mux21 U4118 ( .Y(n7069), .A0(larray[41]), .A1(n____return792_11_), .S0(n6983) );
  inv01 U4119 ( .Y(n7070), .A(larray[42]) );
  inv01 U4120 ( .Y(n7071), .A(larray[43]) );
  inv01 U4121 ( .Y(n7072), .A(larray[44]) );
  inv01 U4122 ( .Y(n7073), .A(larray[45]) );
  inv01 U4123 ( .Y(n7074), .A(larray[46]) );
  inv01 U4124 ( .Y(n7075), .A(larray[47]) );
  inv01 U4125 ( .Y(n7076), .A(larray[48]) );
  inv01 U4126 ( .Y(n7077), .A(larray[49]) );
  inv01 U4127 ( .Y(n7078), .A(larray[50]) );
  inv01 U4128 ( .Y(n7079), .A(larray[51]) );
  inv01 U4129 ( .Y(n7080), .A(larray[52]) );
  inv01 U4130 ( .Y(n7081), .A(larray[53]) );
  inv01 U4131 ( .Y(n4618), .A(n7082) );
  mux21 U4132 ( .Y(n7082), .A0(larray[54]), .A1(n____return1150_0_), .S0(n6982) );
  inv01 U4133 ( .Y(n4617), .A(n7083) );
  mux21 U4134 ( .Y(n7083), .A0(larray[55]), .A1(n____return1150_1_), .S0(n6984) );
  inv01 U4135 ( .Y(n4616), .A(n7084) );
  mux21 U4136 ( .Y(n7084), .A0(larray[56]), .A1(n____return1150_2_), .S0(n6983) );
  inv01 U4137 ( .Y(n4615), .A(n7085) );
  mux21 U4138 ( .Y(n7085), .A0(larray[57]), .A1(n____return1150_3_), .S0(n6982) );
  inv01 U4139 ( .Y(n4614), .A(n7086) );
  mux21 U4140 ( .Y(n7086), .A0(larray[58]), .A1(n____return1150_4_), .S0(n6984) );
  inv01 U4141 ( .Y(n4613), .A(n7087) );
  mux21 U4142 ( .Y(n7087), .A0(larray[59]), .A1(n____return1150_5_), .S0(n6983) );
  inv01 U4143 ( .Y(n4612), .A(n7088) );
  mux21 U4144 ( .Y(n7088), .A0(larray[60]), .A1(n____return1150_6_), .S0(n6982) );
  inv01 U4145 ( .Y(n4611), .A(n7089) );
  mux21 U4146 ( .Y(n7089), .A0(larray[61]), .A1(n____return1150_7_), .S0(n6984) );
  inv01 U4147 ( .Y(n4610), .A(n7090) );
  mux21 U4148 ( .Y(n7090), .A0(larray[62]), .A1(n____return1150_8_), .S0(n6983) );
  inv01 U4149 ( .Y(n4609), .A(n7091) );
  mux21 U4150 ( .Y(n7091), .A0(larray[63]), .A1(n____return1150_9_), .S0(n6982) );
  inv01 U4151 ( .Y(n4608), .A(n7092) );
  mux21 U4152 ( .Y(n7092), .A0(larray[64]), .A1(n____return1150_10_), .S0(
        n6984) );
  inv01 U4153 ( .Y(n4607), .A(n7093) );
  mux21 U4154 ( .Y(n7093), .A0(larray[65]), .A1(n____return1150_11_), .S0(
        n6983) );
  inv01 U4155 ( .Y(n7094), .A(larray[66]) );
  inv01 U4156 ( .Y(n7095), .A(larray[67]) );
  inv01 U4157 ( .Y(n7096), .A(larray[68]) );
  inv01 U4158 ( .Y(n7097), .A(larray[69]) );
  inv01 U4159 ( .Y(n7098), .A(larray[70]) );
  inv01 U4160 ( .Y(n7099), .A(larray[71]) );
  inv01 U4161 ( .Y(n4600), .A(n7100) );
  mux21 U4162 ( .Y(n7100), .A0(larray[72]), .A1(n____return1508_0_), .S0(n6982) );
  inv01 U4163 ( .Y(n4599), .A(n7101) );
  mux21 U4164 ( .Y(n7101), .A0(larray[73]), .A1(n____return1508_1_), .S0(n6984) );
  inv01 U4165 ( .Y(n4598), .A(n7102) );
  mux21 U4166 ( .Y(n7102), .A0(larray[74]), .A1(n____return1508_2_), .S0(n6983) );
  inv01 U4167 ( .Y(n4597), .A(n7103) );
  mux21 U4168 ( .Y(n7103), .A0(larray[75]), .A1(n____return1508_3_), .S0(n6982) );
  inv01 U4169 ( .Y(n4596), .A(n7104) );
  mux21 U4170 ( .Y(n7104), .A0(larray[76]), .A1(n____return1508_4_), .S0(n6984) );
  inv01 U4171 ( .Y(n4595), .A(n7105) );
  mux21 U4172 ( .Y(n7105), .A0(larray[77]), .A1(n____return1508_5_), .S0(n6983) );
  inv01 U4173 ( .Y(n4594), .A(n7106) );
  mux21 U4174 ( .Y(n7106), .A0(larray[78]), .A1(n____return1508_6_), .S0(n6982) );
  inv01 U4175 ( .Y(n4593), .A(n7107) );
  mux21 U4176 ( .Y(n7107), .A0(larray[79]), .A1(n____return1508_7_), .S0(n6984) );
  inv01 U4177 ( .Y(n4592), .A(n7108) );
  mux21 U4178 ( .Y(n7108), .A0(larray[80]), .A1(n____return1508_8_), .S0(n6983) );
  inv01 U4179 ( .Y(n4591), .A(n7109) );
  mux21 U4180 ( .Y(n7109), .A0(larray[81]), .A1(n____return1508_9_), .S0(n6982) );
  inv01 U4181 ( .Y(n4590), .A(n7110) );
  mux21 U4182 ( .Y(n7110), .A0(larray[82]), .A1(n____return1508_10_), .S0(
        n6984) );
  inv01 U4183 ( .Y(n4589), .A(n7111) );
  mux21 U4184 ( .Y(n7111), .A0(larray[83]), .A1(n____return1508_11_), .S0(
        n6983) );
  inv01 U4185 ( .Y(n7112), .A(larray[84]) );
  inv01 U4186 ( .Y(n7113), .A(larray[85]) );
  inv01 U4187 ( .Y(n7114), .A(larray[86]) );
  inv01 U4188 ( .Y(n7115), .A(larray[87]) );
  inv01 U4189 ( .Y(n7116), .A(larray[88]) );
  inv01 U4190 ( .Y(n7117), .A(larray[89]) );
  inv01 U4191 ( .Y(n7118), .A(larray[90]) );
  inv01 U4192 ( .Y(n7119), .A(larray[91]) );
  inv01 U4193 ( .Y(n7120), .A(larray[92]) );
  inv01 U4194 ( .Y(n7121), .A(larray[93]) );
  inv01 U4195 ( .Y(n7122), .A(larray[94]) );
  inv01 U4196 ( .Y(n7123), .A(larray[95]) );
  inv01 U4197 ( .Y(n7125), .A(larray[96]) );
  inv01 U4198 ( .Y(n7126), .A(larray[97]) );
  inv01 U4199 ( .Y(n7127), .A(larray[98]) );
  inv01 U4200 ( .Y(n7128), .A(larray[99]) );
  inv01 U4201 ( .Y(n7129), .A(larray[100]) );
  inv01 U4202 ( .Y(n7130), .A(larray[101]) );
  inv01 U4203 ( .Y(n7131), .A(larray[102]) );
  inv01 U4204 ( .Y(n7132), .A(larray[103]) );
  inv01 U4205 ( .Y(n7133), .A(larray[104]) );
  inv01 U4206 ( .Y(n7134), .A(larray[105]) );
  inv01 U4207 ( .Y(n7135), .A(larray[106]) );
  inv01 U4208 ( .Y(n7136), .A(larray[107]) );
  inv01 U4209 ( .Y(n4564), .A(n7137) );
  mux21 U4210 ( .Y(n7137), .A0(larray[108]), .A1(n____return437_0_), .S0(n6992) );
  inv01 U4211 ( .Y(n4563), .A(n7138) );
  mux21 U4212 ( .Y(n7138), .A0(larray[109]), .A1(n____return437_1_), .S0(n6990) );
  inv01 U4213 ( .Y(n4562), .A(n7139) );
  mux21 U4214 ( .Y(n7139), .A0(larray[110]), .A1(n____return437_2_), .S0(n6992) );
  inv01 U4215 ( .Y(n4561), .A(n7140) );
  mux21 U4216 ( .Y(n7140), .A0(larray[111]), .A1(n____return437_3_), .S0(n6992) );
  inv01 U4217 ( .Y(n4560), .A(n7141) );
  mux21 U4218 ( .Y(n7141), .A0(larray[112]), .A1(n____return437_4_), .S0(n6991) );
  inv01 U4219 ( .Y(n4559), .A(n7142) );
  mux21 U4220 ( .Y(n7142), .A0(larray[113]), .A1(n____return437_5_), .S0(n6992) );
  inv01 U4221 ( .Y(n4558), .A(n7143) );
  mux21 U4222 ( .Y(n7143), .A0(larray[114]), .A1(n____return437_6_), .S0(n6990) );
  inv01 U4223 ( .Y(n4557), .A(n7144) );
  mux21 U4224 ( .Y(n7144), .A0(larray[115]), .A1(n____return437_7_), .S0(n6991) );
  inv01 U4225 ( .Y(n4556), .A(n7145) );
  mux21 U4226 ( .Y(n7145), .A0(larray[116]), .A1(n____return437_8_), .S0(n6991) );
  inv01 U4227 ( .Y(n4555), .A(n7146) );
  mux21 U4228 ( .Y(n7146), .A0(larray[117]), .A1(n____return437_9_), .S0(n6991) );
  inv01 U4229 ( .Y(n4554), .A(n7147) );
  mux21 U4230 ( .Y(n7147), .A0(larray[118]), .A1(n____return437_10_), .S0(
        n6990) );
  inv01 U4231 ( .Y(n4553), .A(n7148) );
  mux21 U4232 ( .Y(n7148), .A0(larray[119]), .A1(n____return437_11_), .S0(
        n6990) );
  inv01 U4233 ( .Y(n7149), .A(larray[120]) );
  inv01 U4234 ( .Y(n7150), .A(larray[121]) );
  inv01 U4235 ( .Y(n7151), .A(larray[122]) );
  inv01 U4236 ( .Y(n7152), .A(larray[123]) );
  inv01 U4237 ( .Y(n7153), .A(larray[124]) );
  inv01 U4238 ( .Y(n7154), .A(larray[125]) );
  inv01 U4239 ( .Y(n4546), .A(n7155) );
  mux21 U4240 ( .Y(n7155), .A0(larray[126]), .A1(n____return792_0_), .S0(n6990) );
  inv01 U4241 ( .Y(n4545), .A(n7156) );
  mux21 U4242 ( .Y(n7156), .A0(larray[127]), .A1(n____return792_1_), .S0(n6991) );
  inv01 U4243 ( .Y(n4544), .A(n7157) );
  mux21 U4244 ( .Y(n7157), .A0(larray[128]), .A1(n____return792_2_), .S0(n6992) );
  inv01 U4245 ( .Y(n4543), .A(n7158) );
  mux21 U4246 ( .Y(n7158), .A0(larray[129]), .A1(n____return792_3_), .S0(n6991) );
  inv01 U4247 ( .Y(n4542), .A(n7159) );
  mux21 U4248 ( .Y(n7159), .A0(larray[130]), .A1(n____return792_4_), .S0(n6991) );
  inv01 U4249 ( .Y(n4541), .A(n7160) );
  mux21 U4250 ( .Y(n7160), .A0(larray[131]), .A1(n____return792_5_), .S0(n6991) );
  inv01 U4251 ( .Y(n4540), .A(n7161) );
  mux21 U4252 ( .Y(n7161), .A0(larray[132]), .A1(n____return792_6_), .S0(n6990) );
  inv01 U4253 ( .Y(n4539), .A(n7162) );
  mux21 U4254 ( .Y(n7162), .A0(larray[133]), .A1(n____return792_7_), .S0(n6991) );
  inv01 U4255 ( .Y(n4538), .A(n7163) );
  mux21 U4256 ( .Y(n7163), .A0(larray[134]), .A1(n____return792_8_), .S0(n6992) );
  inv01 U4257 ( .Y(n4537), .A(n7164) );
  mux21 U4258 ( .Y(n7164), .A0(larray[135]), .A1(n____return792_9_), .S0(n6990) );
  inv01 U4259 ( .Y(n4536), .A(n7165) );
  mux21 U4260 ( .Y(n7165), .A0(larray[136]), .A1(n____return792_10_), .S0(
        n6991) );
  inv01 U4261 ( .Y(n4535), .A(n7166) );
  mux21 U4262 ( .Y(n7166), .A0(larray[137]), .A1(n____return792_11_), .S0(
        n6991) );
  inv01 U4263 ( .Y(n7167), .A(larray[138]) );
  inv01 U4264 ( .Y(n7168), .A(larray[139]) );
  inv01 U4265 ( .Y(n7169), .A(larray[140]) );
  inv01 U4266 ( .Y(n7170), .A(larray[141]) );
  inv01 U4267 ( .Y(n7171), .A(larray[142]) );
  inv01 U4268 ( .Y(n7172), .A(larray[143]) );
  inv01 U4269 ( .Y(n7173), .A(larray[144]) );
  inv01 U4270 ( .Y(n7174), .A(larray[145]) );
  inv01 U4271 ( .Y(n7175), .A(larray[146]) );
  inv01 U4272 ( .Y(n7176), .A(larray[147]) );
  inv01 U4273 ( .Y(n7177), .A(larray[148]) );
  inv01 U4274 ( .Y(n7178), .A(larray[149]) );
  inv01 U4275 ( .Y(n4522), .A(n7179) );
  mux21 U4276 ( .Y(n7179), .A0(larray[150]), .A1(n____return1150_0_), .S0(
        n6992) );
  inv01 U4277 ( .Y(n4521), .A(n7180) );
  mux21 U4278 ( .Y(n7180), .A0(larray[151]), .A1(n____return1150_1_), .S0(
        n6990) );
  inv01 U4279 ( .Y(n4520), .A(n7181) );
  mux21 U4280 ( .Y(n7181), .A0(larray[152]), .A1(n____return1150_2_), .S0(
        n6992) );
  inv01 U4281 ( .Y(n4519), .A(n7182) );
  mux21 U4282 ( .Y(n7182), .A0(larray[153]), .A1(n____return1150_3_), .S0(
        n6991) );
  inv01 U4283 ( .Y(n4518), .A(n7183) );
  mux21 U4284 ( .Y(n7183), .A0(larray[154]), .A1(n____return1150_4_), .S0(
        n6991) );
  inv01 U4285 ( .Y(n4517), .A(n7184) );
  mux21 U4286 ( .Y(n7184), .A0(larray[155]), .A1(n____return1150_5_), .S0(
        n6991) );
  inv01 U4287 ( .Y(n4516), .A(n7185) );
  mux21 U4288 ( .Y(n7185), .A0(larray[156]), .A1(n____return1150_6_), .S0(
        n6992) );
  inv01 U4289 ( .Y(n4515), .A(n7186) );
  mux21 U4290 ( .Y(n7186), .A0(larray[157]), .A1(n____return1150_7_), .S0(
        n6990) );
  inv01 U4291 ( .Y(n4514), .A(n7187) );
  mux21 U4292 ( .Y(n7187), .A0(larray[158]), .A1(n____return1150_8_), .S0(
        n6990) );
  inv01 U4293 ( .Y(n4513), .A(n7188) );
  mux21 U4294 ( .Y(n7188), .A0(larray[159]), .A1(n____return1150_9_), .S0(
        n6992) );
  inv01 U4295 ( .Y(n4512), .A(n7189) );
  mux21 U4296 ( .Y(n7189), .A0(larray[160]), .A1(n____return1150_10_), .S0(
        n6992) );
  inv01 U4297 ( .Y(n4511), .A(n7190) );
  mux21 U4298 ( .Y(n7190), .A0(larray[161]), .A1(n____return1150_11_), .S0(
        n6990) );
  inv01 U4299 ( .Y(n7191), .A(larray[162]) );
  inv01 U4300 ( .Y(n7192), .A(larray[163]) );
  inv01 U4301 ( .Y(n7193), .A(larray[164]) );
  inv01 U4302 ( .Y(n7194), .A(larray[165]) );
  inv01 U4303 ( .Y(n7195), .A(larray[166]) );
  inv01 U4304 ( .Y(n7196), .A(larray[167]) );
  inv01 U4305 ( .Y(n4504), .A(n7197) );
  mux21 U4306 ( .Y(n7197), .A0(larray[168]), .A1(n____return1508_0_), .S0(
        n6990) );
  inv01 U4307 ( .Y(n4503), .A(n7198) );
  mux21 U4308 ( .Y(n7198), .A0(larray[169]), .A1(n____return1508_1_), .S0(
        n6990) );
  inv01 U4309 ( .Y(n4502), .A(n7199) );
  mux21 U4310 ( .Y(n7199), .A0(larray[170]), .A1(n____return1508_2_), .S0(
        n6992) );
  inv01 U4311 ( .Y(n4501), .A(n7200) );
  mux21 U4312 ( .Y(n7200), .A0(larray[171]), .A1(n____return1508_3_), .S0(
        n6991) );
  inv01 U4313 ( .Y(n4500), .A(n7201) );
  mux21 U4314 ( .Y(n7201), .A0(larray[172]), .A1(n____return1508_4_), .S0(
        n6990) );
  inv01 U4315 ( .Y(n4499), .A(n7202) );
  mux21 U4316 ( .Y(n7202), .A0(larray[173]), .A1(n____return1508_5_), .S0(
        n6992) );
  inv01 U4317 ( .Y(n4498), .A(n7203) );
  mux21 U4318 ( .Y(n7203), .A0(larray[174]), .A1(n____return1508_6_), .S0(
        n6990) );
  inv01 U4319 ( .Y(n4497), .A(n7204) );
  mux21 U4320 ( .Y(n7204), .A0(larray[175]), .A1(n____return1508_7_), .S0(
        n6992) );
  inv01 U4321 ( .Y(n4496), .A(n7205) );
  mux21 U4322 ( .Y(n7205), .A0(larray[176]), .A1(n____return1508_8_), .S0(
        n6990) );
  inv01 U4323 ( .Y(n4495), .A(n7206) );
  mux21 U4324 ( .Y(n7206), .A0(larray[177]), .A1(n____return1508_9_), .S0(
        n6992) );
  inv01 U4325 ( .Y(n4494), .A(n7207) );
  mux21 U4326 ( .Y(n7207), .A0(larray[178]), .A1(n____return1508_10_), .S0(
        n6992) );
  inv01 U4327 ( .Y(n4493), .A(n7208) );
  mux21 U4328 ( .Y(n7208), .A0(larray[179]), .A1(n____return1508_11_), .S0(
        n6991) );
  inv01 U4329 ( .Y(n7209), .A(larray[180]) );
  inv01 U4330 ( .Y(n7210), .A(larray[181]) );
  inv01 U4331 ( .Y(n7211), .A(larray[182]) );
  inv01 U4332 ( .Y(n7212), .A(larray[183]) );
  inv01 U4333 ( .Y(n7213), .A(larray[184]) );
  inv01 U4334 ( .Y(n7214), .A(larray[185]) );
  inv01 U4335 ( .Y(n7215), .A(larray[186]) );
  inv01 U4336 ( .Y(n7216), .A(larray[187]) );
  inv01 U4337 ( .Y(n7217), .A(larray[188]) );
  inv01 U4338 ( .Y(n7218), .A(larray[189]) );
  inv01 U4339 ( .Y(n7219), .A(larray[190]) );
  inv01 U4340 ( .Y(n7220), .A(larray[191]) );
  mux21 U4341 ( .Y(n4468), .A0(n7234), .A1(n7235), .S0(n6988) );
  mux21 U4342 ( .Y(n4467), .A0(n7236), .A1(n7237), .S0(n6987) );
  mux21 U4343 ( .Y(n4466), .A0(n7238), .A1(n7239), .S0(n6986) );
  mux21 U4344 ( .Y(n4465), .A0(n7240), .A1(n7241), .S0(n6988) );
  mux21 U4345 ( .Y(n4464), .A0(n7242), .A1(n7243), .S0(n6987) );
  mux21 U4346 ( .Y(n4462), .A0(n7246), .A1(n7247), .S0(n6988) );
  mux21 U4347 ( .Y(n4461), .A0(n7248), .A1(n7249), .S0(n6987) );
  mux21 U4348 ( .Y(n4460), .A0(n7250), .A1(n7251), .S0(n6986) );
  mux21 U4349 ( .Y(n4459), .A0(n7252), .A1(n7253), .S0(n6988) );
  mux21 U4350 ( .Y(n4458), .A0(n7254), .A1(n7255), .S0(n6987) );
  mux21 U4351 ( .Y(n4457), .A0(n7256), .A1(n7257), .S0(n6986) );
  mux21 U4352 ( .Y(n4450), .A0(n7264), .A1(n7265), .S0(n6988) );
  mux21 U4353 ( .Y(n4449), .A0(n7266), .A1(n7267), .S0(n6987) );
  mux21 U4354 ( .Y(n4447), .A0(n7270), .A1(n7271), .S0(n6988) );
  mux21 U4355 ( .Y(n4446), .A0(n7272), .A1(n7273), .S0(n6987) );
  mux21 U4356 ( .Y(n4445), .A0(n7274), .A1(n7275), .S0(n6986) );
  mux21 U4357 ( .Y(n4444), .A0(n7276), .A1(n7277), .S0(n6988) );
  mux21 U4358 ( .Y(n4443), .A0(n7278), .A1(n7279), .S0(n6987) );
  mux21 U4359 ( .Y(n4442), .A0(n7280), .A1(n7281), .S0(n6986) );
  mux21 U4360 ( .Y(n4441), .A0(n7282), .A1(n7283), .S0(n6988) );
  mux21 U4361 ( .Y(n4440), .A0(n7284), .A1(n7285), .S0(n6987) );
  mux21 U4362 ( .Y(n4439), .A0(n7286), .A1(n7287), .S0(n6986) );
  mux21 U4363 ( .Y(n4426), .A0(n7300), .A1(n7301), .S0(n6988) );
  mux21 U4364 ( .Y(n4425), .A0(n7302), .A1(n7303), .S0(n6987) );
  mux21 U4365 ( .Y(n4424), .A0(n7304), .A1(n7305), .S0(n6986) );
  mux21 U4366 ( .Y(n4423), .A0(n7306), .A1(n7307), .S0(n6988) );
  mux21 U4367 ( .Y(n4422), .A0(n7308), .A1(n7309), .S0(n6987) );
  mux21 U4368 ( .Y(n4420), .A0(n7312), .A1(n7313), .S0(n6988) );
  mux21 U4369 ( .Y(n4419), .A0(n7314), .A1(n7315), .S0(n6987) );
  mux21 U4370 ( .Y(n4418), .A0(n7316), .A1(n7317), .S0(n6986) );
  mux21 U4371 ( .Y(n4417), .A0(n7318), .A1(n7319), .S0(n6988) );
  mux21 U4372 ( .Y(n4416), .A0(n7320), .A1(n7321), .S0(n6987) );
  mux21 U4373 ( .Y(n4415), .A0(n7322), .A1(n7323), .S0(n6986) );
  mux21 U4374 ( .Y(n4407), .A0(n7332), .A1(n7333), .S0(n6987) );
  mux21 U4375 ( .Y(n4406), .A0(n7334), .A1(n7335), .S0(n6986) );
  mux21 U4376 ( .Y(n4405), .A0(n7336), .A1(n7337), .S0(n6988) );
  mux21 U4377 ( .Y(n4403), .A0(n7340), .A1(n7341), .S0(n6986) );
  mux21 U4378 ( .Y(n4402), .A0(n7342), .A1(n7343), .S0(n6988) );
  mux21 U4379 ( .Y(n4400), .A0(n7346), .A1(n7347), .S0(n6986) );
  mux21 U4380 ( .Y(n4399), .A0(n7348), .A1(n7349), .S0(n6988) );
  mux21 U4381 ( .Y(n4398), .A0(n7350), .A1(n7351), .S0(n6987) );
  mux21 U4382 ( .Y(n4397), .A0(n7352), .A1(n7353), .S0(n6986) );
  mux21 U4383 ( .Y(n4372), .A0(n7379), .A1(n7235), .S0(n6948) );
  inv01 U4384 ( .Y(n7235), .A(n____return437_0_) );
  mux21 U4385 ( .Y(n4371), .A0(n7380), .A1(n7237), .S0(n6950) );
  inv01 U4386 ( .Y(n7237), .A(n____return437_1_) );
  mux21 U4387 ( .Y(n4370), .A0(n7381), .A1(n7239), .S0(n6950) );
  inv01 U4388 ( .Y(n7239), .A(n____return437_2_) );
  mux21 U4389 ( .Y(n4369), .A0(n7382), .A1(n7241), .S0(n6948) );
  inv01 U4390 ( .Y(n7241), .A(n____return437_3_) );
  mux21 U4391 ( .Y(n4368), .A0(n7383), .A1(n7243), .S0(n6948) );
  inv01 U4392 ( .Y(n7243), .A(n____return437_4_) );
  mux21 U4393 ( .Y(n4367), .A0(n7384), .A1(n7245), .S0(n6948) );
  inv01 U4394 ( .Y(n7245), .A(n____return437_5_) );
  mux21 U4395 ( .Y(n4366), .A0(n7385), .A1(n7247), .S0(n6950) );
  inv01 U4396 ( .Y(n7247), .A(n____return437_6_) );
  mux21 U4397 ( .Y(n4365), .A0(n7386), .A1(n7249), .S0(n6950) );
  inv01 U4398 ( .Y(n7249), .A(n____return437_7_) );
  mux21 U4399 ( .Y(n4364), .A0(n7387), .A1(n7251), .S0(n6949) );
  inv01 U4400 ( .Y(n7251), .A(n____return437_8_) );
  mux21 U4401 ( .Y(n4363), .A0(n7388), .A1(n7253), .S0(n6949) );
  inv01 U4402 ( .Y(n7253), .A(n____return437_9_) );
  mux21 U4403 ( .Y(n4362), .A0(n7389), .A1(n7255), .S0(n6948) );
  inv01 U4404 ( .Y(n7255), .A(n____return437_10_) );
  inv01 U4405 ( .Y(n7257), .A(n____return437_11_) );
  mux21 U4406 ( .Y(n4354), .A0(n7397), .A1(n7265), .S0(n6948) );
  inv01 U4407 ( .Y(n7265), .A(n____return792_0_) );
  mux21 U4408 ( .Y(n4353), .A0(n7398), .A1(n7267), .S0(n6949) );
  inv01 U4409 ( .Y(n7267), .A(n____return792_1_) );
  mux21 U4410 ( .Y(n4352), .A0(n7399), .A1(n7269), .S0(n6949) );
  inv01 U4411 ( .Y(n7269), .A(n____return792_2_) );
  mux21 U4412 ( .Y(n4351), .A0(n7400), .A1(n7271), .S0(n6948) );
  inv01 U4413 ( .Y(n7271), .A(n____return792_3_) );
  inv01 U4414 ( .Y(n7273), .A(n____return792_4_) );
  mux21 U4415 ( .Y(n4349), .A0(n7402), .A1(n7275), .S0(n6950) );
  inv01 U4416 ( .Y(n7275), .A(n____return792_5_) );
  mux21 U4417 ( .Y(n4348), .A0(n7403), .A1(n7277), .S0(n6948) );
  inv01 U4418 ( .Y(n7277), .A(n____return792_6_) );
  mux21 U4419 ( .Y(n4347), .A0(n7404), .A1(n7279), .S0(n6949) );
  inv01 U4420 ( .Y(n7279), .A(n____return792_7_) );
  mux21 U4421 ( .Y(n4346), .A0(n7405), .A1(n7281), .S0(n6948) );
  inv01 U4422 ( .Y(n7281), .A(n____return792_8_) );
  mux21 U4423 ( .Y(n4345), .A0(n7406), .A1(n7283), .S0(n6950) );
  inv01 U4424 ( .Y(n7283), .A(n____return792_9_) );
  mux21 U4425 ( .Y(n4344), .A0(n7407), .A1(n7285), .S0(n6949) );
  inv01 U4426 ( .Y(n7285), .A(n____return792_10_) );
  mux21 U4427 ( .Y(n4343), .A0(n7408), .A1(n7287), .S0(n6950) );
  inv01 U4428 ( .Y(n7287), .A(n____return792_11_) );
  inv01 U4429 ( .Y(n7301), .A(n____return1150_0_) );
  mux21 U4430 ( .Y(n4329), .A0(n7422), .A1(n7303), .S0(n6949) );
  inv01 U4431 ( .Y(n7303), .A(n____return1150_1_) );
  inv01 U4432 ( .Y(n7305), .A(n____return1150_2_) );
  mux21 U4433 ( .Y(n4327), .A0(n7424), .A1(n7307), .S0(n6950) );
  inv01 U4434 ( .Y(n7307), .A(n____return1150_3_) );
  mux21 U4435 ( .Y(n4326), .A0(n7425), .A1(n7309), .S0(n6949) );
  inv01 U4436 ( .Y(n7309), .A(n____return1150_4_) );
  mux21 U4437 ( .Y(n4325), .A0(n7426), .A1(n7311), .S0(n6948) );
  inv01 U4438 ( .Y(n7311), .A(n____return1150_5_) );
  mux21 U4439 ( .Y(n4324), .A0(n7427), .A1(n7313), .S0(n6949) );
  inv01 U4440 ( .Y(n7313), .A(n____return1150_6_) );
  mux21 U4441 ( .Y(n4323), .A0(n7428), .A1(n7315), .S0(n6949) );
  inv01 U4442 ( .Y(n7315), .A(n____return1150_7_) );
  mux21 U4443 ( .Y(n4322), .A0(n7429), .A1(n7317), .S0(n6949) );
  inv01 U4444 ( .Y(n7317), .A(n____return1150_8_) );
  mux21 U4445 ( .Y(n4321), .A0(n7430), .A1(n7319), .S0(n6948) );
  inv01 U4446 ( .Y(n7319), .A(n____return1150_9_) );
  mux21 U4447 ( .Y(n4320), .A0(n7431), .A1(n7321), .S0(n6950) );
  inv01 U4448 ( .Y(n7321), .A(n____return1150_10_) );
  mux21 U4449 ( .Y(n4319), .A0(n7432), .A1(n7323), .S0(n6949) );
  inv01 U4450 ( .Y(n7323), .A(n____return1150_11_) );
  mux21 U4451 ( .Y(n4312), .A0(n7439), .A1(n7331), .S0(n6950) );
  inv01 U4452 ( .Y(n7331), .A(n____return1508_0_) );
  mux21 U4453 ( .Y(n4311), .A0(n7440), .A1(n7333), .S0(n6948) );
  inv01 U4454 ( .Y(n7333), .A(n____return1508_1_) );
  mux21 U4455 ( .Y(n4310), .A0(n7441), .A1(n7335), .S0(n6949) );
  inv01 U4456 ( .Y(n7335), .A(n____return1508_2_) );
  mux21 U4457 ( .Y(n4309), .A0(n7442), .A1(n7337), .S0(n6950) );
  inv01 U4458 ( .Y(n7337), .A(n____return1508_3_) );
  mux21 U4459 ( .Y(n4308), .A0(n7443), .A1(n7339), .S0(n6948) );
  inv01 U4460 ( .Y(n7339), .A(n____return1508_4_) );
  mux21 U4461 ( .Y(n4307), .A0(n7444), .A1(n7341), .S0(n6948) );
  inv01 U4462 ( .Y(n7341), .A(n____return1508_5_) );
  mux21 U4463 ( .Y(n4306), .A0(n7445), .A1(n7343), .S0(n6950) );
  inv01 U4464 ( .Y(n7343), .A(n____return1508_6_) );
  mux21 U4465 ( .Y(n4305), .A0(n7446), .A1(n7345), .S0(n6950) );
  inv01 U4466 ( .Y(n7345), .A(n____return1508_7_) );
  mux21 U4467 ( .Y(n4304), .A0(n7447), .A1(n7347), .S0(n6950) );
  inv01 U4468 ( .Y(n7347), .A(n____return1508_8_) );
  mux21 U4469 ( .Y(n4303), .A0(n7448), .A1(n7349), .S0(n6949) );
  inv01 U4470 ( .Y(n7349), .A(n____return1508_9_) );
  mux21 U4471 ( .Y(n4302), .A0(n7449), .A1(n7351), .S0(n6950) );
  inv01 U4472 ( .Y(n7351), .A(n____return1508_10_) );
  inv01 U4473 ( .Y(n7353), .A(n____return1508_11_) );
  aoi22 U4474 ( .Y(n7463), .A0(n7464), .A1(n6891), .B0(n6936), .B1(n7465) );
  ao22 U4475 ( .Y(n7464), .A0(n7366), .A1(n6936), .B0(s_state), .B1(n6949) );
  nand02 U4476 ( .Y(n7467), .A0(n6945), .A1(n6303) );
  nand02 U4477 ( .Y(n7466), .A0(n7465), .A1(n6994) );
  ao21 U4478 ( .Y(n7465), .A0(n6890), .A1(n7221), .B0(n6995) );
  nand02 U4479 ( .Y(n7469), .A0(n6303), .A1(n6892) );
  nand03 U4480 ( .Y(n6996), .A0(n7221), .A1(n7366), .A2(n6936) );
  nand02 U4481 ( .Y(n7468), .A0(n6995), .A1(n6994) );
  aoi22 U4482 ( .Y(member996_4__4_), .A0(n3564), .A1(n6940), .B0(n3576), .B1(
        n7366) );
  aoi22 U4483 ( .Y(member996_4__1_), .A0(n3561), .A1(n6940), .B0(n3573), .B1(
        n7366) );
  aoi22 U4484 ( .Y(member638_2__3_), .A0(n3569), .A1(n6940), .B0(n3581), .B1(
        n7366) );
  aoi22 U4485 ( .Y(member360_1__3_), .A0(n3545), .A1(n6946), .B0(n3557), .B1(
        n7221) );
  aoi22 U4486 ( .Y(member360_1__1_), .A0(n3543), .A1(n6946), .B0(n3555), .B1(
        n7221) );
  inv01 U4487 ( .Y(n7348), .A(larray[273]) );
  inv01 U4488 ( .Y(n7448), .A(larray[369]) );
  inv01 U4489 ( .Y(n7346), .A(larray[272]) );
  inv01 U4490 ( .Y(n7447), .A(larray[368]) );
  inv01 U4491 ( .Y(n7344), .A(larray[271]) );
  inv01 U4492 ( .Y(n7446), .A(larray[367]) );
  inv01 U4493 ( .Y(n7342), .A(larray[270]) );
  inv01 U4494 ( .Y(n7445), .A(larray[366]) );
  inv01 U4495 ( .Y(n7340), .A(larray[269]) );
  inv01 U4496 ( .Y(n7444), .A(larray[365]) );
  inv01 U4497 ( .Y(n7338), .A(larray[268]) );
  inv01 U4498 ( .Y(n7443), .A(larray[364]) );
  inv01 U4499 ( .Y(n7336), .A(larray[267]) );
  inv01 U4500 ( .Y(n7442), .A(larray[363]) );
  inv01 U4501 ( .Y(n7334), .A(larray[266]) );
  inv01 U4502 ( .Y(n7441), .A(larray[362]) );
  inv01 U4503 ( .Y(n7365), .A(larray[287]) );
  inv01 U4504 ( .Y(n7462), .A(larray[383]) );
  inv01 U4505 ( .Y(n7364), .A(larray[286]) );
  inv01 U4506 ( .Y(n7461), .A(larray[382]) );
  inv01 U4507 ( .Y(n7363), .A(larray[285]) );
  inv01 U4508 ( .Y(n7460), .A(larray[381]) );
  inv01 U4509 ( .Y(n7362), .A(larray[284]) );
  inv01 U4510 ( .Y(n7459), .A(larray[380]) );
  inv01 U4511 ( .Y(n7332), .A(larray[265]) );
  inv01 U4512 ( .Y(n7440), .A(larray[361]) );
  inv01 U4513 ( .Y(n7361), .A(larray[283]) );
  inv01 U4514 ( .Y(n7458), .A(larray[379]) );
  inv01 U4515 ( .Y(n7360), .A(larray[282]) );
  inv01 U4516 ( .Y(n7457), .A(larray[378]) );
  inv01 U4517 ( .Y(n7359), .A(larray[281]) );
  inv01 U4518 ( .Y(n7456), .A(larray[377]) );
  inv01 U4519 ( .Y(n7358), .A(larray[280]) );
  inv01 U4520 ( .Y(n7455), .A(larray[376]) );
  inv01 U4521 ( .Y(n7357), .A(larray[279]) );
  inv01 U4522 ( .Y(n7454), .A(larray[375]) );
  inv01 U4523 ( .Y(n7356), .A(larray[278]) );
  inv01 U4524 ( .Y(n7453), .A(larray[374]) );
  inv01 U4525 ( .Y(n7355), .A(larray[277]) );
  inv01 U4526 ( .Y(n7452), .A(larray[373]) );
  inv01 U4527 ( .Y(n7354), .A(larray[276]) );
  inv01 U4528 ( .Y(n7451), .A(larray[372]) );
  inv01 U4529 ( .Y(n7352), .A(larray[275]) );
  inv01 U4530 ( .Y(n7450), .A(larray[371]) );
  inv01 U4531 ( .Y(n7350), .A(larray[274]) );
  inv01 U4532 ( .Y(n7449), .A(larray[370]) );
  inv01 U4533 ( .Y(n7330), .A(larray[264]) );
  inv01 U4534 ( .Y(n7439), .A(larray[360]) );
  inv01 U4535 ( .Y(n7306), .A(larray[249]) );
  inv01 U4536 ( .Y(n7424), .A(larray[345]) );
  inv01 U4537 ( .Y(n7304), .A(larray[248]) );
  inv01 U4538 ( .Y(n7423), .A(larray[344]) );
  inv01 U4539 ( .Y(n7302), .A(larray[247]) );
  inv01 U4540 ( .Y(n7422), .A(larray[343]) );
  inv01 U4541 ( .Y(n7300), .A(larray[246]) );
  inv01 U4542 ( .Y(n7421), .A(larray[342]) );
  inv01 U4543 ( .Y(n7299), .A(larray[245]) );
  inv01 U4544 ( .Y(n7420), .A(larray[341]) );
  inv01 U4545 ( .Y(n7298), .A(larray[244]) );
  inv01 U4546 ( .Y(n7419), .A(larray[340]) );
  inv01 U4547 ( .Y(n7297), .A(larray[243]) );
  inv01 U4548 ( .Y(n7418), .A(larray[339]) );
  inv01 U4549 ( .Y(n7296), .A(larray[242]) );
  inv01 U4550 ( .Y(n7417), .A(larray[338]) );
  inv01 U4551 ( .Y(n7329), .A(larray[263]) );
  inv01 U4552 ( .Y(n7438), .A(larray[359]) );
  inv01 U4553 ( .Y(n7328), .A(larray[262]) );
  inv01 U4554 ( .Y(n7437), .A(larray[358]) );
  inv01 U4555 ( .Y(n7327), .A(larray[261]) );
  inv01 U4556 ( .Y(n7436), .A(larray[357]) );
  inv01 U4557 ( .Y(n7326), .A(larray[260]) );
  inv01 U4558 ( .Y(n7435), .A(larray[356]) );
  inv01 U4559 ( .Y(n7295), .A(larray[241]) );
  inv01 U4560 ( .Y(n7416), .A(larray[337]) );
  inv01 U4561 ( .Y(n7325), .A(larray[259]) );
  inv01 U4562 ( .Y(n7434), .A(larray[355]) );
  inv01 U4563 ( .Y(n7324), .A(larray[258]) );
  inv01 U4564 ( .Y(n7433), .A(larray[354]) );
  inv01 U4565 ( .Y(n7322), .A(larray[257]) );
  inv01 U4566 ( .Y(n7432), .A(larray[353]) );
  inv01 U4567 ( .Y(n7320), .A(larray[256]) );
  inv01 U4568 ( .Y(n7431), .A(larray[352]) );
  inv01 U4569 ( .Y(n7318), .A(larray[255]) );
  inv01 U4570 ( .Y(n7430), .A(larray[351]) );
  inv01 U4571 ( .Y(n7316), .A(larray[254]) );
  inv01 U4572 ( .Y(n7429), .A(larray[350]) );
  inv01 U4573 ( .Y(n7314), .A(larray[253]) );
  inv01 U4574 ( .Y(n7428), .A(larray[349]) );
  inv01 U4575 ( .Y(n7312), .A(larray[252]) );
  inv01 U4576 ( .Y(n7427), .A(larray[348]) );
  inv01 U4577 ( .Y(n7310), .A(larray[251]) );
  inv01 U4578 ( .Y(n7426), .A(larray[347]) );
  inv01 U4579 ( .Y(n7308), .A(larray[250]) );
  inv01 U4580 ( .Y(n7425), .A(larray[346]) );
  inv01 U4581 ( .Y(n7294), .A(larray[240]) );
  inv01 U4582 ( .Y(n7415), .A(larray[336]) );
  inv01 U4583 ( .Y(n7270), .A(larray[225]) );
  inv01 U4584 ( .Y(n7400), .A(larray[321]) );
  inv01 U4585 ( .Y(n7268), .A(larray[224]) );
  inv01 U4586 ( .Y(n7399), .A(larray[320]) );
  inv01 U4587 ( .Y(n7266), .A(larray[223]) );
  inv01 U4588 ( .Y(n7398), .A(larray[319]) );
  inv01 U4589 ( .Y(n7264), .A(larray[222]) );
  inv01 U4590 ( .Y(n7397), .A(larray[318]) );
  inv01 U4591 ( .Y(n7263), .A(larray[221]) );
  inv01 U4592 ( .Y(n7396), .A(larray[317]) );
  inv01 U4593 ( .Y(n7262), .A(larray[220]) );
  inv01 U4594 ( .Y(n7395), .A(larray[316]) );
  inv01 U4595 ( .Y(n7261), .A(larray[219]) );
  inv01 U4596 ( .Y(n7394), .A(larray[315]) );
  inv01 U4597 ( .Y(n7260), .A(larray[218]) );
  inv01 U4598 ( .Y(n7393), .A(larray[314]) );
  inv01 U4599 ( .Y(n7293), .A(larray[239]) );
  inv01 U4600 ( .Y(n7414), .A(larray[335]) );
  inv01 U4601 ( .Y(n7292), .A(larray[238]) );
  inv01 U4602 ( .Y(n7413), .A(larray[334]) );
  inv01 U4603 ( .Y(n7291), .A(larray[237]) );
  inv01 U4604 ( .Y(n7412), .A(larray[333]) );
  inv01 U4605 ( .Y(n7290), .A(larray[236]) );
  inv01 U4606 ( .Y(n7411), .A(larray[332]) );
  inv01 U4607 ( .Y(n7259), .A(larray[217]) );
  inv01 U4608 ( .Y(n7392), .A(larray[313]) );
  inv01 U4609 ( .Y(n7289), .A(larray[235]) );
  inv01 U4610 ( .Y(n7410), .A(larray[331]) );
  inv01 U4611 ( .Y(n7288), .A(larray[234]) );
  inv01 U4612 ( .Y(n7409), .A(larray[330]) );
  inv01 U4613 ( .Y(n7286), .A(larray[233]) );
  inv01 U4614 ( .Y(n7408), .A(larray[329]) );
  inv01 U4615 ( .Y(n7284), .A(larray[232]) );
  inv01 U4616 ( .Y(n7407), .A(larray[328]) );
  inv01 U4617 ( .Y(n7282), .A(larray[231]) );
  inv01 U4618 ( .Y(n7406), .A(larray[327]) );
  inv01 U4619 ( .Y(n7280), .A(larray[230]) );
  inv01 U4620 ( .Y(n7405), .A(larray[326]) );
  inv01 U4621 ( .Y(n7278), .A(larray[229]) );
  inv01 U4622 ( .Y(n7404), .A(larray[325]) );
  inv01 U4623 ( .Y(n7276), .A(larray[228]) );
  inv01 U4624 ( .Y(n7403), .A(larray[324]) );
  inv01 U4625 ( .Y(n7274), .A(larray[227]) );
  inv01 U4626 ( .Y(n7402), .A(larray[323]) );
  inv01 U4627 ( .Y(n7272), .A(larray[226]) );
  inv01 U4628 ( .Y(n7401), .A(larray[322]) );
  inv01 U4629 ( .Y(n7258), .A(larray[216]) );
  inv01 U4630 ( .Y(n7391), .A(larray[312]) );
  inv01 U4631 ( .Y(n7231), .A(larray[201]) );
  inv01 U4632 ( .Y(n7376), .A(larray[297]) );
  inv01 U4633 ( .Y(n7230), .A(larray[200]) );
  inv01 U4634 ( .Y(n7375), .A(larray[296]) );
  inv01 U4635 ( .Y(n7229), .A(larray[199]) );
  inv01 U4636 ( .Y(n7374), .A(larray[295]) );
  inv01 U4637 ( .Y(n7228), .A(larray[198]) );
  inv01 U4638 ( .Y(n7373), .A(larray[294]) );
  inv01 U4639 ( .Y(n7227), .A(larray[197]) );
  inv01 U4640 ( .Y(n7372), .A(larray[293]) );
  inv01 U4641 ( .Y(n7226), .A(larray[196]) );
  inv01 U4642 ( .Y(n7371), .A(larray[292]) );
  inv01 U4643 ( .Y(n7225), .A(larray[195]) );
  inv01 U4644 ( .Y(n7370), .A(larray[291]) );
  inv01 U4645 ( .Y(n7224), .A(larray[194]) );
  inv01 U4646 ( .Y(n7369), .A(larray[290]) );
  inv01 U4647 ( .Y(n7256), .A(larray[215]) );
  inv01 U4648 ( .Y(n7390), .A(larray[311]) );
  inv01 U4649 ( .Y(n7254), .A(larray[214]) );
  inv01 U4650 ( .Y(n7389), .A(larray[310]) );
  inv01 U4651 ( .Y(n7252), .A(larray[213]) );
  inv01 U4652 ( .Y(n7388), .A(larray[309]) );
  inv01 U4653 ( .Y(n7250), .A(larray[212]) );
  inv01 U4654 ( .Y(n7387), .A(larray[308]) );
  inv01 U4655 ( .Y(n7223), .A(larray[193]) );
  inv01 U4656 ( .Y(n7368), .A(larray[289]) );
  inv01 U4657 ( .Y(n7248), .A(larray[211]) );
  inv01 U4658 ( .Y(n7386), .A(larray[307]) );
  inv01 U4659 ( .Y(n7246), .A(larray[210]) );
  inv01 U4660 ( .Y(n7385), .A(larray[306]) );
  inv01 U4661 ( .Y(n7244), .A(larray[209]) );
  inv01 U4662 ( .Y(n7384), .A(larray[305]) );
  inv01 U4663 ( .Y(n7242), .A(larray[208]) );
  inv01 U4664 ( .Y(n7383), .A(larray[304]) );
  inv01 U4665 ( .Y(n7240), .A(larray[207]) );
  inv01 U4666 ( .Y(n7382), .A(larray[303]) );
  inv01 U4667 ( .Y(n7238), .A(larray[206]) );
  inv01 U4668 ( .Y(n7381), .A(larray[302]) );
  inv01 U4669 ( .Y(n7236), .A(larray[205]) );
  inv01 U4670 ( .Y(n7380), .A(larray[301]) );
  inv01 U4671 ( .Y(n7234), .A(larray[204]) );
  inv01 U4672 ( .Y(n7379), .A(larray[300]) );
  inv01 U4673 ( .Y(n7233), .A(larray[203]) );
  inv01 U4674 ( .Y(n7378), .A(larray[299]) );
  inv01 U4675 ( .Y(n7232), .A(larray[202]) );
  inv01 U4676 ( .Y(n7377), .A(larray[298]) );
  nor02 U4677 ( .Y(n7022), .A0(n7221), .A1(n6938) );
  inv01 U4678 ( .Y(n7222), .A(larray[192]) );
  nand02 U4679 ( .Y(n7024), .A0(n6939), .A1(n6946) );
  inv01 U4680 ( .Y(n7367), .A(larray[288]) );
  nand02 U4681 ( .Y(n7026), .A0(n6938), .A1(n7221) );
  aoi22 U4682 ( .Y(n7534), .A0(n7366), .A1(n6946), .B0(n6940), .B1(n7221) );
  mul_24_DW01_add_48_2 add_0_root_add_223_plus_plus_228 ( .A({
        n____return2374_47_, n____return2374_46_, n____return2374_45_, 
        n____return2374_44_, n____return2374_43_, n____return2374_42_, 
        n____return2374_41_, n____return2374_40_, n____return2374_39_, 
        n____return2374_38_, n____return2374_37_, n____return2374_36_, 
        n____return2374_35_, n____return2374_34_, n____return2374_33_, 
        n____return2374_32_, n____return2374_31_, n____return2374_30_, 
        n____return2374_29_, n____return2374_28_, n____return2374_27_, 
        n____return2374_26_, n____return2374_25_, n____return2374_24_, 
        n____return2374_23_, n____return2374_22_, n____return2374_21_, 
        n____return2374_20_, n____return2374_19_, n____return2374_18_, 
        n____return2374_17_, n____return2374_16_, n____return2374_15_, 
        n____return2374_14_, n____return2374_13_, n____return2374_12_, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        n____return2414_36_, n____return2414_35_, n____return2414_34_, 
        n____return2414_33_, n____return2414_32_, n____return2414_31_, 
        n____return2414_30_, n____return2414_29_, n____return2414_28_, 
        n____return2414_27_, n____return2414_26_, n____return2414_25_, 
        n____return2414_24_, n____return2414_23_, n____return2414_22_, 
        n____return2414_21_, n____return2414_20_, n____return2414_19_, 
        n____return2414_18_, n____return2414_17_, n____return2414_16_, 
        n____return2414_15_, n____return2414_14_, n____return2414_13_, 
        n____return2414_12_, n____return2414_11_, n____return2414_10_, 
        n____return2414_9_, n____return2414_8_, n____return2414_7_, 
        n____return2414_6_, n____return2414_5_, n____return2414_4_, 
        n____return2414_3_, n____return2414_2_, n____return2414_1_, 
        n____return2414_0_}), .CI(1'b0), .SUM(fract_o) );
  mul_24_DW01_add_48_1 add_1_root_add_223_plus_plus_228 ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, prod_a_b_2__35_, 
        prod_a_b_2__34_, prod_a_b_2__33_, prod_a_b_2__32_, prod_a_b_2__31_, 
        prod_a_b_2__30_, prod_a_b_2__29_, prod_a_b_2__28_, prod_a_b_2__27_, 
        prod_a_b_2__26_, prod_a_b_2__25_, prod_a_b_2__24_, prod_a_b_2__23_, 
        prod_a_b_2__22_, prod_a_b_2__21_, prod_a_b_2__20_, prod_a_b_2__19_, 
        prod_a_b_2__18_, prod_a_b_2__17_, prod_a_b_2__16_, prod_a_b_2__15_, 
        prod_a_b_2__14_, prod_a_b_2__13_, prod_a_b_2__12_, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        prod_a_b_3__23_, prod_a_b_3__22_, prod_a_b_3__21_, prod_a_b_3__20_, 
        prod_a_b_3__19_, prod_a_b_3__18_, prod_a_b_3__17_, prod_a_b_3__16_, 
        prod_a_b_3__15_, prod_a_b_3__14_, prod_a_b_3__13_, prod_a_b_3__12_, 
        prod_a_b_3__11_, prod_a_b_3__10_, prod_a_b_3__9_, prod_a_b_3__8_, 
        prod_a_b_3__7_, prod_a_b_3__6_, prod_a_b_3__5_, prod_a_b_3__4_, 
        prod_a_b_3__3_, prod_a_b_3__2_, prod_a_b_3__1_, prod_a_b_3__0_}), .CI(
        1'b0), .SUM({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, n____return2414_36_, n____return2414_35_, 
        n____return2414_34_, n____return2414_33_, n____return2414_32_, 
        n____return2414_31_, n____return2414_30_, n____return2414_29_, 
        n____return2414_28_, n____return2414_27_, n____return2414_26_, 
        n____return2414_25_, n____return2414_24_, n____return2414_23_, 
        n____return2414_22_, n____return2414_21_, n____return2414_20_, 
        n____return2414_19_, n____return2414_18_, n____return2414_17_, 
        n____return2414_16_, n____return2414_15_, n____return2414_14_, 
        n____return2414_13_, n____return2414_12_, n____return2414_11_, 
        n____return2414_10_, n____return2414_9_, n____return2414_8_, 
        n____return2414_7_, n____return2414_6_, n____return2414_5_, 
        n____return2414_4_, n____return2414_3_, n____return2414_2_, 
        n____return2414_1_, n____return2414_0_}) );
  mul_24_DW01_add_48_0 add_2_root_add_223_plus_plus_228 ( .A({prod_a_b_0__47_, 
        prod_a_b_0__46_, prod_a_b_0__45_, prod_a_b_0__44_, prod_a_b_0__43_, 
        prod_a_b_0__42_, prod_a_b_0__41_, prod_a_b_0__40_, prod_a_b_0__39_, 
        prod_a_b_0__38_, prod_a_b_0__37_, prod_a_b_0__36_, prod_a_b_0__35_, 
        prod_a_b_0__34_, prod_a_b_0__33_, prod_a_b_0__32_, prod_a_b_0__31_, 
        prod_a_b_0__30_, prod_a_b_0__29_, prod_a_b_0__28_, prod_a_b_0__27_, 
        prod_a_b_0__26_, prod_a_b_0__25_, prod_a_b_0__24_, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        prod_a_b_1__35_, prod_a_b_1__34_, prod_a_b_1__33_, prod_a_b_1__32_, 
        prod_a_b_1__31_, prod_a_b_1__30_, prod_a_b_1__29_, prod_a_b_1__28_, 
        prod_a_b_1__27_, prod_a_b_1__26_, prod_a_b_1__25_, prod_a_b_1__24_, 
        prod_a_b_1__23_, prod_a_b_1__22_, prod_a_b_1__21_, prod_a_b_1__20_, 
        prod_a_b_1__19_, prod_a_b_1__18_, prod_a_b_1__17_, prod_a_b_1__16_, 
        prod_a_b_1__15_, prod_a_b_1__14_, prod_a_b_1__13_, prod_a_b_1__12_, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({n____return2374_47_, n____return2374_46_, 
        n____return2374_45_, n____return2374_44_, n____return2374_43_, 
        n____return2374_42_, n____return2374_41_, n____return2374_40_, 
        n____return2374_39_, n____return2374_38_, n____return2374_37_, 
        n____return2374_36_, n____return2374_35_, n____return2374_34_, 
        n____return2374_33_, n____return2374_32_, n____return2374_31_, 
        n____return2374_30_, n____return2374_29_, n____return2374_28_, 
        n____return2374_27_, n____return2374_26_, n____return2374_25_, 
        n____return2374_24_, n____return2374_23_, n____return2374_22_, 
        n____return2374_21_, n____return2374_20_, n____return2374_19_, 
        n____return2374_18_, n____return2374_17_, n____return2374_16_, 
        n____return2374_15_, n____return2374_14_, n____return2374_13_, 
        n____return2374_12_, SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23}) );
  mul_24_DW01_add_24_2 add_0_root_add_208_plus_plus_218 ( .A({
        n____return1960_23_, n____return1960_22_, n____return1960_21_, 
        n____return1960_20_, n____return1960_19_, n____return1960_18_, 
        n____return1960_17_, n____return1960_16_, n____return1960_15_, 
        n____return1960_14_, n____return1960_13_, n____return1960_12_, 
        n____return1960_11_, n____return1960_10_, n____return1960_9_, 
        n____return1960_8_, n____return1960_7_, n____return1960_6_, 
        n____return1960_5_, n____return1960_4_, n____return1960_3_, 
        n____return1960_2_, n____return1960_1_, n____return1960_0_}), .B({
        n____return2087_23_, n____return2087_22_, n____return2087_21_, 
        n____return2087_20_, n____return2087_19_, n____return2087_18_, 
        n____return2087_17_, n____return2087_16_, n____return2087_15_, 
        n____return2087_14_, n____return2087_13_, n____return2087_12_, 
        n____return2087_11_, n____return2087_10_, n____return2087_9_, 
        n____return2087_8_, n____return2087_7_, n____return2087_6_, 
        n____return2087_5_, n____return2087_4_, n____return2087_3_, 
        n____return2087_2_, n____return2087_1_, n____return2087_0_}), .CI(1'b0), .SUM({n____return2214_23_, n____return2214_22_, n____return2214_21_, 
        n____return2214_20_, n____return2214_19_, n____return2214_18_, 
        n____return2214_17_, n____return2214_16_, n____return2214_15_, 
        n____return2214_14_, n____return2214_13_, n____return2214_12_, 
        n____return2214_11_, n____return2214_10_, n____return2214_9_, 
        n____return2214_8_, n____return2214_7_, n____return2214_6_, 
        n____return2214_5_, n____return2214_4_, n____return2214_3_, 
        n____return2214_2_, n____return2214_1_, n____return2214_0_}) );
  mul_24_DW01_add_24_1 add_1_root_add_208_plus_plus_218 ( .A({
        member2010_2__23_, member2010_2__22_, member2010_2__21_, 
        member2010_2__20_, member2010_2__19_, member2010_2__18_, 
        member2010_2__17_, member2010_2__16_, member2010_2__15_, 
        member2010_2__14_, member2010_2__13_, member2010_2__12_, 
        member2010_2__11_, member2010_2__10_, member2010_2__9_, 
        member2010_2__8_, member2010_2__7_, member2010_2__6_, member2010_2__5_, 
        member2010_2__4_, member2010_2__3_, member2010_2__2_, member2010_2__1_, 
        member2010_2__0_}), .B({member2137_3__23_, member2137_3__22_, 
        member2137_3__21_, member2137_3__20_, member2137_3__19_, 
        member2137_3__18_, member2137_3__17_, member2137_3__16_, 
        member2137_3__15_, member2137_3__14_, member2137_3__13_, 
        member2137_3__12_, member2137_3__11_, member2137_3__10_, 
        member2137_3__9_, member2137_3__8_, member2137_3__7_, member2137_3__6_, 
        member2137_3__5_, member2137_3__4_, member2137_3__3_, member2137_3__2_, 
        member2137_3__1_, member2137_3__0_}), .CI(1'b0), .SUM({
        n____return2087_23_, n____return2087_22_, n____return2087_21_, 
        n____return2087_20_, n____return2087_19_, n____return2087_18_, 
        n____return2087_17_, n____return2087_16_, n____return2087_15_, 
        n____return2087_14_, n____return2087_13_, n____return2087_12_, 
        n____return2087_11_, n____return2087_10_, n____return2087_9_, 
        n____return2087_8_, n____return2087_7_, n____return2087_6_, 
        n____return2087_5_, n____return2087_4_, n____return2087_3_, 
        n____return2087_2_, n____return2087_1_, n____return2087_0_}) );
  mul_24_DW01_add_24_0 add_2_root_add_208_plus_plus_218 ( .A({
        member1796_0__23_, member1796_0__22_, member1796_0__21_, 
        member1796_0__20_, member1796_0__19_, member1796_0__18_, 
        member1796_0__17_, member1796_0__16_, member1796_0__15_, 
        member1796_0__14_, member1796_0__13_, member1796_0__12_, 
        member1796_0__11_, member1796_0__10_, member1796_0__9_, 
        member1796_0__8_, member1796_0__7_, member1796_0__6_, member1796_0__5_, 
        member1796_0__4_, member1796_0__3_, member1796_0__2_, member1796_0__1_, 
        member1796_0__0_}), .B({member1883_1__23_, member1883_1__22_, 
        member1883_1__21_, member1883_1__20_, member1883_1__19_, 
        member1883_1__18_, member1883_1__17_, member1883_1__16_, 
        member1883_1__15_, member1883_1__14_, member1883_1__13_, 
        member1883_1__12_, member1883_1__11_, member1883_1__10_, 
        member1883_1__9_, member1883_1__8_, member1883_1__7_, member1883_1__6_, 
        member1883_1__5_, member1883_1__4_, member1883_1__3_, member1883_1__2_, 
        member1883_1__1_, member1883_1__0_}), .CI(1'b0), .SUM({
        n____return1960_23_, n____return1960_22_, n____return1960_21_, 
        n____return1960_20_, n____return1960_19_, n____return1960_18_, 
        n____return1960_17_, n____return1960_16_, n____return1960_15_, 
        n____return1960_14_, n____return1960_13_, n____return1960_12_, 
        n____return1960_11_, n____return1960_10_, n____return1960_9_, 
        n____return1960_8_, n____return1960_7_, n____return1960_6_, 
        n____return1960_5_, n____return1960_4_, n____return1960_3_, 
        n____return1960_2_, n____return1960_1_, n____return1960_0_}) );
  mul_24_DW02_mult_6_6_3 mul_197_mult_mult ( .A({n6910, n6893, n6934, n6894, 
        n6898, n6924}), .B({n6920, n6900, n6922, n6914, n6902, n6916}), .TC(
        1'b0), .PRODUCT({n____return1508_11_, n____return1508_10_, 
        n____return1508_9_, n____return1508_8_, n____return1508_7_, 
        n____return1508_6_, n____return1508_5_, n____return1508_4_, 
        n____return1508_3_, n____return1508_2_, n____return1508_1_, 
        n____return1508_0_}) );
  mul_24_DW02_mult_6_6_2 mul_196_mult_mult ( .A({n6910, n6893, n6934, n6894, 
        n6898, n6924}), .B({n6908, n6918, n6896, n6904, n6895, n6906}), .TC(
        1'b0), .PRODUCT({n____return1150_11_, n____return1150_10_, 
        n____return1150_9_, n____return1150_8_, n____return1150_7_, 
        n____return1150_6_, n____return1150_5_, n____return1150_4_, 
        n____return1150_3_, n____return1150_2_, n____return1150_1_, 
        n____return1150_0_}) );
  mul_24_DW02_mult_6_6_1 mul_195_mult_mult ( .A({n6932, n6926, n6897, n6928, 
        n6912, n6930}), .B({n6920, n6900, n6922, n6914, n6902, n6916}), .TC(
        1'b0), .PRODUCT({n____return792_11_, n____return792_10_, 
        n____return792_9_, n____return792_8_, n____return792_7_, 
        n____return792_6_, n____return792_5_, n____return792_4_, 
        n____return792_3_, n____return792_2_, n____return792_1_, 
        n____return792_0_}) );
  mul_24_DW02_mult_6_6_0 mul_194_mult_mult ( .A({n6932, n6926, n6897, n6928, 
        n6912, n6930}), .B({n6908, n6918, n6896, n6904, n6895, n6906}), .TC(
        1'b0), .PRODUCT({n____return437_11_, n____return437_10_, 
        n____return437_9_, n____return437_8_, n____return437_7_, 
        n____return437_6_, n____return437_5_, n____return437_4_, 
        n____return437_3_, n____return437_2_, n____return437_1_, 
        n____return437_0_}) );
endmodule


module serial_mul_DW01_add_48_0 ( A, B, CI, SUM, CO );
  input [47:0] A;
  input [47:0] B;
  output [47:0] SUM;
  input CI;
  output CO;
  wire   carry_47_, carry_46_, carry_45_, carry_44_, carry_43_, carry_42_,
         carry_41_, carry_40_, carry_39_, carry_38_, carry_37_, carry_36_,
         carry_35_, carry_34_, carry_33_, carry_32_, carry_31_, carry_30_,
         carry_29_, carry_28_, carry_27_, carry_26_, carry_25_, carry_24_,
         carry_23_, carry_22_, carry_21_, carry_20_, carry_19_, carry_18_,
         carry_17_, carry_16_, carry_15_, carry_14_, carry_13_, carry_12_,
         carry_11_, carry_10_, carry_9_, carry_8_, carry_7_, carry_6_,
         carry_5_, carry_4_, carry_3_, carry_2_, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621;

  nand02 U4 ( .Y(SUM[46]), .A0(n1), .A1(n2) );
  nand02 U5 ( .Y(carry_47_), .A0(n3), .A1(n4) );
  inv01 U6 ( .Y(n5), .A(carry_46_) );
  inv01 U7 ( .Y(n6), .A(A[46]) );
  inv01 U8 ( .Y(n7), .A(B[46]) );
  nand02 U9 ( .Y(n8), .A0(n6), .A1(n9) );
  nand02 U10 ( .Y(n10), .A0(n7), .A1(n11) );
  nand02 U11 ( .Y(n12), .A0(n7), .A1(n13) );
  nand02 U12 ( .Y(n14), .A0(carry_46_), .A1(n15) );
  nand02 U13 ( .Y(n16), .A0(A[46]), .A1(carry_46_) );
  nand02 U14 ( .Y(n17), .A0(B[46]), .A1(carry_46_) );
  nand02 U15 ( .Y(n3), .A0(B[46]), .A1(A[46]) );
  nand02 U16 ( .Y(n18), .A0(B[46]), .A1(n5) );
  inv01 U17 ( .Y(n9), .A(n18) );
  nand02 U18 ( .Y(n19), .A0(A[46]), .A1(n5) );
  inv01 U19 ( .Y(n11), .A(n19) );
  nand02 U20 ( .Y(n20), .A0(carry_46_), .A1(n6) );
  inv01 U21 ( .Y(n13), .A(n20) );
  nand02 U22 ( .Y(n21), .A0(B[46]), .A1(A[46]) );
  inv01 U23 ( .Y(n15), .A(n21) );
  nand02 U24 ( .Y(n22), .A0(n8), .A1(n10) );
  inv01 U25 ( .Y(n1), .A(n22) );
  nand02 U26 ( .Y(n23), .A0(n12), .A1(n14) );
  inv01 U27 ( .Y(n2), .A(n23) );
  nand02 U28 ( .Y(n24), .A0(n16), .A1(n17) );
  inv01 U29 ( .Y(n4), .A(n24) );
  nand02 U30 ( .Y(n25), .A0(A[0]), .A1(B[0]) );
  inv02 U31 ( .Y(n26), .A(n25) );
  inv01 U32 ( .Y(SUM[45]), .A(n27) );
  inv02 U33 ( .Y(carry_46_), .A(n28) );
  inv02 U34 ( .Y(n29), .A(B[45]) );
  inv02 U35 ( .Y(n30), .A(A[45]) );
  inv02 U36 ( .Y(n31), .A(carry_45_) );
  nor02 U37 ( .Y(n32), .A0(n29), .A1(n33) );
  nor02 U38 ( .Y(n34), .A0(n30), .A1(n35) );
  nor02 U39 ( .Y(n36), .A0(n31), .A1(n37) );
  nor02 U40 ( .Y(n38), .A0(n31), .A1(n39) );
  nor02 U41 ( .Y(n27), .A0(n40), .A1(n41) );
  nor02 U42 ( .Y(n42), .A0(n30), .A1(n31) );
  nor02 U43 ( .Y(n43), .A0(n29), .A1(n31) );
  nor02 U44 ( .Y(n44), .A0(n29), .A1(n30) );
  nor02 U45 ( .Y(n28), .A0(n44), .A1(n45) );
  nor02 U46 ( .Y(n46), .A0(A[45]), .A1(carry_45_) );
  inv01 U47 ( .Y(n33), .A(n46) );
  nor02 U48 ( .Y(n47), .A0(B[45]), .A1(carry_45_) );
  inv01 U49 ( .Y(n35), .A(n47) );
  nor02 U50 ( .Y(n48), .A0(B[45]), .A1(A[45]) );
  inv01 U51 ( .Y(n37), .A(n48) );
  nor02 U52 ( .Y(n49), .A0(n29), .A1(n30) );
  inv01 U53 ( .Y(n39), .A(n49) );
  nor02 U54 ( .Y(n50), .A0(n32), .A1(n34) );
  inv01 U55 ( .Y(n40), .A(n50) );
  nor02 U56 ( .Y(n51), .A0(n36), .A1(n38) );
  inv01 U57 ( .Y(n41), .A(n51) );
  nor02 U58 ( .Y(n52), .A0(n42), .A1(n43) );
  inv01 U59 ( .Y(n45), .A(n52) );
  inv01 U60 ( .Y(SUM[44]), .A(n53) );
  inv02 U61 ( .Y(carry_45_), .A(n54) );
  inv02 U62 ( .Y(n55), .A(B[44]) );
  inv02 U63 ( .Y(n56), .A(A[44]) );
  inv02 U64 ( .Y(n57), .A(carry_44_) );
  nor02 U65 ( .Y(n58), .A0(n55), .A1(n59) );
  nor02 U66 ( .Y(n60), .A0(n56), .A1(n61) );
  nor02 U67 ( .Y(n62), .A0(n57), .A1(n63) );
  nor02 U68 ( .Y(n64), .A0(n57), .A1(n65) );
  nor02 U69 ( .Y(n53), .A0(n66), .A1(n67) );
  nor02 U70 ( .Y(n68), .A0(n56), .A1(n57) );
  nor02 U71 ( .Y(n69), .A0(n55), .A1(n57) );
  nor02 U72 ( .Y(n70), .A0(n55), .A1(n56) );
  nor02 U73 ( .Y(n54), .A0(n70), .A1(n71) );
  nor02 U74 ( .Y(n72), .A0(A[44]), .A1(carry_44_) );
  inv01 U75 ( .Y(n59), .A(n72) );
  nor02 U76 ( .Y(n73), .A0(B[44]), .A1(carry_44_) );
  inv01 U77 ( .Y(n61), .A(n73) );
  nor02 U78 ( .Y(n74), .A0(B[44]), .A1(A[44]) );
  inv01 U79 ( .Y(n63), .A(n74) );
  nor02 U80 ( .Y(n75), .A0(n55), .A1(n56) );
  inv01 U81 ( .Y(n65), .A(n75) );
  nor02 U82 ( .Y(n76), .A0(n58), .A1(n60) );
  inv01 U83 ( .Y(n66), .A(n76) );
  nor02 U84 ( .Y(n77), .A0(n62), .A1(n64) );
  inv01 U85 ( .Y(n67), .A(n77) );
  nor02 U86 ( .Y(n78), .A0(n68), .A1(n69) );
  inv01 U87 ( .Y(n71), .A(n78) );
  inv01 U88 ( .Y(SUM[43]), .A(n79) );
  inv02 U89 ( .Y(carry_44_), .A(n80) );
  inv02 U90 ( .Y(n81), .A(B[43]) );
  inv02 U91 ( .Y(n82), .A(A[43]) );
  inv02 U92 ( .Y(n83), .A(carry_43_) );
  nor02 U93 ( .Y(n84), .A0(n81), .A1(n85) );
  nor02 U94 ( .Y(n86), .A0(n82), .A1(n87) );
  nor02 U95 ( .Y(n88), .A0(n83), .A1(n89) );
  nor02 U96 ( .Y(n90), .A0(n83), .A1(n91) );
  nor02 U97 ( .Y(n79), .A0(n92), .A1(n93) );
  nor02 U98 ( .Y(n94), .A0(n82), .A1(n83) );
  nor02 U99 ( .Y(n95), .A0(n81), .A1(n83) );
  nor02 U100 ( .Y(n96), .A0(n81), .A1(n82) );
  nor02 U101 ( .Y(n80), .A0(n96), .A1(n97) );
  nor02 U102 ( .Y(n98), .A0(A[43]), .A1(carry_43_) );
  inv01 U103 ( .Y(n85), .A(n98) );
  nor02 U104 ( .Y(n99), .A0(B[43]), .A1(carry_43_) );
  inv01 U105 ( .Y(n87), .A(n99) );
  nor02 U106 ( .Y(n100), .A0(B[43]), .A1(A[43]) );
  inv01 U107 ( .Y(n89), .A(n100) );
  nor02 U108 ( .Y(n101), .A0(n81), .A1(n82) );
  inv01 U109 ( .Y(n91), .A(n101) );
  nor02 U110 ( .Y(n102), .A0(n84), .A1(n86) );
  inv01 U111 ( .Y(n92), .A(n102) );
  nor02 U112 ( .Y(n103), .A0(n88), .A1(n90) );
  inv01 U113 ( .Y(n93), .A(n103) );
  nor02 U114 ( .Y(n104), .A0(n94), .A1(n95) );
  inv01 U115 ( .Y(n97), .A(n104) );
  inv01 U116 ( .Y(SUM[42]), .A(n105) );
  inv02 U117 ( .Y(carry_43_), .A(n106) );
  inv02 U118 ( .Y(n107), .A(B[42]) );
  inv02 U119 ( .Y(n108), .A(A[42]) );
  inv02 U120 ( .Y(n109), .A(carry_42_) );
  nor02 U121 ( .Y(n110), .A0(n107), .A1(n111) );
  nor02 U122 ( .Y(n112), .A0(n108), .A1(n113) );
  nor02 U123 ( .Y(n114), .A0(n109), .A1(n115) );
  nor02 U124 ( .Y(n116), .A0(n109), .A1(n117) );
  nor02 U125 ( .Y(n105), .A0(n118), .A1(n119) );
  nor02 U126 ( .Y(n120), .A0(n108), .A1(n109) );
  nor02 U127 ( .Y(n121), .A0(n107), .A1(n109) );
  nor02 U128 ( .Y(n122), .A0(n107), .A1(n108) );
  nor02 U129 ( .Y(n106), .A0(n122), .A1(n123) );
  nor02 U130 ( .Y(n124), .A0(A[42]), .A1(carry_42_) );
  inv01 U131 ( .Y(n111), .A(n124) );
  nor02 U132 ( .Y(n125), .A0(B[42]), .A1(carry_42_) );
  inv01 U133 ( .Y(n113), .A(n125) );
  nor02 U134 ( .Y(n126), .A0(B[42]), .A1(A[42]) );
  inv01 U135 ( .Y(n115), .A(n126) );
  nor02 U136 ( .Y(n127), .A0(n107), .A1(n108) );
  inv01 U137 ( .Y(n117), .A(n127) );
  nor02 U138 ( .Y(n128), .A0(n110), .A1(n112) );
  inv01 U139 ( .Y(n118), .A(n128) );
  nor02 U140 ( .Y(n129), .A0(n114), .A1(n116) );
  inv01 U141 ( .Y(n119), .A(n129) );
  nor02 U142 ( .Y(n130), .A0(n120), .A1(n121) );
  inv01 U143 ( .Y(n123), .A(n130) );
  inv01 U144 ( .Y(SUM[41]), .A(n131) );
  inv02 U145 ( .Y(carry_42_), .A(n132) );
  inv02 U146 ( .Y(n133), .A(B[41]) );
  inv02 U147 ( .Y(n134), .A(A[41]) );
  inv02 U148 ( .Y(n135), .A(carry_41_) );
  nor02 U149 ( .Y(n136), .A0(n133), .A1(n137) );
  nor02 U150 ( .Y(n138), .A0(n134), .A1(n139) );
  nor02 U151 ( .Y(n140), .A0(n135), .A1(n141) );
  nor02 U152 ( .Y(n142), .A0(n135), .A1(n143) );
  nor02 U153 ( .Y(n131), .A0(n144), .A1(n145) );
  nor02 U154 ( .Y(n146), .A0(n134), .A1(n135) );
  nor02 U155 ( .Y(n147), .A0(n133), .A1(n135) );
  nor02 U156 ( .Y(n148), .A0(n133), .A1(n134) );
  nor02 U157 ( .Y(n132), .A0(n148), .A1(n149) );
  nor02 U158 ( .Y(n150), .A0(A[41]), .A1(carry_41_) );
  inv01 U159 ( .Y(n137), .A(n150) );
  nor02 U160 ( .Y(n151), .A0(B[41]), .A1(carry_41_) );
  inv01 U161 ( .Y(n139), .A(n151) );
  nor02 U162 ( .Y(n152), .A0(B[41]), .A1(A[41]) );
  inv01 U163 ( .Y(n141), .A(n152) );
  nor02 U164 ( .Y(n153), .A0(n133), .A1(n134) );
  inv01 U165 ( .Y(n143), .A(n153) );
  nor02 U166 ( .Y(n154), .A0(n136), .A1(n138) );
  inv01 U167 ( .Y(n144), .A(n154) );
  nor02 U168 ( .Y(n155), .A0(n140), .A1(n142) );
  inv01 U169 ( .Y(n145), .A(n155) );
  nor02 U170 ( .Y(n156), .A0(n146), .A1(n147) );
  inv01 U171 ( .Y(n149), .A(n156) );
  inv01 U172 ( .Y(SUM[40]), .A(n157) );
  inv02 U173 ( .Y(carry_41_), .A(n158) );
  inv02 U174 ( .Y(n159), .A(B[40]) );
  inv02 U175 ( .Y(n160), .A(A[40]) );
  inv02 U176 ( .Y(n161), .A(carry_40_) );
  nor02 U177 ( .Y(n162), .A0(n159), .A1(n163) );
  nor02 U178 ( .Y(n164), .A0(n160), .A1(n165) );
  nor02 U179 ( .Y(n166), .A0(n161), .A1(n167) );
  nor02 U180 ( .Y(n168), .A0(n161), .A1(n169) );
  nor02 U181 ( .Y(n157), .A0(n170), .A1(n171) );
  nor02 U182 ( .Y(n172), .A0(n160), .A1(n161) );
  nor02 U183 ( .Y(n173), .A0(n159), .A1(n161) );
  nor02 U184 ( .Y(n174), .A0(n159), .A1(n160) );
  nor02 U185 ( .Y(n158), .A0(n174), .A1(n175) );
  nor02 U186 ( .Y(n176), .A0(A[40]), .A1(carry_40_) );
  inv01 U187 ( .Y(n163), .A(n176) );
  nor02 U188 ( .Y(n177), .A0(B[40]), .A1(carry_40_) );
  inv01 U189 ( .Y(n165), .A(n177) );
  nor02 U190 ( .Y(n178), .A0(B[40]), .A1(A[40]) );
  inv01 U191 ( .Y(n167), .A(n178) );
  nor02 U192 ( .Y(n179), .A0(n159), .A1(n160) );
  inv01 U193 ( .Y(n169), .A(n179) );
  nor02 U194 ( .Y(n180), .A0(n162), .A1(n164) );
  inv01 U195 ( .Y(n170), .A(n180) );
  nor02 U196 ( .Y(n181), .A0(n166), .A1(n168) );
  inv01 U197 ( .Y(n171), .A(n181) );
  nor02 U198 ( .Y(n182), .A0(n172), .A1(n173) );
  inv01 U199 ( .Y(n175), .A(n182) );
  inv01 U200 ( .Y(SUM[39]), .A(n183) );
  inv02 U201 ( .Y(carry_40_), .A(n184) );
  inv02 U202 ( .Y(n185), .A(B[39]) );
  inv02 U203 ( .Y(n186), .A(A[39]) );
  inv02 U204 ( .Y(n187), .A(carry_39_) );
  nor02 U205 ( .Y(n188), .A0(n185), .A1(n189) );
  nor02 U206 ( .Y(n190), .A0(n186), .A1(n191) );
  nor02 U207 ( .Y(n192), .A0(n187), .A1(n193) );
  nor02 U208 ( .Y(n194), .A0(n187), .A1(n195) );
  nor02 U209 ( .Y(n183), .A0(n196), .A1(n197) );
  nor02 U210 ( .Y(n198), .A0(n186), .A1(n187) );
  nor02 U211 ( .Y(n199), .A0(n185), .A1(n187) );
  nor02 U212 ( .Y(n200), .A0(n185), .A1(n186) );
  nor02 U213 ( .Y(n184), .A0(n200), .A1(n201) );
  nor02 U214 ( .Y(n202), .A0(A[39]), .A1(carry_39_) );
  inv01 U215 ( .Y(n189), .A(n202) );
  nor02 U216 ( .Y(n203), .A0(B[39]), .A1(carry_39_) );
  inv01 U217 ( .Y(n191), .A(n203) );
  nor02 U218 ( .Y(n204), .A0(B[39]), .A1(A[39]) );
  inv01 U219 ( .Y(n193), .A(n204) );
  nor02 U220 ( .Y(n205), .A0(n185), .A1(n186) );
  inv01 U221 ( .Y(n195), .A(n205) );
  nor02 U222 ( .Y(n206), .A0(n188), .A1(n190) );
  inv01 U223 ( .Y(n196), .A(n206) );
  nor02 U224 ( .Y(n207), .A0(n192), .A1(n194) );
  inv01 U225 ( .Y(n197), .A(n207) );
  nor02 U226 ( .Y(n208), .A0(n198), .A1(n199) );
  inv01 U227 ( .Y(n201), .A(n208) );
  inv01 U228 ( .Y(SUM[38]), .A(n209) );
  inv02 U229 ( .Y(carry_39_), .A(n210) );
  inv02 U230 ( .Y(n211), .A(B[38]) );
  inv02 U231 ( .Y(n212), .A(A[38]) );
  inv02 U232 ( .Y(n213), .A(carry_38_) );
  nor02 U233 ( .Y(n214), .A0(n211), .A1(n215) );
  nor02 U234 ( .Y(n216), .A0(n212), .A1(n217) );
  nor02 U235 ( .Y(n218), .A0(n213), .A1(n219) );
  nor02 U236 ( .Y(n220), .A0(n213), .A1(n221) );
  nor02 U237 ( .Y(n209), .A0(n222), .A1(n223) );
  nor02 U238 ( .Y(n224), .A0(n212), .A1(n213) );
  nor02 U239 ( .Y(n225), .A0(n211), .A1(n213) );
  nor02 U240 ( .Y(n226), .A0(n211), .A1(n212) );
  nor02 U241 ( .Y(n210), .A0(n226), .A1(n227) );
  nor02 U242 ( .Y(n228), .A0(A[38]), .A1(carry_38_) );
  inv01 U243 ( .Y(n215), .A(n228) );
  nor02 U244 ( .Y(n229), .A0(B[38]), .A1(carry_38_) );
  inv01 U245 ( .Y(n217), .A(n229) );
  nor02 U246 ( .Y(n230), .A0(B[38]), .A1(A[38]) );
  inv01 U247 ( .Y(n219), .A(n230) );
  nor02 U248 ( .Y(n231), .A0(n211), .A1(n212) );
  inv01 U249 ( .Y(n221), .A(n231) );
  nor02 U250 ( .Y(n232), .A0(n214), .A1(n216) );
  inv01 U251 ( .Y(n222), .A(n232) );
  nor02 U252 ( .Y(n233), .A0(n218), .A1(n220) );
  inv01 U253 ( .Y(n223), .A(n233) );
  nor02 U254 ( .Y(n234), .A0(n224), .A1(n225) );
  inv01 U255 ( .Y(n227), .A(n234) );
  inv01 U256 ( .Y(SUM[37]), .A(n235) );
  inv02 U257 ( .Y(carry_38_), .A(n236) );
  inv02 U258 ( .Y(n237), .A(B[37]) );
  inv02 U259 ( .Y(n238), .A(A[37]) );
  inv02 U260 ( .Y(n239), .A(carry_37_) );
  nor02 U261 ( .Y(n240), .A0(n237), .A1(n241) );
  nor02 U262 ( .Y(n242), .A0(n238), .A1(n243) );
  nor02 U263 ( .Y(n244), .A0(n239), .A1(n245) );
  nor02 U264 ( .Y(n246), .A0(n239), .A1(n247) );
  nor02 U265 ( .Y(n235), .A0(n248), .A1(n249) );
  nor02 U266 ( .Y(n250), .A0(n238), .A1(n239) );
  nor02 U267 ( .Y(n251), .A0(n237), .A1(n239) );
  nor02 U268 ( .Y(n252), .A0(n237), .A1(n238) );
  nor02 U269 ( .Y(n236), .A0(n252), .A1(n253) );
  nor02 U270 ( .Y(n254), .A0(A[37]), .A1(carry_37_) );
  inv01 U271 ( .Y(n241), .A(n254) );
  nor02 U272 ( .Y(n255), .A0(B[37]), .A1(carry_37_) );
  inv01 U273 ( .Y(n243), .A(n255) );
  nor02 U274 ( .Y(n256), .A0(B[37]), .A1(A[37]) );
  inv01 U275 ( .Y(n245), .A(n256) );
  nor02 U276 ( .Y(n257), .A0(n237), .A1(n238) );
  inv01 U277 ( .Y(n247), .A(n257) );
  nor02 U278 ( .Y(n258), .A0(n240), .A1(n242) );
  inv01 U279 ( .Y(n248), .A(n258) );
  nor02 U280 ( .Y(n259), .A0(n244), .A1(n246) );
  inv01 U281 ( .Y(n249), .A(n259) );
  nor02 U282 ( .Y(n260), .A0(n250), .A1(n251) );
  inv01 U283 ( .Y(n253), .A(n260) );
  inv01 U284 ( .Y(SUM[36]), .A(n261) );
  inv02 U285 ( .Y(carry_37_), .A(n262) );
  inv02 U286 ( .Y(n263), .A(B[36]) );
  inv02 U287 ( .Y(n264), .A(A[36]) );
  inv02 U288 ( .Y(n265), .A(carry_36_) );
  nor02 U289 ( .Y(n266), .A0(n263), .A1(n267) );
  nor02 U290 ( .Y(n268), .A0(n264), .A1(n269) );
  nor02 U291 ( .Y(n270), .A0(n265), .A1(n271) );
  nor02 U292 ( .Y(n272), .A0(n265), .A1(n273) );
  nor02 U293 ( .Y(n261), .A0(n274), .A1(n275) );
  nor02 U294 ( .Y(n276), .A0(n264), .A1(n265) );
  nor02 U295 ( .Y(n277), .A0(n263), .A1(n265) );
  nor02 U296 ( .Y(n278), .A0(n263), .A1(n264) );
  nor02 U297 ( .Y(n262), .A0(n278), .A1(n279) );
  nor02 U298 ( .Y(n280), .A0(A[36]), .A1(carry_36_) );
  inv01 U299 ( .Y(n267), .A(n280) );
  nor02 U300 ( .Y(n281), .A0(B[36]), .A1(carry_36_) );
  inv01 U301 ( .Y(n269), .A(n281) );
  nor02 U302 ( .Y(n282), .A0(B[36]), .A1(A[36]) );
  inv01 U303 ( .Y(n271), .A(n282) );
  nor02 U304 ( .Y(n283), .A0(n263), .A1(n264) );
  inv01 U305 ( .Y(n273), .A(n283) );
  nor02 U306 ( .Y(n284), .A0(n266), .A1(n268) );
  inv01 U307 ( .Y(n274), .A(n284) );
  nor02 U308 ( .Y(n285), .A0(n270), .A1(n272) );
  inv01 U309 ( .Y(n275), .A(n285) );
  nor02 U310 ( .Y(n286), .A0(n276), .A1(n277) );
  inv01 U311 ( .Y(n279), .A(n286) );
  inv01 U312 ( .Y(SUM[35]), .A(n287) );
  inv02 U313 ( .Y(carry_36_), .A(n288) );
  inv02 U314 ( .Y(n289), .A(B[35]) );
  inv02 U315 ( .Y(n290), .A(A[35]) );
  inv02 U316 ( .Y(n291), .A(carry_35_) );
  nor02 U317 ( .Y(n292), .A0(n289), .A1(n293) );
  nor02 U318 ( .Y(n294), .A0(n290), .A1(n295) );
  nor02 U319 ( .Y(n296), .A0(n291), .A1(n297) );
  nor02 U320 ( .Y(n298), .A0(n291), .A1(n299) );
  nor02 U321 ( .Y(n287), .A0(n300), .A1(n301) );
  nor02 U322 ( .Y(n302), .A0(n290), .A1(n291) );
  nor02 U323 ( .Y(n303), .A0(n289), .A1(n291) );
  nor02 U324 ( .Y(n304), .A0(n289), .A1(n290) );
  nor02 U325 ( .Y(n288), .A0(n304), .A1(n305) );
  nor02 U326 ( .Y(n306), .A0(A[35]), .A1(carry_35_) );
  inv01 U327 ( .Y(n293), .A(n306) );
  nor02 U328 ( .Y(n307), .A0(B[35]), .A1(carry_35_) );
  inv01 U329 ( .Y(n295), .A(n307) );
  nor02 U330 ( .Y(n308), .A0(B[35]), .A1(A[35]) );
  inv01 U331 ( .Y(n297), .A(n308) );
  nor02 U332 ( .Y(n309), .A0(n289), .A1(n290) );
  inv01 U333 ( .Y(n299), .A(n309) );
  nor02 U334 ( .Y(n310), .A0(n292), .A1(n294) );
  inv01 U335 ( .Y(n300), .A(n310) );
  nor02 U336 ( .Y(n311), .A0(n296), .A1(n298) );
  inv01 U337 ( .Y(n301), .A(n311) );
  nor02 U338 ( .Y(n312), .A0(n302), .A1(n303) );
  inv01 U339 ( .Y(n305), .A(n312) );
  inv01 U340 ( .Y(SUM[34]), .A(n313) );
  inv02 U341 ( .Y(carry_35_), .A(n314) );
  inv02 U342 ( .Y(n315), .A(B[34]) );
  inv02 U343 ( .Y(n316), .A(A[34]) );
  inv02 U344 ( .Y(n317), .A(carry_34_) );
  nor02 U345 ( .Y(n318), .A0(n315), .A1(n319) );
  nor02 U346 ( .Y(n320), .A0(n316), .A1(n321) );
  nor02 U347 ( .Y(n322), .A0(n317), .A1(n323) );
  nor02 U348 ( .Y(n324), .A0(n317), .A1(n325) );
  nor02 U349 ( .Y(n313), .A0(n326), .A1(n327) );
  nor02 U350 ( .Y(n328), .A0(n316), .A1(n317) );
  nor02 U351 ( .Y(n329), .A0(n315), .A1(n317) );
  nor02 U352 ( .Y(n330), .A0(n315), .A1(n316) );
  nor02 U353 ( .Y(n314), .A0(n330), .A1(n331) );
  nor02 U354 ( .Y(n332), .A0(A[34]), .A1(carry_34_) );
  inv01 U355 ( .Y(n319), .A(n332) );
  nor02 U356 ( .Y(n333), .A0(B[34]), .A1(carry_34_) );
  inv01 U357 ( .Y(n321), .A(n333) );
  nor02 U358 ( .Y(n334), .A0(B[34]), .A1(A[34]) );
  inv01 U359 ( .Y(n323), .A(n334) );
  nor02 U360 ( .Y(n335), .A0(n315), .A1(n316) );
  inv01 U361 ( .Y(n325), .A(n335) );
  nor02 U362 ( .Y(n336), .A0(n318), .A1(n320) );
  inv01 U363 ( .Y(n326), .A(n336) );
  nor02 U364 ( .Y(n337), .A0(n322), .A1(n324) );
  inv01 U365 ( .Y(n327), .A(n337) );
  nor02 U366 ( .Y(n338), .A0(n328), .A1(n329) );
  inv01 U367 ( .Y(n331), .A(n338) );
  inv01 U368 ( .Y(SUM[33]), .A(n339) );
  inv02 U369 ( .Y(carry_34_), .A(n340) );
  inv02 U370 ( .Y(n341), .A(B[33]) );
  inv02 U371 ( .Y(n342), .A(A[33]) );
  inv02 U372 ( .Y(n343), .A(carry_33_) );
  nor02 U373 ( .Y(n344), .A0(n341), .A1(n345) );
  nor02 U374 ( .Y(n346), .A0(n342), .A1(n347) );
  nor02 U375 ( .Y(n348), .A0(n343), .A1(n349) );
  nor02 U376 ( .Y(n350), .A0(n343), .A1(n351) );
  nor02 U377 ( .Y(n339), .A0(n352), .A1(n353) );
  nor02 U378 ( .Y(n354), .A0(n342), .A1(n343) );
  nor02 U379 ( .Y(n355), .A0(n341), .A1(n343) );
  nor02 U380 ( .Y(n356), .A0(n341), .A1(n342) );
  nor02 U381 ( .Y(n340), .A0(n356), .A1(n357) );
  nor02 U382 ( .Y(n358), .A0(A[33]), .A1(carry_33_) );
  inv01 U383 ( .Y(n345), .A(n358) );
  nor02 U384 ( .Y(n359), .A0(B[33]), .A1(carry_33_) );
  inv01 U385 ( .Y(n347), .A(n359) );
  nor02 U386 ( .Y(n360), .A0(B[33]), .A1(A[33]) );
  inv01 U387 ( .Y(n349), .A(n360) );
  nor02 U388 ( .Y(n361), .A0(n341), .A1(n342) );
  inv01 U389 ( .Y(n351), .A(n361) );
  nor02 U390 ( .Y(n362), .A0(n344), .A1(n346) );
  inv01 U391 ( .Y(n352), .A(n362) );
  nor02 U392 ( .Y(n363), .A0(n348), .A1(n350) );
  inv01 U393 ( .Y(n353), .A(n363) );
  nor02 U394 ( .Y(n364), .A0(n354), .A1(n355) );
  inv01 U395 ( .Y(n357), .A(n364) );
  inv01 U396 ( .Y(SUM[32]), .A(n365) );
  inv02 U397 ( .Y(carry_33_), .A(n366) );
  inv02 U398 ( .Y(n367), .A(B[32]) );
  inv02 U399 ( .Y(n368), .A(A[32]) );
  inv02 U400 ( .Y(n369), .A(carry_32_) );
  nor02 U401 ( .Y(n370), .A0(n367), .A1(n371) );
  nor02 U402 ( .Y(n372), .A0(n368), .A1(n373) );
  nor02 U403 ( .Y(n374), .A0(n369), .A1(n375) );
  nor02 U404 ( .Y(n376), .A0(n369), .A1(n377) );
  nor02 U405 ( .Y(n365), .A0(n378), .A1(n379) );
  nor02 U406 ( .Y(n380), .A0(n368), .A1(n369) );
  nor02 U407 ( .Y(n381), .A0(n367), .A1(n369) );
  nor02 U408 ( .Y(n382), .A0(n367), .A1(n368) );
  nor02 U409 ( .Y(n366), .A0(n382), .A1(n383) );
  nor02 U410 ( .Y(n384), .A0(A[32]), .A1(carry_32_) );
  inv01 U411 ( .Y(n371), .A(n384) );
  nor02 U412 ( .Y(n385), .A0(B[32]), .A1(carry_32_) );
  inv01 U413 ( .Y(n373), .A(n385) );
  nor02 U414 ( .Y(n386), .A0(B[32]), .A1(A[32]) );
  inv01 U415 ( .Y(n375), .A(n386) );
  nor02 U416 ( .Y(n387), .A0(n367), .A1(n368) );
  inv01 U417 ( .Y(n377), .A(n387) );
  nor02 U418 ( .Y(n388), .A0(n370), .A1(n372) );
  inv01 U419 ( .Y(n378), .A(n388) );
  nor02 U420 ( .Y(n389), .A0(n374), .A1(n376) );
  inv01 U421 ( .Y(n379), .A(n389) );
  nor02 U422 ( .Y(n390), .A0(n380), .A1(n381) );
  inv01 U423 ( .Y(n383), .A(n390) );
  inv01 U424 ( .Y(SUM[31]), .A(n391) );
  inv02 U425 ( .Y(carry_32_), .A(n392) );
  inv02 U426 ( .Y(n393), .A(B[31]) );
  inv02 U427 ( .Y(n394), .A(A[31]) );
  inv02 U428 ( .Y(n395), .A(carry_31_) );
  nor02 U429 ( .Y(n396), .A0(n393), .A1(n397) );
  nor02 U430 ( .Y(n398), .A0(n394), .A1(n399) );
  nor02 U431 ( .Y(n400), .A0(n395), .A1(n401) );
  nor02 U432 ( .Y(n402), .A0(n395), .A1(n403) );
  nor02 U433 ( .Y(n391), .A0(n404), .A1(n405) );
  nor02 U434 ( .Y(n406), .A0(n394), .A1(n395) );
  nor02 U435 ( .Y(n407), .A0(n393), .A1(n395) );
  nor02 U436 ( .Y(n408), .A0(n393), .A1(n394) );
  nor02 U437 ( .Y(n392), .A0(n408), .A1(n409) );
  nor02 U438 ( .Y(n410), .A0(A[31]), .A1(carry_31_) );
  inv01 U439 ( .Y(n397), .A(n410) );
  nor02 U440 ( .Y(n411), .A0(B[31]), .A1(carry_31_) );
  inv01 U441 ( .Y(n399), .A(n411) );
  nor02 U442 ( .Y(n412), .A0(B[31]), .A1(A[31]) );
  inv01 U443 ( .Y(n401), .A(n412) );
  nor02 U444 ( .Y(n413), .A0(n393), .A1(n394) );
  inv01 U445 ( .Y(n403), .A(n413) );
  nor02 U446 ( .Y(n414), .A0(n396), .A1(n398) );
  inv01 U447 ( .Y(n404), .A(n414) );
  nor02 U448 ( .Y(n415), .A0(n400), .A1(n402) );
  inv01 U449 ( .Y(n405), .A(n415) );
  nor02 U450 ( .Y(n416), .A0(n406), .A1(n407) );
  inv01 U451 ( .Y(n409), .A(n416) );
  inv01 U452 ( .Y(SUM[30]), .A(n417) );
  inv02 U453 ( .Y(carry_31_), .A(n418) );
  inv02 U454 ( .Y(n419), .A(B[30]) );
  inv02 U455 ( .Y(n420), .A(A[30]) );
  inv02 U456 ( .Y(n421), .A(carry_30_) );
  nor02 U457 ( .Y(n422), .A0(n419), .A1(n423) );
  nor02 U458 ( .Y(n424), .A0(n420), .A1(n425) );
  nor02 U459 ( .Y(n426), .A0(n421), .A1(n427) );
  nor02 U460 ( .Y(n428), .A0(n421), .A1(n429) );
  nor02 U461 ( .Y(n417), .A0(n430), .A1(n431) );
  nor02 U462 ( .Y(n432), .A0(n420), .A1(n421) );
  nor02 U463 ( .Y(n433), .A0(n419), .A1(n421) );
  nor02 U464 ( .Y(n434), .A0(n419), .A1(n420) );
  nor02 U465 ( .Y(n418), .A0(n434), .A1(n435) );
  nor02 U466 ( .Y(n436), .A0(A[30]), .A1(carry_30_) );
  inv01 U467 ( .Y(n423), .A(n436) );
  nor02 U468 ( .Y(n437), .A0(B[30]), .A1(carry_30_) );
  inv01 U469 ( .Y(n425), .A(n437) );
  nor02 U470 ( .Y(n438), .A0(B[30]), .A1(A[30]) );
  inv01 U471 ( .Y(n427), .A(n438) );
  nor02 U472 ( .Y(n439), .A0(n419), .A1(n420) );
  inv01 U473 ( .Y(n429), .A(n439) );
  nor02 U474 ( .Y(n440), .A0(n422), .A1(n424) );
  inv01 U475 ( .Y(n430), .A(n440) );
  nor02 U476 ( .Y(n441), .A0(n426), .A1(n428) );
  inv01 U477 ( .Y(n431), .A(n441) );
  nor02 U478 ( .Y(n442), .A0(n432), .A1(n433) );
  inv01 U479 ( .Y(n435), .A(n442) );
  inv01 U480 ( .Y(SUM[29]), .A(n443) );
  inv02 U481 ( .Y(carry_30_), .A(n444) );
  inv02 U482 ( .Y(n445), .A(B[29]) );
  inv02 U483 ( .Y(n446), .A(A[29]) );
  inv02 U484 ( .Y(n447), .A(carry_29_) );
  nor02 U485 ( .Y(n448), .A0(n445), .A1(n449) );
  nor02 U486 ( .Y(n450), .A0(n446), .A1(n451) );
  nor02 U487 ( .Y(n452), .A0(n447), .A1(n453) );
  nor02 U488 ( .Y(n454), .A0(n447), .A1(n455) );
  nor02 U489 ( .Y(n443), .A0(n456), .A1(n457) );
  nor02 U490 ( .Y(n458), .A0(n446), .A1(n447) );
  nor02 U491 ( .Y(n459), .A0(n445), .A1(n447) );
  nor02 U492 ( .Y(n460), .A0(n445), .A1(n446) );
  nor02 U493 ( .Y(n444), .A0(n460), .A1(n461) );
  nor02 U494 ( .Y(n462), .A0(A[29]), .A1(carry_29_) );
  inv01 U495 ( .Y(n449), .A(n462) );
  nor02 U496 ( .Y(n463), .A0(B[29]), .A1(carry_29_) );
  inv01 U497 ( .Y(n451), .A(n463) );
  nor02 U498 ( .Y(n464), .A0(B[29]), .A1(A[29]) );
  inv01 U499 ( .Y(n453), .A(n464) );
  nor02 U500 ( .Y(n465), .A0(n445), .A1(n446) );
  inv01 U501 ( .Y(n455), .A(n465) );
  nor02 U502 ( .Y(n466), .A0(n448), .A1(n450) );
  inv01 U503 ( .Y(n456), .A(n466) );
  nor02 U504 ( .Y(n467), .A0(n452), .A1(n454) );
  inv01 U505 ( .Y(n457), .A(n467) );
  nor02 U506 ( .Y(n468), .A0(n458), .A1(n459) );
  inv01 U507 ( .Y(n461), .A(n468) );
  inv01 U508 ( .Y(SUM[28]), .A(n469) );
  inv02 U509 ( .Y(carry_29_), .A(n470) );
  inv02 U510 ( .Y(n471), .A(B[28]) );
  inv02 U511 ( .Y(n472), .A(A[28]) );
  inv02 U512 ( .Y(n473), .A(carry_28_) );
  nor02 U513 ( .Y(n474), .A0(n471), .A1(n475) );
  nor02 U514 ( .Y(n476), .A0(n472), .A1(n477) );
  nor02 U515 ( .Y(n478), .A0(n473), .A1(n479) );
  nor02 U516 ( .Y(n480), .A0(n473), .A1(n481) );
  nor02 U517 ( .Y(n469), .A0(n482), .A1(n483) );
  nor02 U518 ( .Y(n484), .A0(n472), .A1(n473) );
  nor02 U519 ( .Y(n485), .A0(n471), .A1(n473) );
  nor02 U520 ( .Y(n486), .A0(n471), .A1(n472) );
  nor02 U521 ( .Y(n470), .A0(n486), .A1(n487) );
  nor02 U522 ( .Y(n488), .A0(A[28]), .A1(carry_28_) );
  inv01 U523 ( .Y(n475), .A(n488) );
  nor02 U524 ( .Y(n489), .A0(B[28]), .A1(carry_28_) );
  inv01 U525 ( .Y(n477), .A(n489) );
  nor02 U526 ( .Y(n490), .A0(B[28]), .A1(A[28]) );
  inv01 U527 ( .Y(n479), .A(n490) );
  nor02 U528 ( .Y(n491), .A0(n471), .A1(n472) );
  inv01 U529 ( .Y(n481), .A(n491) );
  nor02 U530 ( .Y(n492), .A0(n474), .A1(n476) );
  inv01 U531 ( .Y(n482), .A(n492) );
  nor02 U532 ( .Y(n493), .A0(n478), .A1(n480) );
  inv01 U533 ( .Y(n483), .A(n493) );
  nor02 U534 ( .Y(n494), .A0(n484), .A1(n485) );
  inv01 U535 ( .Y(n487), .A(n494) );
  inv01 U536 ( .Y(SUM[27]), .A(n495) );
  inv02 U537 ( .Y(carry_28_), .A(n496) );
  inv02 U538 ( .Y(n497), .A(B[27]) );
  inv02 U539 ( .Y(n498), .A(A[27]) );
  inv02 U540 ( .Y(n499), .A(carry_27_) );
  nor02 U541 ( .Y(n500), .A0(n497), .A1(n501) );
  nor02 U542 ( .Y(n502), .A0(n498), .A1(n503) );
  nor02 U543 ( .Y(n504), .A0(n499), .A1(n505) );
  nor02 U544 ( .Y(n506), .A0(n499), .A1(n507) );
  nor02 U545 ( .Y(n495), .A0(n508), .A1(n509) );
  nor02 U546 ( .Y(n510), .A0(n498), .A1(n499) );
  nor02 U547 ( .Y(n511), .A0(n497), .A1(n499) );
  nor02 U548 ( .Y(n512), .A0(n497), .A1(n498) );
  nor02 U549 ( .Y(n496), .A0(n512), .A1(n513) );
  nor02 U550 ( .Y(n514), .A0(A[27]), .A1(carry_27_) );
  inv01 U551 ( .Y(n501), .A(n514) );
  nor02 U552 ( .Y(n515), .A0(B[27]), .A1(carry_27_) );
  inv01 U553 ( .Y(n503), .A(n515) );
  nor02 U554 ( .Y(n516), .A0(B[27]), .A1(A[27]) );
  inv01 U555 ( .Y(n505), .A(n516) );
  nor02 U556 ( .Y(n517), .A0(n497), .A1(n498) );
  inv01 U557 ( .Y(n507), .A(n517) );
  nor02 U558 ( .Y(n518), .A0(n500), .A1(n502) );
  inv01 U559 ( .Y(n508), .A(n518) );
  nor02 U560 ( .Y(n519), .A0(n504), .A1(n506) );
  inv01 U561 ( .Y(n509), .A(n519) );
  nor02 U562 ( .Y(n520), .A0(n510), .A1(n511) );
  inv01 U563 ( .Y(n513), .A(n520) );
  inv01 U564 ( .Y(SUM[26]), .A(n521) );
  inv02 U565 ( .Y(carry_27_), .A(n522) );
  inv02 U566 ( .Y(n523), .A(B[26]) );
  inv02 U567 ( .Y(n524), .A(A[26]) );
  inv02 U568 ( .Y(n525), .A(carry_26_) );
  nor02 U569 ( .Y(n526), .A0(n523), .A1(n527) );
  nor02 U570 ( .Y(n528), .A0(n524), .A1(n529) );
  nor02 U571 ( .Y(n530), .A0(n525), .A1(n531) );
  nor02 U572 ( .Y(n532), .A0(n525), .A1(n533) );
  nor02 U573 ( .Y(n521), .A0(n534), .A1(n535) );
  nor02 U574 ( .Y(n536), .A0(n524), .A1(n525) );
  nor02 U575 ( .Y(n537), .A0(n523), .A1(n525) );
  nor02 U576 ( .Y(n538), .A0(n523), .A1(n524) );
  nor02 U577 ( .Y(n522), .A0(n538), .A1(n539) );
  nor02 U578 ( .Y(n540), .A0(A[26]), .A1(carry_26_) );
  inv01 U579 ( .Y(n527), .A(n540) );
  nor02 U580 ( .Y(n541), .A0(B[26]), .A1(carry_26_) );
  inv01 U581 ( .Y(n529), .A(n541) );
  nor02 U582 ( .Y(n542), .A0(B[26]), .A1(A[26]) );
  inv01 U583 ( .Y(n531), .A(n542) );
  nor02 U584 ( .Y(n543), .A0(n523), .A1(n524) );
  inv01 U585 ( .Y(n533), .A(n543) );
  nor02 U586 ( .Y(n544), .A0(n526), .A1(n528) );
  inv01 U587 ( .Y(n534), .A(n544) );
  nor02 U588 ( .Y(n545), .A0(n530), .A1(n532) );
  inv01 U589 ( .Y(n535), .A(n545) );
  nor02 U590 ( .Y(n546), .A0(n536), .A1(n537) );
  inv01 U591 ( .Y(n539), .A(n546) );
  inv01 U592 ( .Y(SUM[25]), .A(n547) );
  inv02 U593 ( .Y(carry_26_), .A(n548) );
  inv02 U594 ( .Y(n549), .A(B[25]) );
  inv02 U595 ( .Y(n550), .A(A[25]) );
  inv02 U596 ( .Y(n551), .A(carry_25_) );
  nor02 U597 ( .Y(n552), .A0(n549), .A1(n553) );
  nor02 U598 ( .Y(n554), .A0(n550), .A1(n555) );
  nor02 U599 ( .Y(n556), .A0(n551), .A1(n557) );
  nor02 U600 ( .Y(n558), .A0(n551), .A1(n559) );
  nor02 U601 ( .Y(n547), .A0(n560), .A1(n561) );
  nor02 U602 ( .Y(n562), .A0(n550), .A1(n551) );
  nor02 U603 ( .Y(n563), .A0(n549), .A1(n551) );
  nor02 U604 ( .Y(n564), .A0(n549), .A1(n550) );
  nor02 U605 ( .Y(n548), .A0(n564), .A1(n565) );
  nor02 U606 ( .Y(n566), .A0(A[25]), .A1(carry_25_) );
  inv01 U607 ( .Y(n553), .A(n566) );
  nor02 U608 ( .Y(n567), .A0(B[25]), .A1(carry_25_) );
  inv01 U609 ( .Y(n555), .A(n567) );
  nor02 U610 ( .Y(n568), .A0(B[25]), .A1(A[25]) );
  inv01 U611 ( .Y(n557), .A(n568) );
  nor02 U612 ( .Y(n569), .A0(n549), .A1(n550) );
  inv01 U613 ( .Y(n559), .A(n569) );
  nor02 U614 ( .Y(n570), .A0(n552), .A1(n554) );
  inv01 U615 ( .Y(n560), .A(n570) );
  nor02 U616 ( .Y(n571), .A0(n556), .A1(n558) );
  inv01 U617 ( .Y(n561), .A(n571) );
  nor02 U618 ( .Y(n572), .A0(n562), .A1(n563) );
  inv01 U619 ( .Y(n565), .A(n572) );
  inv01 U620 ( .Y(SUM[24]), .A(n573) );
  inv02 U621 ( .Y(carry_25_), .A(n574) );
  inv02 U622 ( .Y(n575), .A(B[24]) );
  inv02 U623 ( .Y(n576), .A(A[24]) );
  inv02 U624 ( .Y(n577), .A(n599) );
  nor02 U625 ( .Y(n578), .A0(n575), .A1(n579) );
  nor02 U626 ( .Y(n580), .A0(n576), .A1(n581) );
  nor02 U627 ( .Y(n582), .A0(n577), .A1(n583) );
  nor02 U628 ( .Y(n584), .A0(n577), .A1(n585) );
  nor02 U629 ( .Y(n573), .A0(n586), .A1(n587) );
  nor02 U630 ( .Y(n588), .A0(n576), .A1(n577) );
  nor02 U631 ( .Y(n589), .A0(n575), .A1(n577) );
  nor02 U632 ( .Y(n590), .A0(n575), .A1(n576) );
  nor02 U633 ( .Y(n574), .A0(n590), .A1(n591) );
  nor02 U634 ( .Y(n592), .A0(A[24]), .A1(n599) );
  inv01 U635 ( .Y(n579), .A(n592) );
  nor02 U636 ( .Y(n593), .A0(B[24]), .A1(n599) );
  inv01 U637 ( .Y(n581), .A(n593) );
  nor02 U638 ( .Y(n594), .A0(B[24]), .A1(A[24]) );
  inv01 U639 ( .Y(n583), .A(n594) );
  nor02 U640 ( .Y(n595), .A0(n575), .A1(n576) );
  inv01 U641 ( .Y(n585), .A(n595) );
  nor02 U642 ( .Y(n596), .A0(n578), .A1(n580) );
  inv01 U643 ( .Y(n586), .A(n596) );
  nor02 U644 ( .Y(n597), .A0(n582), .A1(n584) );
  inv01 U645 ( .Y(n587), .A(n597) );
  nor02 U646 ( .Y(n598), .A0(n588), .A1(n589) );
  inv01 U647 ( .Y(n591), .A(n598) );
  buf02 U648 ( .Y(n599), .A(carry_24_) );
  buf02 U649 ( .Y(n600), .A(carry_23_) );
  buf02 U650 ( .Y(n601), .A(carry_22_) );
  buf02 U651 ( .Y(n602), .A(carry_21_) );
  buf02 U652 ( .Y(n603), .A(carry_20_) );
  buf02 U653 ( .Y(n604), .A(carry_19_) );
  buf02 U654 ( .Y(n605), .A(carry_18_) );
  buf02 U655 ( .Y(n606), .A(carry_17_) );
  buf02 U656 ( .Y(n607), .A(carry_16_) );
  buf02 U657 ( .Y(n608), .A(carry_15_) );
  buf02 U658 ( .Y(n609), .A(carry_14_) );
  buf02 U659 ( .Y(n610), .A(carry_13_) );
  buf02 U660 ( .Y(n611), .A(carry_12_) );
  buf02 U661 ( .Y(n612), .A(carry_11_) );
  buf02 U662 ( .Y(n613), .A(carry_10_) );
  buf02 U663 ( .Y(n614), .A(carry_9_) );
  buf02 U664 ( .Y(n615), .A(carry_8_) );
  buf02 U665 ( .Y(n616), .A(carry_7_) );
  buf02 U666 ( .Y(n617), .A(carry_6_) );
  buf02 U667 ( .Y(n618), .A(carry_5_) );
  buf02 U668 ( .Y(n619), .A(carry_4_) );
  buf02 U669 ( .Y(n620), .A(carry_3_) );
  buf02 U670 ( .Y(n621), .A(carry_2_) );
  xor2 U671 ( .Y(SUM[47]), .A0(B[47]), .A1(carry_47_) );
  xor2 U672 ( .Y(SUM[0]), .A0(B[0]), .A1(A[0]) );
  fadd1 U1_1 ( .S(SUM[1]), .CO(carry_2_), .A(A[1]), .B(B[1]), .CI(n26) );
  fadd1 U1_2 ( .S(SUM[2]), .CO(carry_3_), .A(A[2]), .B(B[2]), .CI(n621) );
  fadd1 U1_3 ( .S(SUM[3]), .CO(carry_4_), .A(A[3]), .B(B[3]), .CI(n620) );
  fadd1 U1_4 ( .S(SUM[4]), .CO(carry_5_), .A(A[4]), .B(B[4]), .CI(n619) );
  fadd1 U1_5 ( .S(SUM[5]), .CO(carry_6_), .A(A[5]), .B(B[5]), .CI(n618) );
  fadd1 U1_6 ( .S(SUM[6]), .CO(carry_7_), .A(A[6]), .B(B[6]), .CI(n617) );
  fadd1 U1_7 ( .S(SUM[7]), .CO(carry_8_), .A(A[7]), .B(B[7]), .CI(n616) );
  fadd1 U1_8 ( .S(SUM[8]), .CO(carry_9_), .A(A[8]), .B(B[8]), .CI(n615) );
  fadd1 U1_9 ( .S(SUM[9]), .CO(carry_10_), .A(A[9]), .B(B[9]), .CI(n614) );
  fadd1 U1_10 ( .S(SUM[10]), .CO(carry_11_), .A(A[10]), .B(B[10]), .CI(n613)
         );
  fadd1 U1_11 ( .S(SUM[11]), .CO(carry_12_), .A(A[11]), .B(B[11]), .CI(n612)
         );
  fadd1 U1_12 ( .S(SUM[12]), .CO(carry_13_), .A(A[12]), .B(B[12]), .CI(n611)
         );
  fadd1 U1_13 ( .S(SUM[13]), .CO(carry_14_), .A(A[13]), .B(B[13]), .CI(n610)
         );
  fadd1 U1_14 ( .S(SUM[14]), .CO(carry_15_), .A(A[14]), .B(B[14]), .CI(n609)
         );
  fadd1 U1_15 ( .S(SUM[15]), .CO(carry_16_), .A(A[15]), .B(B[15]), .CI(n608)
         );
  fadd1 U1_16 ( .S(SUM[16]), .CO(carry_17_), .A(A[16]), .B(B[16]), .CI(n607)
         );
  fadd1 U1_17 ( .S(SUM[17]), .CO(carry_18_), .A(A[17]), .B(B[17]), .CI(n606)
         );
  fadd1 U1_18 ( .S(SUM[18]), .CO(carry_19_), .A(A[18]), .B(B[18]), .CI(n605)
         );
  fadd1 U1_19 ( .S(SUM[19]), .CO(carry_20_), .A(A[19]), .B(B[19]), .CI(n604)
         );
  fadd1 U1_20 ( .S(SUM[20]), .CO(carry_21_), .A(A[20]), .B(B[20]), .CI(n603)
         );
  fadd1 U1_21 ( .S(SUM[21]), .CO(carry_22_), .A(A[21]), .B(B[21]), .CI(n602)
         );
  fadd1 U1_22 ( .S(SUM[22]), .CO(carry_23_), .A(A[22]), .B(B[22]), .CI(n601)
         );
  fadd1 U1_23 ( .S(SUM[23]), .CO(carry_24_), .A(A[23]), .B(B[23]), .CI(n600)
         );
endmodule


module serial_mul_DW01_inc_5_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   carry_4_, carry_3_, carry_2_;

  inv01 U5 ( .Y(SUM[0]), .A(A[0]) );
  xor2 U6 ( .Y(SUM[4]), .A0(carry_4_), .A1(A[4]) );
  hadd1 U1_1_1 ( .S(SUM[1]), .CO(carry_2_), .A(A[1]), .B(A[0]) );
  hadd1 U1_1_2 ( .S(SUM[2]), .CO(carry_3_), .A(A[2]), .B(carry_2_) );
  hadd1 U1_1_3 ( .S(SUM[3]), .CO(carry_4_), .A(A[3]), .B(carry_3_) );
endmodule


module serial_mul ( clk_i, fracta_i, fractb_i, signa_i, signb_i, start_i, 
        fract_o, sign_o, ready_o );
  input [23:0] fracta_i;
  input [23:0] fractb_i;
  output [47:0] fract_o;
  input clk_i, signa_i, signb_i, start_i;
  output sign_o, ready_o;
  wire   s_sign_o, s_ready_o, s_fracta_i_23_, s_fracta_i_0_, s_fractb_i_21_,
         s_fractb_i_20_, s_fractb_i_19_, s_fractb_i_18_, s_fractb_i_13_,
         s_fractb_i_12_, s_fractb_i_11_, s_fractb_i_10_, s_fractb_i_5_,
         s_fractb_i_3_, v_prod_shl239_38_, v_prod_shl239_37_,
         v_prod_shl239_36_, v_prod_shl239_35_, v_prod_shl239_34_,
         v_prod_shl239_33_, v_prod_shl239_32_, v_prod_shl239_31_,
         v_prod_shl239_30_, v_prod_shl239_29_, v_prod_shl239_28_,
         v_prod_shl239_27_, v_prod_shl239_26_, v_prod_shl239_25_,
         v_prod_shl239_24_, v_prod_shl239_23_, v_prod_shl239_22_,
         v_prod_shl239_21_, v_prod_shl239_20_, v_prod_shl239_19_,
         v_prod_shl239_18_, v_prod_shl239_17_, v_prod_shl239_16_,
         v_prod_shl239_15_, v_prod_shl239_14_, v_prod_shl239_13_,
         v_prod_shl239_12_, v_prod_shl239_11_, v_prod_shl239_7_,
         v_prod_shl239_0_, s_state132, sum218_4_, sum218_3_, sum218_2_,
         sum218_1_, sum218_0_, n313_0_, n____return527_47_, n____return527_46_,
         n____return527_45_, n____return527_44_, n____return527_43_,
         n____return527_42_, n____return527_41_, n____return527_40_,
         n____return527_39_, n____return527_38_, n____return527_37_,
         n____return527_36_, n____return527_35_, n____return527_34_,
         n____return527_33_, n____return527_32_, n____return527_31_,
         n____return527_30_, n____return527_29_, n____return527_28_,
         n____return527_27_, n____return527_26_, n____return527_25_,
         n____return527_24_, n____return527_23_, n____return527_22_,
         n____return527_21_, n____return527_20_, n____return527_19_,
         n____return527_18_, n____return527_17_, n____return527_16_,
         n____return527_15_, n____return527_14_, n____return527_13_,
         n____return527_12_, n____return527_11_, n____return527_10_,
         n____return527_9_, n____return527_8_, n____return527_7_,
         n____return527_6_, n____return527_5_, n____return527_4_,
         n____return527_3_, n____return527_2_, n____return527_1_,
         n____return527_0_, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056;
  wire   [47:0] s_fract_o;
  wire   [4:0] s_count;

  dff s_count_reg_0_ ( .Q(s_count[0]), .QB(n1753), .D(n985), .CLK(clk_i) );
  dff s_count_reg_1_ ( .Q(s_count[1]), .D(n986), .CLK(clk_i) );
  dff s_count_reg_2_ ( .Q(s_count[2]), .QB(n1361), .D(n987), .CLK(clk_i) );
  dff s_count_reg_3_ ( .Q(s_count[3]), .QB(n1892), .D(n988), .CLK(clk_i) );
  dff s_count_reg_4_ ( .Q(s_count[4]), .D(n989), .CLK(clk_i) );
  dff s_fract_o_reg_47_ ( .Q(s_fract_o[47]), .D(n990), .CLK(clk_i) );
  dff s_fract_o_reg_46_ ( .Q(s_fract_o[46]), .D(n991), .CLK(clk_i) );
  dff s_fract_o_reg_45_ ( .Q(s_fract_o[45]), .D(n992), .CLK(clk_i) );
  dff s_fract_o_reg_44_ ( .Q(s_fract_o[44]), .D(n993), .CLK(clk_i) );
  dff s_fract_o_reg_43_ ( .Q(s_fract_o[43]), .D(n994), .CLK(clk_i) );
  dff s_fract_o_reg_42_ ( .Q(s_fract_o[42]), .D(n995), .CLK(clk_i) );
  dff s_fract_o_reg_41_ ( .Q(s_fract_o[41]), .D(n996), .CLK(clk_i) );
  dff s_fract_o_reg_40_ ( .Q(s_fract_o[40]), .D(n997), .CLK(clk_i) );
  dff s_fract_o_reg_39_ ( .Q(s_fract_o[39]), .D(n998), .CLK(clk_i) );
  dff s_fract_o_reg_38_ ( .Q(s_fract_o[38]), .D(n999), .CLK(clk_i) );
  dff s_fract_o_reg_37_ ( .Q(s_fract_o[37]), .D(n1000), .CLK(clk_i) );
  dff s_fract_o_reg_36_ ( .Q(s_fract_o[36]), .D(n1001), .CLK(clk_i) );
  dff s_fract_o_reg_35_ ( .Q(s_fract_o[35]), .D(n1002), .CLK(clk_i) );
  dff s_fract_o_reg_34_ ( .Q(s_fract_o[34]), .D(n1003), .CLK(clk_i) );
  dff s_fract_o_reg_33_ ( .Q(s_fract_o[33]), .D(n1004), .CLK(clk_i) );
  dff s_fract_o_reg_32_ ( .Q(s_fract_o[32]), .D(n1005), .CLK(clk_i) );
  dff s_fract_o_reg_31_ ( .Q(s_fract_o[31]), .D(n1006), .CLK(clk_i) );
  dff s_fract_o_reg_30_ ( .Q(s_fract_o[30]), .D(n1007), .CLK(clk_i) );
  dff s_fract_o_reg_29_ ( .Q(s_fract_o[29]), .D(n1008), .CLK(clk_i) );
  dff s_fract_o_reg_28_ ( .Q(s_fract_o[28]), .D(n1009), .CLK(clk_i) );
  dff s_fract_o_reg_27_ ( .Q(s_fract_o[27]), .D(n1010), .CLK(clk_i) );
  dff s_fract_o_reg_26_ ( .Q(s_fract_o[26]), .D(n1011), .CLK(clk_i) );
  dff s_fract_o_reg_25_ ( .Q(s_fract_o[25]), .D(n1012), .CLK(clk_i) );
  dff s_fract_o_reg_24_ ( .Q(s_fract_o[24]), .D(n1013), .CLK(clk_i) );
  dff s_fract_o_reg_23_ ( .Q(s_fract_o[23]), .QB(n2040), .D(n1014), .CLK(clk_i) );
  dff s_fract_o_reg_22_ ( .Q(s_fract_o[22]), .QB(n2041), .D(n1015), .CLK(clk_i) );
  dff s_fract_o_reg_21_ ( .Q(s_fract_o[21]), .QB(n2042), .D(n1016), .CLK(clk_i) );
  dff s_fract_o_reg_20_ ( .Q(s_fract_o[20]), .QB(n2043), .D(n1017), .CLK(clk_i) );
  dff s_fract_o_reg_19_ ( .Q(s_fract_o[19]), .QB(n2045), .D(n1018), .CLK(clk_i) );
  dff s_fract_o_reg_18_ ( .Q(s_fract_o[18]), .QB(n2046), .D(n1019), .CLK(clk_i) );
  dff s_fract_o_reg_17_ ( .Q(s_fract_o[17]), .QB(n2047), .D(n1020), .CLK(clk_i) );
  dff s_fract_o_reg_16_ ( .Q(s_fract_o[16]), .QB(n2048), .D(n1021), .CLK(clk_i) );
  dff s_fract_o_reg_15_ ( .Q(s_fract_o[15]), .QB(n2049), .D(n1022), .CLK(clk_i) );
  dff s_fract_o_reg_14_ ( .Q(s_fract_o[14]), .QB(n2050), .D(n1023), .CLK(clk_i) );
  dff s_fract_o_reg_13_ ( .Q(s_fract_o[13]), .QB(n2051), .D(n1024), .CLK(clk_i) );
  dff s_fract_o_reg_12_ ( .Q(s_fract_o[12]), .QB(n2052), .D(n1025), .CLK(clk_i) );
  dff s_fract_o_reg_11_ ( .Q(s_fract_o[11]), .QB(n2053), .D(n1026), .CLK(clk_i) );
  dff s_fract_o_reg_10_ ( .Q(s_fract_o[10]), .QB(n2054), .D(n1027), .CLK(clk_i) );
  dff s_fract_o_reg_9_ ( .Q(s_fract_o[9]), .QB(n2032), .D(n1028), .CLK(clk_i)
         );
  dff s_fract_o_reg_8_ ( .Q(s_fract_o[8]), .QB(n2033), .D(n1029), .CLK(clk_i)
         );
  dff s_fract_o_reg_7_ ( .Q(s_fract_o[7]), .QB(n2034), .D(n1030), .CLK(clk_i)
         );
  dff s_fract_o_reg_6_ ( .Q(s_fract_o[6]), .QB(n2035), .D(n1031), .CLK(clk_i)
         );
  dff s_fract_o_reg_5_ ( .Q(s_fract_o[5]), .QB(n2036), .D(n1032), .CLK(clk_i)
         );
  dff s_fract_o_reg_4_ ( .Q(s_fract_o[4]), .QB(n2037), .D(n1033), .CLK(clk_i)
         );
  dff s_fract_o_reg_3_ ( .Q(s_fract_o[3]), .QB(n2038), .D(n1034), .CLK(clk_i)
         );
  dff s_fract_o_reg_2_ ( .Q(s_fract_o[2]), .QB(n2039), .D(n1035), .CLK(clk_i)
         );
  dff s_fract_o_reg_1_ ( .Q(s_fract_o[1]), .QB(n2044), .D(n1036), .CLK(clk_i)
         );
  dff s_fract_o_reg_0_ ( .Q(s_fract_o[0]), .QB(n2055), .D(n1037), .CLK(clk_i)
         );
  dff s_state_reg ( .Q(n313_0_), .D(n1038), .CLK(clk_i) );
  dff s_ready_o_reg ( .Q(s_ready_o), .QB(n2031), .D(n1039), .CLK(clk_i) );
  dff s_fracta_i_reg_23_ ( .Q(s_fracta_i_23_), .D(fracta_i[23]), .CLK(clk_i)
         );
  dff s_fracta_i_reg_22_ ( .Q(n724), .D(fracta_i[22]), .CLK(clk_i) );
  dff s_fracta_i_reg_21_ ( .Q(n723), .D(fracta_i[21]), .CLK(clk_i) );
  dff s_fracta_i_reg_20_ ( .Q(n722), .D(fracta_i[20]), .CLK(clk_i) );
  dff s_fracta_i_reg_19_ ( .Q(n721), .D(fracta_i[19]), .CLK(clk_i) );
  dff s_fracta_i_reg_18_ ( .Q(n720), .D(fracta_i[18]), .CLK(clk_i) );
  dff s_fracta_i_reg_17_ ( .Q(n719), .D(fracta_i[17]), .CLK(clk_i) );
  dff s_fracta_i_reg_16_ ( .Q(n718), .D(fracta_i[16]), .CLK(clk_i) );
  dff s_fracta_i_reg_15_ ( .Q(n717), .D(fracta_i[15]), .CLK(clk_i) );
  dff s_fracta_i_reg_14_ ( .Q(n716), .D(fracta_i[14]), .CLK(clk_i) );
  dff s_fracta_i_reg_13_ ( .Q(n715), .D(fracta_i[13]), .CLK(clk_i) );
  dff s_fracta_i_reg_12_ ( .Q(n714), .D(fracta_i[12]), .CLK(clk_i) );
  dff s_fracta_i_reg_11_ ( .Q(n713), .D(fracta_i[11]), .CLK(clk_i) );
  dff s_fracta_i_reg_10_ ( .Q(n712), .D(fracta_i[10]), .CLK(clk_i) );
  dff s_fracta_i_reg_9_ ( .Q(n711), .D(fracta_i[9]), .CLK(clk_i) );
  dff s_fracta_i_reg_8_ ( .Q(n710), .D(fracta_i[8]), .CLK(clk_i) );
  dff s_fracta_i_reg_7_ ( .Q(n709), .D(fracta_i[7]), .CLK(clk_i) );
  dff s_fracta_i_reg_6_ ( .Q(n708), .D(fracta_i[6]), .CLK(clk_i) );
  dff s_fracta_i_reg_5_ ( .Q(n707), .D(fracta_i[5]), .CLK(clk_i) );
  dff s_fracta_i_reg_4_ ( .Q(n706), .D(fracta_i[4]), .CLK(clk_i) );
  dff s_fracta_i_reg_3_ ( .Q(n705), .D(fracta_i[3]), .CLK(clk_i) );
  dff s_fracta_i_reg_2_ ( .Q(n704), .D(fracta_i[2]), .CLK(clk_i) );
  dff s_fracta_i_reg_1_ ( .Q(n703), .D(fracta_i[1]), .CLK(clk_i) );
  dff s_fracta_i_reg_0_ ( .Q(s_fracta_i_0_), .D(fracta_i[0]), .CLK(clk_i) );
  dff s_fractb_i_reg_23_ ( .QB(n702), .D(fractb_i[23]), .CLK(clk_i) );
  dff s_fractb_i_reg_22_ ( .QB(n701), .D(fractb_i[22]), .CLK(clk_i) );
  dff s_fractb_i_reg_21_ ( .Q(s_fractb_i_21_), .D(fractb_i[21]), .CLK(clk_i)
         );
  dff s_fractb_i_reg_20_ ( .Q(s_fractb_i_20_), .D(fractb_i[20]), .CLK(clk_i)
         );
  dff s_fractb_i_reg_19_ ( .Q(s_fractb_i_19_), .D(fractb_i[19]), .CLK(clk_i)
         );
  dff s_fractb_i_reg_18_ ( .Q(s_fractb_i_18_), .D(fractb_i[18]), .CLK(clk_i)
         );
  dff s_fractb_i_reg_17_ ( .QB(n700), .D(fractb_i[17]), .CLK(clk_i) );
  dff s_fractb_i_reg_16_ ( .QB(n699), .D(fractb_i[16]), .CLK(clk_i) );
  dff s_fractb_i_reg_15_ ( .QB(n698), .D(fractb_i[15]), .CLK(clk_i) );
  dff s_fractb_i_reg_14_ ( .QB(n697), .D(fractb_i[14]), .CLK(clk_i) );
  dff s_fractb_i_reg_13_ ( .Q(s_fractb_i_13_), .D(fractb_i[13]), .CLK(clk_i)
         );
  dff s_fractb_i_reg_12_ ( .Q(s_fractb_i_12_), .D(fractb_i[12]), .CLK(clk_i)
         );
  dff s_fractb_i_reg_11_ ( .Q(s_fractb_i_11_), .D(fractb_i[11]), .CLK(clk_i)
         );
  dff s_fractb_i_reg_10_ ( .Q(s_fractb_i_10_), .D(fractb_i[10]), .CLK(clk_i)
         );
  dff s_fractb_i_reg_9_ ( .QB(n696), .D(fractb_i[9]), .CLK(clk_i) );
  dff s_fractb_i_reg_8_ ( .QB(n695), .D(fractb_i[8]), .CLK(clk_i) );
  dff s_fractb_i_reg_7_ ( .QB(n694), .D(fractb_i[7]), .CLK(clk_i) );
  dff s_fractb_i_reg_6_ ( .QB(n693), .D(fractb_i[6]), .CLK(clk_i) );
  dff s_fractb_i_reg_5_ ( .Q(s_fractb_i_5_), .D(fractb_i[5]), .CLK(clk_i) );
  dff s_fractb_i_reg_4_ ( .QB(n692), .D(fractb_i[4]), .CLK(clk_i) );
  dff s_fractb_i_reg_3_ ( .Q(s_fractb_i_3_), .D(fractb_i[3]), .CLK(clk_i) );
  dff s_fractb_i_reg_2_ ( .QB(n691), .D(fractb_i[2]), .CLK(clk_i) );
  dff s_fractb_i_reg_1_ ( .QB(n690), .D(fractb_i[1]), .CLK(clk_i) );
  dff s_fractb_i_reg_0_ ( .Q(n2056), .D(fractb_i[0]), .CLK(clk_i) );
  dff fract_o_reg_47_ ( .Q(fract_o[47]), .D(s_fract_o[47]), .CLK(clk_i) );
  dff fract_o_reg_46_ ( .Q(fract_o[46]), .D(s_fract_o[46]), .CLK(clk_i) );
  dff fract_o_reg_45_ ( .Q(fract_o[45]), .D(s_fract_o[45]), .CLK(clk_i) );
  dff fract_o_reg_44_ ( .Q(fract_o[44]), .D(s_fract_o[44]), .CLK(clk_i) );
  dff fract_o_reg_43_ ( .Q(fract_o[43]), .D(s_fract_o[43]), .CLK(clk_i) );
  dff fract_o_reg_42_ ( .Q(fract_o[42]), .D(s_fract_o[42]), .CLK(clk_i) );
  dff fract_o_reg_41_ ( .Q(fract_o[41]), .D(s_fract_o[41]), .CLK(clk_i) );
  dff fract_o_reg_40_ ( .Q(fract_o[40]), .D(s_fract_o[40]), .CLK(clk_i) );
  dff fract_o_reg_39_ ( .Q(fract_o[39]), .D(s_fract_o[39]), .CLK(clk_i) );
  dff fract_o_reg_38_ ( .Q(fract_o[38]), .D(s_fract_o[38]), .CLK(clk_i) );
  dff fract_o_reg_37_ ( .Q(fract_o[37]), .D(s_fract_o[37]), .CLK(clk_i) );
  dff fract_o_reg_36_ ( .Q(fract_o[36]), .D(s_fract_o[36]), .CLK(clk_i) );
  dff fract_o_reg_35_ ( .Q(fract_o[35]), .D(s_fract_o[35]), .CLK(clk_i) );
  dff fract_o_reg_34_ ( .Q(fract_o[34]), .D(s_fract_o[34]), .CLK(clk_i) );
  dff fract_o_reg_33_ ( .Q(fract_o[33]), .D(s_fract_o[33]), .CLK(clk_i) );
  dff fract_o_reg_32_ ( .Q(fract_o[32]), .D(s_fract_o[32]), .CLK(clk_i) );
  dff fract_o_reg_31_ ( .Q(fract_o[31]), .D(s_fract_o[31]), .CLK(clk_i) );
  dff fract_o_reg_30_ ( .Q(fract_o[30]), .D(s_fract_o[30]), .CLK(clk_i) );
  dff fract_o_reg_29_ ( .Q(fract_o[29]), .D(s_fract_o[29]), .CLK(clk_i) );
  dff fract_o_reg_28_ ( .Q(fract_o[28]), .D(s_fract_o[28]), .CLK(clk_i) );
  dff fract_o_reg_27_ ( .Q(fract_o[27]), .D(s_fract_o[27]), .CLK(clk_i) );
  dff fract_o_reg_26_ ( .Q(fract_o[26]), .D(s_fract_o[26]), .CLK(clk_i) );
  dff fract_o_reg_25_ ( .Q(fract_o[25]), .D(s_fract_o[25]), .CLK(clk_i) );
  dff fract_o_reg_24_ ( .Q(fract_o[24]), .D(s_fract_o[24]), .CLK(clk_i) );
  dff fract_o_reg_23_ ( .Q(fract_o[23]), .D(s_fract_o[23]), .CLK(clk_i) );
  dff fract_o_reg_22_ ( .Q(fract_o[22]), .D(s_fract_o[22]), .CLK(clk_i) );
  dff fract_o_reg_21_ ( .Q(fract_o[21]), .D(s_fract_o[21]), .CLK(clk_i) );
  dff fract_o_reg_20_ ( .Q(fract_o[20]), .D(s_fract_o[20]), .CLK(clk_i) );
  dff fract_o_reg_19_ ( .Q(fract_o[19]), .D(s_fract_o[19]), .CLK(clk_i) );
  dff fract_o_reg_18_ ( .Q(fract_o[18]), .D(s_fract_o[18]), .CLK(clk_i) );
  dff fract_o_reg_17_ ( .Q(fract_o[17]), .D(s_fract_o[17]), .CLK(clk_i) );
  dff fract_o_reg_16_ ( .Q(fract_o[16]), .D(s_fract_o[16]), .CLK(clk_i) );
  dff fract_o_reg_15_ ( .Q(fract_o[15]), .D(s_fract_o[15]), .CLK(clk_i) );
  dff fract_o_reg_14_ ( .Q(fract_o[14]), .D(s_fract_o[14]), .CLK(clk_i) );
  dff fract_o_reg_13_ ( .Q(fract_o[13]), .D(s_fract_o[13]), .CLK(clk_i) );
  dff fract_o_reg_12_ ( .Q(fract_o[12]), .D(s_fract_o[12]), .CLK(clk_i) );
  dff fract_o_reg_11_ ( .Q(fract_o[11]), .D(s_fract_o[11]), .CLK(clk_i) );
  dff fract_o_reg_10_ ( .Q(fract_o[10]), .D(s_fract_o[10]), .CLK(clk_i) );
  dff fract_o_reg_9_ ( .Q(fract_o[9]), .D(s_fract_o[9]), .CLK(clk_i) );
  dff fract_o_reg_8_ ( .Q(fract_o[8]), .D(s_fract_o[8]), .CLK(clk_i) );
  dff fract_o_reg_7_ ( .Q(fract_o[7]), .D(s_fract_o[7]), .CLK(clk_i) );
  dff fract_o_reg_6_ ( .Q(fract_o[6]), .D(s_fract_o[6]), .CLK(clk_i) );
  dff fract_o_reg_5_ ( .Q(fract_o[5]), .D(s_fract_o[5]), .CLK(clk_i) );
  dff fract_o_reg_4_ ( .Q(fract_o[4]), .D(s_fract_o[4]), .CLK(clk_i) );
  dff fract_o_reg_3_ ( .Q(fract_o[3]), .D(s_fract_o[3]), .CLK(clk_i) );
  dff fract_o_reg_2_ ( .Q(fract_o[2]), .D(s_fract_o[2]), .CLK(clk_i) );
  dff fract_o_reg_1_ ( .Q(fract_o[1]), .D(s_fract_o[1]), .CLK(clk_i) );
  dff fract_o_reg_0_ ( .Q(fract_o[0]), .D(s_fract_o[0]), .CLK(clk_i) );
  dff s_start_i_reg ( .Q(s_state132), .D(start_i), .CLK(clk_i) );
  dff sign_o_reg ( .Q(sign_o), .D(s_sign_o), .CLK(clk_i) );
  dff ready_o_reg ( .Q(ready_o), .D(s_ready_o), .CLK(clk_i) );
  ao22 U511 ( .Y(n1041), .A0(n1903), .A1(n719), .B0(n1909), .B1(n720) );
  inv01 U512 ( .Y(n1042), .A(n1041) );
  ao22 U513 ( .Y(n1043), .A0(n1903), .A1(n715), .B0(n1909), .B1(n716) );
  inv01 U514 ( .Y(n1044), .A(n1043) );
  ao22 U515 ( .Y(n1045), .A0(n1903), .A1(n724), .B0(n1907), .B1(s_fracta_i_23_) );
  inv01 U516 ( .Y(n1046), .A(n1045) );
  inv01 U517 ( .Y(n1999), .A(n1047) );
  nor02 U518 ( .Y(n1048), .A0(n1868), .A1(n1898) );
  nor02 U519 ( .Y(n1049), .A0(n1854), .A1(n1983) );
  nor02 U520 ( .Y(n1047), .A0(n1048), .A1(n1049) );
  inv01 U521 ( .Y(n1868), .A(n1867) );
  inv01 U522 ( .Y(n1050), .A(n2018) );
  buf02 U523 ( .Y(n1051), .A(n2005) );
  buf02 U524 ( .Y(n1052), .A(n1977) );
  buf02 U525 ( .Y(n1053), .A(v_prod_shl239_15_) );
  buf02 U526 ( .Y(n1054), .A(n2010) );
  ao22 U527 ( .Y(n1055), .A0(n1903), .A1(s_fracta_i_0_), .B0(n1908), .B1(n703)
         );
  inv01 U528 ( .Y(n1056), .A(n1055) );
  nand02 U529 ( .Y(n1963), .A0(n1057), .A1(n1058) );
  inv01 U530 ( .Y(n1059), .A(n1916) );
  inv01 U531 ( .Y(n1060), .A(n1902) );
  inv01 U532 ( .Y(n1061), .A(n1729) );
  inv01 U533 ( .Y(n1062), .A(n____return527_2_) );
  nand02 U534 ( .Y(n1063), .A0(n1059), .A1(n1060) );
  nand02 U535 ( .Y(n1064), .A0(n1059), .A1(n1061) );
  nand02 U536 ( .Y(n1065), .A0(n1060), .A1(n1062) );
  nand02 U537 ( .Y(n1066), .A0(n1061), .A1(n1062) );
  nand02 U538 ( .Y(n1067), .A0(n1063), .A1(n1064) );
  inv01 U539 ( .Y(n1057), .A(n1067) );
  nand02 U540 ( .Y(n1068), .A0(n1065), .A1(n1066) );
  inv01 U541 ( .Y(n1058), .A(n1068) );
  nand02 U542 ( .Y(n1965), .A0(n1069), .A1(n1070) );
  inv01 U543 ( .Y(n1071), .A(n1916) );
  inv01 U544 ( .Y(n1072), .A(n1902) );
  inv01 U545 ( .Y(n1073), .A(n1744) );
  inv01 U546 ( .Y(n1074), .A(n____return527_4_) );
  nand02 U547 ( .Y(n1075), .A0(n1071), .A1(n1072) );
  nand02 U548 ( .Y(n1076), .A0(n1071), .A1(n1073) );
  nand02 U549 ( .Y(n1077), .A0(n1072), .A1(n1074) );
  nand02 U550 ( .Y(n1078), .A0(n1073), .A1(n1074) );
  nand02 U551 ( .Y(n1079), .A0(n1075), .A1(n1076) );
  inv01 U552 ( .Y(n1069), .A(n1079) );
  nand02 U553 ( .Y(n1080), .A0(n1077), .A1(n1078) );
  inv01 U554 ( .Y(n1070), .A(n1080) );
  nand02 U555 ( .Y(n1976), .A0(n1081), .A1(n1082) );
  inv01 U556 ( .Y(n1083), .A(n1916) );
  inv01 U557 ( .Y(n1084), .A(n1902) );
  inv01 U558 ( .Y(n1085), .A(n1640) );
  inv01 U559 ( .Y(n1086), .A(n____return527_10_) );
  nand02 U560 ( .Y(n1087), .A0(n1083), .A1(n1084) );
  nand02 U561 ( .Y(n1088), .A0(n1083), .A1(n1085) );
  nand02 U562 ( .Y(n1089), .A0(n1084), .A1(n1086) );
  nand02 U563 ( .Y(n1090), .A0(n1085), .A1(n1086) );
  nand02 U564 ( .Y(n1091), .A0(n1087), .A1(n1088) );
  inv01 U565 ( .Y(n1081), .A(n1091) );
  nand02 U566 ( .Y(n1092), .A0(n1089), .A1(n1090) );
  inv01 U567 ( .Y(n1082), .A(n1092) );
  ao22 U568 ( .Y(n1093), .A0(n1738), .A1(n1902), .B0(n____return527_3_), .B1(
        n1916) );
  inv01 U569 ( .Y(n1094), .A(n1093) );
  inv02 U570 ( .Y(n1640), .A(n1639) );
  nand02 U571 ( .Y(n1969), .A0(n1095), .A1(n1096) );
  inv01 U572 ( .Y(n1097), .A(n1916) );
  inv01 U573 ( .Y(n1098), .A(n1902) );
  inv01 U574 ( .Y(n1099), .A(n1741) );
  inv01 U575 ( .Y(n1100), .A(n____return527_6_) );
  nand02 U576 ( .Y(n1101), .A0(n1097), .A1(n1098) );
  nand02 U577 ( .Y(n1102), .A0(n1097), .A1(n1099) );
  nand02 U578 ( .Y(n1103), .A0(n1098), .A1(n1100) );
  nand02 U579 ( .Y(n1104), .A0(n1099), .A1(n1100) );
  nand02 U580 ( .Y(n1105), .A0(n1101), .A1(n1102) );
  inv01 U581 ( .Y(n1095), .A(n1105) );
  nand02 U582 ( .Y(n1106), .A0(n1103), .A1(n1104) );
  inv01 U583 ( .Y(n1096), .A(n1106) );
  nand02 U584 ( .Y(n1971), .A0(n1107), .A1(n1108) );
  inv01 U585 ( .Y(n1109), .A(n1916) );
  inv01 U586 ( .Y(n1110), .A(n1902) );
  inv01 U587 ( .Y(n1111), .A(v_prod_shl239_7_) );
  inv01 U588 ( .Y(n1112), .A(n____return527_7_) );
  nand02 U589 ( .Y(n1113), .A0(n1109), .A1(n1110) );
  nand02 U590 ( .Y(n1114), .A0(n1109), .A1(n1111) );
  nand02 U591 ( .Y(n1115), .A0(n1110), .A1(n1112) );
  nand02 U592 ( .Y(n1116), .A0(n1111), .A1(n1112) );
  nand02 U593 ( .Y(n1117), .A0(n1113), .A1(n1114) );
  inv01 U594 ( .Y(n1107), .A(n1117) );
  nand02 U595 ( .Y(n1118), .A0(n1115), .A1(n1116) );
  inv01 U596 ( .Y(n1108), .A(n1118) );
  nand02 U597 ( .Y(n1967), .A0(n1119), .A1(n1120) );
  inv01 U598 ( .Y(n1121), .A(n1916) );
  inv01 U599 ( .Y(n1122), .A(n1902) );
  inv01 U600 ( .Y(n1123), .A(n1747) );
  inv01 U601 ( .Y(n1124), .A(n____return527_5_) );
  nand02 U602 ( .Y(n1125), .A0(n1121), .A1(n1122) );
  nand02 U603 ( .Y(n1126), .A0(n1121), .A1(n1123) );
  nand02 U604 ( .Y(n1127), .A0(n1122), .A1(n1124) );
  nand02 U605 ( .Y(n1128), .A0(n1123), .A1(n1124) );
  nand02 U606 ( .Y(n1129), .A0(n1125), .A1(n1126) );
  inv01 U607 ( .Y(n1119), .A(n1129) );
  nand02 U608 ( .Y(n1130), .A0(n1127), .A1(n1128) );
  inv01 U609 ( .Y(n1120), .A(n1130) );
  ao22 U610 ( .Y(n1131), .A0(n1735), .A1(n1902), .B0(n____return527_8_), .B1(
        n1916) );
  inv01 U611 ( .Y(n1132), .A(n1131) );
  ao22 U612 ( .Y(n1133), .A0(n1901), .A1(n1943), .B0(n1897), .B1(n1946) );
  inv01 U613 ( .Y(n1134), .A(n1133) );
  nand02 U614 ( .Y(n1975), .A0(n1135), .A1(n1136) );
  inv01 U615 ( .Y(n1137), .A(n1916) );
  inv01 U616 ( .Y(n1138), .A(n1902) );
  inv01 U617 ( .Y(n1139), .A(n1638) );
  inv01 U618 ( .Y(n1140), .A(n____return527_9_) );
  nand02 U619 ( .Y(n1141), .A0(n1137), .A1(n1138) );
  nand02 U620 ( .Y(n1142), .A0(n1137), .A1(n1139) );
  nand02 U621 ( .Y(n1143), .A0(n1138), .A1(n1140) );
  nand02 U622 ( .Y(n1144), .A0(n1139), .A1(n1140) );
  nand02 U623 ( .Y(n1145), .A0(n1141), .A1(n1142) );
  inv01 U624 ( .Y(n1135), .A(n1145) );
  nand02 U625 ( .Y(n1146), .A0(n1143), .A1(n1144) );
  inv01 U626 ( .Y(n1136), .A(n1146) );
  ao22 U627 ( .Y(n1147), .A0(n1732), .A1(n1902), .B0(n____return527_1_), .B1(
        n1916) );
  inv01 U628 ( .Y(n1148), .A(n1147) );
  inv02 U629 ( .Y(n1638), .A(n1637) );
  ao22 U630 ( .Y(n1149), .A0(n1897), .A1(n1943), .B0(n1904), .B1(n1985) );
  inv01 U631 ( .Y(n1150), .A(n1149) );
  buf02 U632 ( .Y(n1151), .A(n2008) );
  ao22 U633 ( .Y(n1152), .A0(n1758), .A1(n1365), .B0(n1862), .B1(n1951) );
  inv01 U634 ( .Y(n1153), .A(n1152) );
  ao22 U635 ( .Y(n1154), .A0(n1902), .A1(n1652), .B0(n____return527_15_), .B1(
        n1916) );
  inv01 U636 ( .Y(n1155), .A(n1154) );
  ao22 U637 ( .Y(n1156), .A0(n1252), .A1(n1759), .B0(n1860), .B1(n1892) );
  inv01 U638 ( .Y(n1157), .A(n1156) );
  ao22 U639 ( .Y(n1158), .A0(n1964), .A1(n1762), .B0(n1942), .B1(n1539) );
  inv01 U640 ( .Y(n1159), .A(n1158) );
  ao22 U641 ( .Y(n1160), .A0(s_fractb_i_20_), .A1(n1904), .B0(s_fractb_i_18_), 
        .B1(n1901) );
  inv01 U642 ( .Y(n1161), .A(n1160) );
  nand02 U643 ( .Y(n2025), .A0(n1162), .A1(n1163) );
  inv01 U644 ( .Y(n1164), .A(n1901) );
  inv01 U645 ( .Y(n1165), .A(n1904) );
  inv01 U646 ( .Y(n1166), .A(s_fractb_i_13_) );
  inv01 U647 ( .Y(n1167), .A(s_fractb_i_11_) );
  nand02 U648 ( .Y(n1168), .A0(n1164), .A1(n1165) );
  nand02 U649 ( .Y(n1169), .A0(n1164), .A1(n1166) );
  nand02 U650 ( .Y(n1170), .A0(n1165), .A1(n1167) );
  nand02 U651 ( .Y(n1171), .A0(n1166), .A1(n1167) );
  nand02 U652 ( .Y(n1172), .A0(n1168), .A1(n1169) );
  inv01 U653 ( .Y(n1162), .A(n1172) );
  nand02 U654 ( .Y(n1173), .A0(n1170), .A1(n1171) );
  inv01 U655 ( .Y(n1163), .A(n1173) );
  nand02 U656 ( .Y(n2026), .A0(n1174), .A1(n1175) );
  inv01 U657 ( .Y(n1176), .A(n1901) );
  inv01 U658 ( .Y(n1177), .A(n1904) );
  inv01 U659 ( .Y(n1178), .A(s_fractb_i_21_) );
  inv01 U660 ( .Y(n1179), .A(s_fractb_i_19_) );
  nand02 U661 ( .Y(n1180), .A0(n1176), .A1(n1177) );
  nand02 U662 ( .Y(n1181), .A0(n1176), .A1(n1178) );
  nand02 U663 ( .Y(n1182), .A0(n1177), .A1(n1179) );
  nand02 U664 ( .Y(n1183), .A0(n1178), .A1(n1179) );
  nand02 U665 ( .Y(n1184), .A0(n1180), .A1(n1181) );
  inv01 U666 ( .Y(n1174), .A(n1184) );
  nand02 U667 ( .Y(n1185), .A0(n1182), .A1(n1183) );
  inv01 U668 ( .Y(n1175), .A(n1185) );
  nand02 U669 ( .Y(n2027), .A0(n1186), .A1(n1187) );
  inv01 U670 ( .Y(n1188), .A(n1901) );
  inv01 U671 ( .Y(n1189), .A(n1904) );
  inv01 U672 ( .Y(n1190), .A(s_fractb_i_5_) );
  inv01 U673 ( .Y(n1191), .A(s_fractb_i_3_) );
  nand02 U674 ( .Y(n1192), .A0(n1188), .A1(n1189) );
  nand02 U675 ( .Y(n1193), .A0(n1188), .A1(n1190) );
  nand02 U676 ( .Y(n1194), .A0(n1189), .A1(n1191) );
  nand02 U677 ( .Y(n1195), .A0(n1190), .A1(n1191) );
  nand02 U678 ( .Y(n1196), .A0(n1192), .A1(n1193) );
  inv01 U679 ( .Y(n1186), .A(n1196) );
  nand02 U680 ( .Y(n1197), .A0(n1194), .A1(n1195) );
  inv01 U681 ( .Y(n1187), .A(n1197) );
  ao22 U682 ( .Y(n1198), .A0(s_fractb_i_12_), .A1(n1904), .B0(s_fractb_i_10_), 
        .B1(n1901) );
  inv01 U683 ( .Y(n1199), .A(n1198) );
  ao22 U684 ( .Y(n1200), .A0(n1897), .A1(n1985), .B0(n1904), .B1(n1626) );
  inv01 U685 ( .Y(n1201), .A(n1200) );
  inv01 U686 ( .Y(n2013), .A(n1202) );
  nor02 U687 ( .Y(n1203), .A0(n1998), .A1(n1629) );
  nor02 U688 ( .Y(n1204), .A0(n1901), .A1(n1629) );
  nor02 U689 ( .Y(n1205), .A0(n1998), .A1(n1897) );
  nor02 U690 ( .Y(n1206), .A0(n1901), .A1(n1897) );
  nor02 U691 ( .Y(n1202), .A0(n1207), .A1(n1208) );
  nor02 U692 ( .Y(n1209), .A0(n1203), .A1(n1204) );
  inv01 U693 ( .Y(n1207), .A(n1209) );
  nor02 U694 ( .Y(n1210), .A0(n1205), .A1(n1206) );
  inv01 U695 ( .Y(n1208), .A(n1210) );
  ao22 U696 ( .Y(n1211), .A0(n1896), .A1(n1998), .B0(n1904), .B1(n1628) );
  inv01 U697 ( .Y(n1212), .A(n1211) );
  inv02 U698 ( .Y(n1998), .A(n1648) );
  ao22 U699 ( .Y(n1213), .A0(n1953), .A1(n1900), .B0(n2055), .B1(n1913) );
  inv01 U700 ( .Y(n1214), .A(n1213) );
  ao22 U701 ( .Y(n1215), .A0(n1902), .A1(v_prod_shl239_19_), .B0(
        n____return527_19_), .B1(n1916) );
  inv01 U702 ( .Y(n1216), .A(n1215) );
  ao22 U703 ( .Y(n1217), .A0(n1902), .A1(v_prod_shl239_17_), .B0(
        n____return527_17_), .B1(n1916) );
  inv01 U704 ( .Y(n1218), .A(n1217) );
  ao22 U705 ( .Y(n1219), .A0(n1902), .A1(v_prod_shl239_18_), .B0(
        n____return527_18_), .B1(n1916) );
  inv01 U706 ( .Y(n1220), .A(n1219) );
  ao22 U707 ( .Y(n1221), .A0(n1902), .A1(v_prod_shl239_21_), .B0(
        n____return527_21_), .B1(n1916) );
  inv01 U708 ( .Y(n1222), .A(n1221) );
  ao22 U709 ( .Y(n1223), .A0(n1902), .A1(v_prod_shl239_22_), .B0(
        n____return527_22_), .B1(n1916) );
  inv01 U710 ( .Y(n1224), .A(n1223) );
  ao22 U711 ( .Y(n1225), .A0(n1902), .A1(v_prod_shl239_20_), .B0(
        n____return527_20_), .B1(n1916) );
  inv01 U712 ( .Y(n1226), .A(n1225) );
  ao22 U713 ( .Y(n1227), .A0(n1902), .A1(v_prod_shl239_23_), .B0(
        n____return527_23_), .B1(n1916) );
  inv01 U714 ( .Y(n1228), .A(n1227) );
  ao22 U715 ( .Y(n1229), .A0(n1902), .A1(v_prod_shl239_13_), .B0(
        n____return527_13_), .B1(n1916) );
  inv01 U716 ( .Y(n1230), .A(n1229) );
  ao22 U717 ( .Y(n1231), .A0(n1902), .A1(v_prod_shl239_11_), .B0(
        n____return527_11_), .B1(n1916) );
  inv01 U718 ( .Y(n1232), .A(n1231) );
  ao22 U719 ( .Y(n1233), .A0(n1902), .A1(v_prod_shl239_14_), .B0(
        n____return527_14_), .B1(n1916) );
  inv01 U720 ( .Y(n1234), .A(n1233) );
  ao22 U721 ( .Y(n1235), .A0(n1902), .A1(v_prod_shl239_12_), .B0(
        n____return527_12_), .B1(n1916) );
  inv01 U722 ( .Y(n1236), .A(n1235) );
  buf02 U723 ( .Y(n1237), .A(n1999) );
  inv02 U724 ( .Y(n1238), .A(n1237) );
  inv01 U725 ( .Y(n2014), .A(n1239) );
  nor02 U726 ( .Y(n1240), .A0(n1910), .A1(n1852) );
  nor02 U727 ( .Y(n1241), .A0(n1950), .A1(n1869) );
  nor02 U728 ( .Y(n1239), .A0(n1240), .A1(n1241) );
  inv01 U729 ( .Y(n1982), .A(n1242) );
  nor02 U730 ( .Y(n1243), .A0(n1950), .A1(n1648) );
  nor02 U731 ( .Y(n1244), .A0(n1910), .A1(n1862) );
  nor02 U732 ( .Y(n1242), .A0(n1243), .A1(n1244) );
  inv04 U733 ( .Y(n1950), .A(n1727) );
  inv01 U734 ( .Y(n1996), .A(n1245) );
  nor02 U735 ( .Y(n1246), .A0(n1898), .A1(n1882) );
  nor02 U736 ( .Y(n1247), .A0(n1983), .A1(n1634) );
  nor02 U737 ( .Y(n1245), .A0(n1246), .A1(n1247) );
  inv08 U738 ( .Y(n1913), .A(n1912) );
  inv01 U739 ( .Y(n1989), .A(n1248) );
  nor02 U740 ( .Y(n1249), .A0(n1910), .A1(n1869) );
  nor02 U741 ( .Y(n1250), .A0(n1898), .A1(n1422) );
  nor02 U742 ( .Y(n1248), .A0(n1249), .A1(n1250) );
  nor02 U743 ( .Y(n1251), .A0(n1898), .A1(n1852) );
  inv02 U744 ( .Y(n1252), .A(n1251) );
  or02 U745 ( .Y(n1253), .A0(n1913), .A1(n1960) );
  inv01 U746 ( .Y(n1254), .A(n1253) );
  buf12 U747 ( .Y(n1914), .A(n1923) );
  inv02 U748 ( .Y(n1923), .A(n2016) );
  inv01 U749 ( .Y(n1039), .A(n1255) );
  nor02 U750 ( .Y(n1256), .A0(s_state132), .A1(n1957) );
  inv01 U751 ( .Y(n1257), .A(n1958) );
  nor02 U752 ( .Y(n1255), .A0(n1256), .A1(n1257) );
  inv01 U753 ( .Y(n1031), .A(n1258) );
  nor02 U754 ( .Y(n1259), .A0(n1900), .A1(n2035) );
  inv01 U755 ( .Y(n1260), .A(n1969) );
  nor02 U756 ( .Y(n1258), .A0(n1259), .A1(n1260) );
  inv01 U757 ( .Y(n1032), .A(n1261) );
  nor02 U758 ( .Y(n1262), .A0(n1900), .A1(n2036) );
  inv01 U759 ( .Y(n1263), .A(n1967) );
  nor02 U760 ( .Y(n1261), .A0(n1262), .A1(n1263) );
  inv01 U761 ( .Y(n1033), .A(n1264) );
  nor02 U762 ( .Y(n1265), .A0(n1900), .A1(n2037) );
  inv01 U763 ( .Y(n1266), .A(n1965) );
  nor02 U764 ( .Y(n1264), .A0(n1265), .A1(n1266) );
  inv01 U765 ( .Y(n1034), .A(n1267) );
  nor02 U766 ( .Y(n1268), .A0(n313_0_), .A1(n2038) );
  inv01 U767 ( .Y(n1269), .A(n1094) );
  nor02 U768 ( .Y(n1267), .A0(n1268), .A1(n1269) );
  inv01 U769 ( .Y(n1036), .A(n1270) );
  nor02 U770 ( .Y(n1271), .A0(n1900), .A1(n2044) );
  inv01 U771 ( .Y(n1272), .A(n1148) );
  nor02 U772 ( .Y(n1270), .A0(n1271), .A1(n1272) );
  inv01 U773 ( .Y(n1035), .A(n1273) );
  nor02 U774 ( .Y(n1274), .A0(n1900), .A1(n2039) );
  inv01 U775 ( .Y(n1275), .A(n1963) );
  nor02 U776 ( .Y(n1273), .A0(n1274), .A1(n1275) );
  inv01 U777 ( .Y(n1029), .A(n1276) );
  nor02 U778 ( .Y(n1277), .A0(n1900), .A1(n2033) );
  inv01 U779 ( .Y(n1278), .A(n1132) );
  nor02 U780 ( .Y(n1276), .A0(n1277), .A1(n1278) );
  inv01 U781 ( .Y(n1021), .A(n1279) );
  nor02 U782 ( .Y(n1280), .A0(n313_0_), .A1(n2048) );
  inv01 U783 ( .Y(n1281), .A(n1052) );
  nor02 U784 ( .Y(n1279), .A0(n1280), .A1(n1281) );
  inv01 U785 ( .Y(n1022), .A(n1282) );
  nor02 U786 ( .Y(n1283), .A0(n1900), .A1(n2049) );
  inv01 U787 ( .Y(n1284), .A(n1155) );
  nor02 U788 ( .Y(n1282), .A0(n1283), .A1(n1284) );
  inv01 U789 ( .Y(n1027), .A(n1285) );
  nor02 U790 ( .Y(n1286), .A0(n313_0_), .A1(n2054) );
  inv01 U791 ( .Y(n1287), .A(n1976) );
  nor02 U792 ( .Y(n1285), .A0(n1286), .A1(n1287) );
  inv01 U793 ( .Y(n1028), .A(n1288) );
  nor02 U794 ( .Y(n1289), .A0(n1900), .A1(n2032) );
  inv01 U795 ( .Y(n1290), .A(n1975) );
  nor02 U796 ( .Y(n1288), .A0(n1289), .A1(n1290) );
  inv01 U797 ( .Y(n1017), .A(n1291) );
  nor02 U798 ( .Y(n1292), .A0(n1900), .A1(n2043) );
  inv01 U799 ( .Y(n1293), .A(n1226) );
  nor02 U800 ( .Y(n1291), .A0(n1292), .A1(n1293) );
  inv01 U801 ( .Y(n1018), .A(n1294) );
  nor02 U802 ( .Y(n1295), .A0(n1900), .A1(n2045) );
  inv01 U803 ( .Y(n1296), .A(n1216) );
  nor02 U804 ( .Y(n1294), .A0(n1295), .A1(n1296) );
  inv01 U805 ( .Y(n1024), .A(n1297) );
  nor02 U806 ( .Y(n1298), .A0(n1900), .A1(n2051) );
  inv01 U807 ( .Y(n1299), .A(n1230) );
  nor02 U808 ( .Y(n1297), .A0(n1298), .A1(n1299) );
  inv01 U809 ( .Y(n1016), .A(n1300) );
  nor02 U810 ( .Y(n1301), .A0(n1900), .A1(n2042) );
  inv01 U811 ( .Y(n1302), .A(n1222) );
  nor02 U812 ( .Y(n1300), .A0(n1301), .A1(n1302) );
  inv01 U813 ( .Y(n1020), .A(n1303) );
  nor02 U814 ( .Y(n1304), .A0(n1900), .A1(n2047) );
  inv01 U815 ( .Y(n1305), .A(n1218) );
  nor02 U816 ( .Y(n1303), .A0(n1304), .A1(n1305) );
  inv01 U817 ( .Y(n1025), .A(n1306) );
  nor02 U818 ( .Y(n1307), .A0(n1900), .A1(n2052) );
  inv01 U819 ( .Y(n1308), .A(n1236) );
  nor02 U820 ( .Y(n1306), .A0(n1307), .A1(n1308) );
  inv01 U821 ( .Y(n1026), .A(n1309) );
  nor02 U822 ( .Y(n1310), .A0(n1900), .A1(n2053) );
  inv01 U823 ( .Y(n1311), .A(n1232) );
  nor02 U824 ( .Y(n1309), .A0(n1310), .A1(n1311) );
  inv01 U825 ( .Y(n1014), .A(n1312) );
  nor02 U826 ( .Y(n1313), .A0(n1900), .A1(n2040) );
  inv01 U827 ( .Y(n1314), .A(n1228) );
  nor02 U828 ( .Y(n1312), .A0(n1313), .A1(n1314) );
  inv01 U829 ( .Y(n1023), .A(n1315) );
  nor02 U830 ( .Y(n1316), .A0(n1900), .A1(n2050) );
  inv01 U831 ( .Y(n1317), .A(n1234) );
  nor02 U832 ( .Y(n1315), .A0(n1316), .A1(n1317) );
  inv01 U833 ( .Y(n1019), .A(n1318) );
  nor02 U834 ( .Y(n1319), .A0(n1900), .A1(n2046) );
  inv01 U835 ( .Y(n1320), .A(n1220) );
  nor02 U836 ( .Y(n1318), .A0(n1319), .A1(n1320) );
  inv01 U837 ( .Y(n1015), .A(n1321) );
  nor02 U838 ( .Y(n1322), .A0(n1900), .A1(n2041) );
  inv01 U839 ( .Y(n1323), .A(n1224) );
  nor02 U840 ( .Y(n1321), .A0(n1322), .A1(n1323) );
  inv01 U841 ( .Y(n1030), .A(n1324) );
  nor02 U842 ( .Y(n1325), .A0(n1900), .A1(n2034) );
  inv01 U843 ( .Y(n1326), .A(n1971) );
  nor02 U844 ( .Y(n1324), .A0(n1325), .A1(n1326) );
  inv02 U845 ( .Y(v_prod_shl239_0_), .A(n1953) );
  ao22 U846 ( .Y(n1327), .A0(n1903), .A1(n716), .B0(n1908), .B1(n717) );
  inv01 U847 ( .Y(n1328), .A(n1327) );
  inv02 U848 ( .Y(n1990), .A(n1328) );
  inv01 U849 ( .Y(n2006), .A(n1329) );
  nor02 U850 ( .Y(n1330), .A0(n1514), .A1(n1898) );
  nor02 U851 ( .Y(n1331), .A0(n1868), .A1(n1983) );
  nor02 U852 ( .Y(n1332), .A0(n1853), .A1(n1950) );
  nor02 U853 ( .Y(n1329), .A0(n1332), .A1(n1333) );
  nor02 U854 ( .Y(n1334), .A0(n1330), .A1(n1331) );
  inv01 U855 ( .Y(n1333), .A(n1334) );
  inv01 U856 ( .Y(n1949), .A(n1335) );
  nor02 U857 ( .Y(n1336), .A0(n1882), .A1(n1910) );
  nor02 U858 ( .Y(n1337), .A0(s_count[2]), .A1(n1926) );
  nor02 U859 ( .Y(n1338), .A0(n1538), .A1(n1950) );
  nor02 U860 ( .Y(n1335), .A0(n1338), .A1(n1339) );
  nor02 U861 ( .Y(n1340), .A0(n1336), .A1(n1337) );
  inv01 U862 ( .Y(n1339), .A(n1340) );
  inv04 U863 ( .Y(n1898), .A(n1897) );
  inv01 U864 ( .Y(n2003), .A(n1341) );
  nor02 U865 ( .Y(n1342), .A0(n1648), .A1(n1898) );
  nor02 U866 ( .Y(n1343), .A0(n1950), .A1(n1757) );
  nor02 U867 ( .Y(n1344), .A0(n1862), .A1(n1983) );
  nor02 U868 ( .Y(n1341), .A0(n1344), .A1(n1345) );
  nor02 U869 ( .Y(n1346), .A0(n1342), .A1(n1343) );
  inv01 U870 ( .Y(n1345), .A(n1346) );
  ao22 U871 ( .Y(n1347), .A0(n1972), .A1(n1760), .B0(n1973), .B1(n1892) );
  inv01 U872 ( .Y(n1348), .A(n1347) );
  inv01 U873 ( .Y(n2029), .A(n1349) );
  nor02 U874 ( .Y(n1350), .A0(n1910), .A1(n693) );
  nor02 U875 ( .Y(n1351), .A0(n1950), .A1(n692) );
  nor02 U876 ( .Y(n1352), .A0(n1983), .A1(n691) );
  nor02 U877 ( .Y(n1349), .A0(n1352), .A1(n1353) );
  nor02 U878 ( .Y(n1354), .A0(n1350), .A1(n1351) );
  inv01 U879 ( .Y(n1353), .A(n1354) );
  ao22 U880 ( .Y(n1355), .A0(n1936), .A1(n1760), .B0(n1937), .B1(n1539) );
  inv01 U881 ( .Y(n1356), .A(n1355) );
  ao22 U882 ( .Y(n1357), .A0(n1933), .A1(n1762), .B0(n1934), .B1(n1892) );
  inv01 U883 ( .Y(n1358), .A(n1357) );
  ao22 U884 ( .Y(n1359), .A0(n1931), .A1(n1760), .B0(n1932), .B1(n1892) );
  inv01 U885 ( .Y(n1360), .A(n1359) );
  inv02 U886 ( .Y(n1362), .A(n1361) );
  buf02 U887 ( .Y(n1363), .A(s_count[1]) );
  buf02 U888 ( .Y(n1366), .A(s_count[1]) );
  buf02 U889 ( .Y(n1364), .A(s_count[1]) );
  buf02 U890 ( .Y(n1365), .A(s_count[1]) );
  inv01 U891 ( .Y(n2022), .A(n1367) );
  nor02 U892 ( .Y(n1368), .A0(n1898), .A1(n690) );
  nor02 U893 ( .Y(n1369), .A0(n1910), .A1(n694) );
  inv01 U894 ( .Y(n1370), .A(n2027) );
  nor02 U895 ( .Y(n1367), .A0(n1370), .A1(n1371) );
  nor02 U896 ( .Y(n1372), .A0(n1368), .A1(n1369) );
  inv01 U897 ( .Y(n1371), .A(n1372) );
  inv01 U898 ( .Y(n2024), .A(n1373) );
  nor02 U899 ( .Y(n1374), .A0(n1898), .A1(n696) );
  nor02 U900 ( .Y(n1375), .A0(n1910), .A1(n698) );
  inv01 U901 ( .Y(n1376), .A(n2025) );
  nor02 U902 ( .Y(n1373), .A0(n1376), .A1(n1377) );
  nor02 U903 ( .Y(n1378), .A0(n1374), .A1(n1375) );
  inv01 U904 ( .Y(n1377), .A(n1378) );
  inv01 U905 ( .Y(n2023), .A(n1379) );
  nor02 U906 ( .Y(n1380), .A0(n1898), .A1(n700) );
  nor02 U907 ( .Y(n1381), .A0(n1910), .A1(n702) );
  inv01 U908 ( .Y(n1382), .A(n2026) );
  nor02 U909 ( .Y(n1379), .A0(n1382), .A1(n1383) );
  nor02 U910 ( .Y(n1384), .A0(n1380), .A1(n1381) );
  inv01 U911 ( .Y(n1383), .A(n1384) );
  inv01 U912 ( .Y(n2030), .A(n1385) );
  nor02 U913 ( .Y(n1386), .A0(n1898), .A1(n699) );
  nor02 U914 ( .Y(n1387), .A0(n1910), .A1(n701) );
  inv01 U915 ( .Y(n1388), .A(n1161) );
  nor02 U916 ( .Y(n1385), .A0(n1388), .A1(n1389) );
  nor02 U917 ( .Y(n1390), .A0(n1386), .A1(n1387) );
  inv01 U918 ( .Y(n1389), .A(n1390) );
  inv01 U919 ( .Y(n2028), .A(n1391) );
  nor02 U920 ( .Y(n1392), .A0(n1898), .A1(n695) );
  nor02 U921 ( .Y(n1393), .A0(n1910), .A1(n697) );
  inv01 U922 ( .Y(n1394), .A(n1199) );
  nor02 U923 ( .Y(n1391), .A0(n1394), .A1(n1395) );
  nor02 U924 ( .Y(n1396), .A0(n1392), .A1(n1393) );
  inv01 U925 ( .Y(n1395), .A(n1396) );
  inv01 U926 ( .Y(n1997), .A(n1397) );
  nor02 U927 ( .Y(n1398), .A0(n1875), .A1(n1983) );
  nor02 U928 ( .Y(n1399), .A0(n1984), .A1(n1898) );
  inv01 U929 ( .Y(n1400), .A(n1212) );
  nor02 U930 ( .Y(n1397), .A0(n1400), .A1(n1401) );
  nor02 U931 ( .Y(n1402), .A0(n1398), .A1(n1399) );
  inv01 U932 ( .Y(n1401), .A(n1402) );
  inv01 U933 ( .Y(n2004), .A(n1403) );
  nor02 U934 ( .Y(n1404), .A0(n1875), .A1(n1950) );
  nor02 U935 ( .Y(n1405), .A0(n1984), .A1(n1983) );
  inv01 U936 ( .Y(n1406), .A(n1051) );
  nor02 U937 ( .Y(n1403), .A0(n1406), .A1(n1407) );
  nor02 U938 ( .Y(n1408), .A0(n1404), .A1(n1405) );
  inv01 U939 ( .Y(n1407), .A(n1408) );
  inv04 U940 ( .Y(n1983), .A(n1901) );
  inv01 U941 ( .Y(n2012), .A(n1409) );
  nor02 U942 ( .Y(n1410), .A0(n1862), .A1(n1950) );
  nor02 U943 ( .Y(n1411), .A0(n1910), .A1(n1758) );
  inv01 U944 ( .Y(n1412), .A(n2013) );
  nor02 U945 ( .Y(n1409), .A0(n1412), .A1(n1413) );
  nor02 U946 ( .Y(n1414), .A0(n1410), .A1(n1411) );
  inv01 U947 ( .Y(n1413), .A(n1414) );
  inv01 U948 ( .Y(n2009), .A(n1415) );
  nor02 U949 ( .Y(n1416), .A0(n1875), .A1(n1910) );
  nor02 U950 ( .Y(n1417), .A0(n1984), .A1(n1950) );
  inv01 U951 ( .Y(n1418), .A(n1054) );
  nor02 U952 ( .Y(n1415), .A0(n1418), .A1(n1419) );
  nor02 U953 ( .Y(n1420), .A0(n1416), .A1(n1417) );
  inv01 U954 ( .Y(n1419), .A(n1420) );
  buf08 U955 ( .Y(n1910), .A(n1922) );
  ao22 U956 ( .Y(n1421), .A0(n1903), .A1(n710), .B0(n1909), .B1(n711) );
  inv02 U957 ( .Y(n1422), .A(n1421) );
  inv02 U958 ( .Y(n2001), .A(n1422) );
  ao22 U959 ( .Y(n1423), .A0(n1903), .A1(n720), .B0(n1907), .B1(n721) );
  inv01 U960 ( .Y(n1424), .A(n1423) );
  nand02 U961 ( .Y(n2021), .A0(n1425), .A1(n1426) );
  inv02 U962 ( .Y(n1427), .A(n2024) );
  inv02 U963 ( .Y(n1428), .A(n2023) );
  inv02 U964 ( .Y(n1429), .A(n2022) );
  inv02 U965 ( .Y(n1430), .A(n1642) );
  inv02 U966 ( .Y(n1431), .A(n1669) );
  nand02 U967 ( .Y(n1432), .A0(n1429), .A1(n1433) );
  nand02 U968 ( .Y(n1434), .A0(n1430), .A1(n1435) );
  nand02 U969 ( .Y(n1436), .A0(n1431), .A1(n1437) );
  nand02 U970 ( .Y(n1438), .A0(n1431), .A1(n1439) );
  nand02 U971 ( .Y(n1440), .A0(n1914), .A1(n1441) );
  nand02 U972 ( .Y(n1442), .A0(n1914), .A1(n1443) );
  nand02 U973 ( .Y(n1444), .A0(n1914), .A1(n1445) );
  nand02 U974 ( .Y(n1446), .A0(n1914), .A1(n1447) );
  nand02 U975 ( .Y(n1448), .A0(n1427), .A1(n1428) );
  inv01 U976 ( .Y(n1433), .A(n1448) );
  nand02 U977 ( .Y(n1449), .A0(n1427), .A1(n1428) );
  inv01 U978 ( .Y(n1435), .A(n1449) );
  nand02 U979 ( .Y(n1450), .A0(n1427), .A1(n1429) );
  inv01 U980 ( .Y(n1437), .A(n1450) );
  nand02 U981 ( .Y(n1451), .A0(n1427), .A1(n1430) );
  inv01 U982 ( .Y(n1439), .A(n1451) );
  nand02 U983 ( .Y(n1452), .A0(n1428), .A1(n1429) );
  inv01 U984 ( .Y(n1441), .A(n1452) );
  nand02 U985 ( .Y(n1453), .A0(n1428), .A1(n1430) );
  inv01 U986 ( .Y(n1443), .A(n1453) );
  nand02 U987 ( .Y(n1454), .A0(n1429), .A1(n1431) );
  inv01 U988 ( .Y(n1445), .A(n1454) );
  nand02 U989 ( .Y(n1455), .A0(n1430), .A1(n1431) );
  inv01 U990 ( .Y(n1447), .A(n1455) );
  nand02 U991 ( .Y(n1456), .A0(n1432), .A1(n1434) );
  inv01 U992 ( .Y(n1457), .A(n1456) );
  nand02 U993 ( .Y(n1458), .A0(n1436), .A1(n1438) );
  inv01 U994 ( .Y(n1459), .A(n1458) );
  nand02 U995 ( .Y(n1460), .A0(n1457), .A1(n1459) );
  inv01 U996 ( .Y(n1425), .A(n1460) );
  nand02 U997 ( .Y(n1461), .A0(n1440), .A1(n1442) );
  inv01 U998 ( .Y(n1462), .A(n1461) );
  nand02 U999 ( .Y(n1463), .A0(n1444), .A1(n1446) );
  inv01 U1000 ( .Y(n1464), .A(n1463) );
  nand02 U1001 ( .Y(n1465), .A0(n1462), .A1(n1464) );
  inv01 U1002 ( .Y(n1426), .A(n1465) );
  nand02 U1003 ( .Y(n2020), .A0(n1466), .A1(n1467) );
  inv02 U1004 ( .Y(n1468), .A(n2030) );
  inv02 U1005 ( .Y(n1469), .A(n2029) );
  inv02 U1006 ( .Y(n1470), .A(n2028) );
  inv02 U1007 ( .Y(n1471), .A(n1642) );
  inv02 U1008 ( .Y(n1472), .A(n1669) );
  nand02 U1009 ( .Y(n1473), .A0(n1470), .A1(n1474) );
  nand02 U1010 ( .Y(n1475), .A0(n1914), .A1(n1476) );
  nand02 U1011 ( .Y(n1477), .A0(n1471), .A1(n1478) );
  nand02 U1012 ( .Y(n1479), .A0(n1471), .A1(n1480) );
  nand02 U1013 ( .Y(n1481), .A0(n1472), .A1(n1482) );
  nand02 U1014 ( .Y(n1483), .A0(n1472), .A1(n1484) );
  nand02 U1015 ( .Y(n1485), .A0(n1472), .A1(n1486) );
  nand02 U1016 ( .Y(n1487), .A0(n1472), .A1(n1488) );
  nand02 U1017 ( .Y(n1489), .A0(n1468), .A1(n1469) );
  inv01 U1018 ( .Y(n1474), .A(n1489) );
  nand02 U1019 ( .Y(n1490), .A0(n1468), .A1(n1469) );
  inv01 U1020 ( .Y(n1476), .A(n1490) );
  nand02 U1021 ( .Y(n1491), .A0(n1468), .A1(n1470) );
  inv01 U1022 ( .Y(n1478), .A(n1491) );
  nand02 U1023 ( .Y(n1492), .A0(n1468), .A1(n1914) );
  inv01 U1024 ( .Y(n1480), .A(n1492) );
  nand02 U1025 ( .Y(n1493), .A0(n1469), .A1(n1470) );
  inv01 U1026 ( .Y(n1482), .A(n1493) );
  nand02 U1027 ( .Y(n1494), .A0(n1469), .A1(n1914) );
  inv01 U1028 ( .Y(n1484), .A(n1494) );
  nand02 U1029 ( .Y(n1495), .A0(n1470), .A1(n1471) );
  inv01 U1030 ( .Y(n1486), .A(n1495) );
  nand02 U1031 ( .Y(n1496), .A0(n1914), .A1(n1471) );
  inv01 U1032 ( .Y(n1488), .A(n1496) );
  nand02 U1033 ( .Y(n1497), .A0(n1473), .A1(n1475) );
  inv01 U1034 ( .Y(n1498), .A(n1497) );
  nand02 U1035 ( .Y(n1499), .A0(n1477), .A1(n1479) );
  inv01 U1036 ( .Y(n1500), .A(n1499) );
  nand02 U1037 ( .Y(n1501), .A0(n1498), .A1(n1500) );
  inv01 U1038 ( .Y(n1466), .A(n1501) );
  nand02 U1039 ( .Y(n1502), .A0(n1481), .A1(n1483) );
  inv01 U1040 ( .Y(n1503), .A(n1502) );
  nand02 U1041 ( .Y(n1504), .A0(n1485), .A1(n1487) );
  inv01 U1042 ( .Y(n1505), .A(n1504) );
  nand02 U1043 ( .Y(n1506), .A0(n1503), .A1(n1505) );
  inv01 U1044 ( .Y(n1467), .A(n1506) );
  inv01 U1045 ( .Y(n1978), .A(n1507) );
  nor02 U1046 ( .Y(n1508), .A0(n1915), .A1(n1509) );
  nor02 U1047 ( .Y(n1510), .A0(n1607), .A1(n1914) );
  nor02 U1048 ( .Y(n1507), .A0(n1508), .A1(n1510) );
  nor02 U1049 ( .Y(n1511), .A0(n1756), .A1(n1898) );
  inv01 U1050 ( .Y(n1509), .A(n1511) );
  inv01 U1051 ( .Y(n1512), .A(n1675) );
  ao22 U1052 ( .Y(n1513), .A0(n1903), .A1(n706), .B0(n1908), .B1(n707) );
  inv02 U1053 ( .Y(n1514), .A(n1513) );
  inv02 U1054 ( .Y(n1987), .A(n1514) );
  inv02 U1055 ( .Y(v_prod_shl239_29_), .A(n1515) );
  nor02 U1056 ( .Y(n1516), .A0(n1751), .A1(n1358) );
  nor02 U1057 ( .Y(n1517), .A0(n1866), .A1(n1915) );
  nor02 U1058 ( .Y(n1515), .A0(n1516), .A1(n1517) );
  buf02 U1059 ( .Y(n1518), .A(v_prod_shl239_35_) );
  inv02 U1060 ( .Y(v_prod_shl239_32_), .A(n1519) );
  nor02 U1061 ( .Y(n1520), .A0(n1920), .A1(n1914) );
  nor02 U1062 ( .Y(n1521), .A0(n1929), .A1(n1915) );
  nor02 U1063 ( .Y(n1519), .A0(n1520), .A1(n1521) );
  inv02 U1064 ( .Y(v_prod_shl239_31_), .A(n1522) );
  nor02 U1065 ( .Y(n1523), .A0(n1850), .A1(n1914) );
  nor02 U1066 ( .Y(n1524), .A0(n1856), .A1(n1915) );
  nor02 U1067 ( .Y(n1522), .A0(n1523), .A1(n1524) );
  inv02 U1068 ( .Y(v_prod_shl239_30_), .A(n1525) );
  nor02 U1069 ( .Y(n1526), .A0(n1751), .A1(n1360) );
  nor02 U1070 ( .Y(n1527), .A0(n1930), .A1(n1915) );
  nor02 U1071 ( .Y(n1525), .A0(n1526), .A1(n1527) );
  inv02 U1072 ( .Y(v_prod_shl239_28_), .A(n1528) );
  nor02 U1073 ( .Y(n1529), .A0(n1751), .A1(n1356) );
  nor02 U1074 ( .Y(n1530), .A0(n1935), .A1(n1915) );
  nor02 U1075 ( .Y(n1528), .A0(n1529), .A1(n1530) );
  inv02 U1076 ( .Y(v_prod_shl239_33_), .A(n1531) );
  nor02 U1077 ( .Y(n1532), .A0(n1919), .A1(n1914) );
  nor02 U1078 ( .Y(n1533), .A0(n1858), .A1(n1915) );
  nor02 U1079 ( .Y(n1531), .A0(n1532), .A1(n1533) );
  inv02 U1080 ( .Y(v_prod_shl239_34_), .A(n1534) );
  nor02 U1081 ( .Y(n1535), .A0(n1918), .A1(n1914) );
  nor02 U1082 ( .Y(n1536), .A0(n1871), .A1(n1915) );
  nor02 U1083 ( .Y(n1534), .A0(n1535), .A1(n1536) );
  ao22 U1084 ( .Y(n1537), .A0(n1903), .A1(n721), .B0(n1906), .B1(n722) );
  inv02 U1085 ( .Y(n1538), .A(n1537) );
  buf02 U1086 ( .Y(n1539), .A(n1892) );
  or02 U1087 ( .Y(n1540), .A0(n1920), .A1(n1915) );
  inv02 U1088 ( .Y(n1541), .A(n1540) );
  or02 U1089 ( .Y(n1542), .A0(n1661), .A1(n1915) );
  inv02 U1090 ( .Y(n1543), .A(n1542) );
  or02 U1091 ( .Y(n1544), .A0(n1850), .A1(n1915) );
  inv02 U1092 ( .Y(n1545), .A(n1544) );
  or02 U1093 ( .Y(n1546), .A0(n1919), .A1(n1915) );
  inv02 U1094 ( .Y(n1547), .A(n1546) );
  or02 U1095 ( .Y(n1548), .A0(n1918), .A1(n1915) );
  inv02 U1096 ( .Y(n1549), .A(n1548) );
  inv02 U1097 ( .Y(v_prod_shl239_27_), .A(n1550) );
  nor02 U1098 ( .Y(n1551), .A0(n1864), .A1(n1914) );
  nor02 U1099 ( .Y(n1552), .A0(n1661), .A1(n1911) );
  nor02 U1100 ( .Y(n1553), .A0(n1873), .A1(n1915) );
  nor02 U1101 ( .Y(n1550), .A0(n1553), .A1(n1554) );
  nor02 U1102 ( .Y(n1555), .A0(n1551), .A1(n1552) );
  inv01 U1103 ( .Y(n1554), .A(n1555) );
  inv01 U1104 ( .Y(n1936), .A(n1556) );
  nor02 U1105 ( .Y(n1557), .A0(n1670), .A1(n1910) );
  nor02 U1106 ( .Y(n1558), .A0(n1882), .A1(n1983) );
  inv01 U1107 ( .Y(n1559), .A(n1150) );
  nor02 U1108 ( .Y(n1556), .A0(n1559), .A1(n1560) );
  nor02 U1109 ( .Y(n1561), .A0(n1557), .A1(n1558) );
  inv01 U1110 ( .Y(n1560), .A(n1561) );
  nand02 U1111 ( .Y(n1933), .A0(n1151), .A1(n1562) );
  inv01 U1112 ( .Y(n1563), .A(n1910) );
  inv01 U1113 ( .Y(n1564), .A(n1328) );
  inv01 U1114 ( .Y(n1565), .A(n1983) );
  inv01 U1115 ( .Y(n1566), .A(n1424) );
  nand02 U1116 ( .Y(n1567), .A0(n1563), .A1(n1564) );
  nand02 U1117 ( .Y(n1568), .A0(n1565), .A1(n1566) );
  nand02 U1118 ( .Y(n1569), .A0(n1567), .A1(n1568) );
  inv01 U1119 ( .Y(n1562), .A(n1569) );
  or02 U1120 ( .Y(n1570), .A0(n1356), .A1(n1895) );
  inv02 U1121 ( .Y(n1571), .A(n1570) );
  inv01 U1122 ( .Y(n1931), .A(n1572) );
  nor02 U1123 ( .Y(n1573), .A0(n1882), .A1(n1950) );
  nor02 U1124 ( .Y(n1574), .A0(n1634), .A1(n1910) );
  inv01 U1125 ( .Y(n1575), .A(n1134) );
  nor02 U1126 ( .Y(n1572), .A0(n1575), .A1(n1576) );
  nor02 U1127 ( .Y(n1577), .A0(n1573), .A1(n1574) );
  inv01 U1128 ( .Y(n1576), .A(n1577) );
  inv02 U1129 ( .Y(v_prod_shl239_25_), .A(n1578) );
  nor02 U1130 ( .Y(n1579), .A0(n1860), .A1(n1915) );
  nor02 U1131 ( .Y(n1580), .A0(n1919), .A1(n1911) );
  nor02 U1132 ( .Y(n1581), .A0(n1858), .A1(n1914) );
  nor02 U1133 ( .Y(n1578), .A0(n1581), .A1(n1582) );
  nor02 U1134 ( .Y(n1583), .A0(n1579), .A1(n1580) );
  inv01 U1135 ( .Y(n1582), .A(n1583) );
  inv02 U1136 ( .Y(v_prod_shl239_26_), .A(n1584) );
  nor02 U1137 ( .Y(n1585), .A0(n1871), .A1(n1914) );
  nor02 U1138 ( .Y(n1586), .A0(n1918), .A1(n1911) );
  nor02 U1139 ( .Y(n1587), .A0(n1942), .A1(n1915) );
  nor02 U1140 ( .Y(n1584), .A0(n1587), .A1(n1588) );
  nor02 U1141 ( .Y(n1589), .A0(n1585), .A1(n1586) );
  inv01 U1142 ( .Y(n1588), .A(n1589) );
  or02 U1143 ( .Y(n1590), .A0(n1360), .A1(n1895) );
  inv02 U1144 ( .Y(n1591), .A(n1590) );
  or02 U1145 ( .Y(n1592), .A0(n1358), .A1(n1895) );
  inv02 U1146 ( .Y(n1593), .A(n1592) );
  inv02 U1147 ( .Y(v_prod_shl239_24_), .A(n1594) );
  nor02 U1148 ( .Y(n1595), .A0(n1929), .A1(n1914) );
  nor02 U1149 ( .Y(n1596), .A0(n1920), .A1(n1911) );
  nor02 U1150 ( .Y(n1597), .A0(n1348), .A1(n1894) );
  nor02 U1151 ( .Y(n1594), .A0(n1597), .A1(n1598) );
  nor02 U1152 ( .Y(n1599), .A0(n1595), .A1(n1596) );
  inv01 U1153 ( .Y(n1598), .A(n1599) );
  inv01 U1154 ( .Y(n1948), .A(n1600) );
  nor02 U1155 ( .Y(n1601), .A0(n1984), .A1(n1910) );
  nor02 U1156 ( .Y(n1602), .A0(n1670), .A1(n1983) );
  inv01 U1157 ( .Y(n1603), .A(n1201) );
  nor02 U1158 ( .Y(n1600), .A0(n1603), .A1(n1604) );
  nor02 U1159 ( .Y(n1605), .A0(n1601), .A1(n1602) );
  inv01 U1160 ( .Y(n1604), .A(n1605) );
  inv02 U1161 ( .Y(n1929), .A(n1948) );
  inv02 U1162 ( .Y(n1920), .A(n1949) );
  ao221 U1163 ( .Y(n1606), .A0(n1629), .A1(n1901), .B0(n1980), .B1(n1897), 
        .C0(n1982) );
  inv01 U1164 ( .Y(n1607), .A(n1606) );
  inv02 U1165 ( .Y(v_prod_shl239_36_), .A(n1608) );
  nor02 U1166 ( .Y(n1609), .A0(n1927), .A1(n1610) );
  nor02 U1167 ( .Y(n1611), .A0(n1928), .A1(n1915) );
  nor02 U1168 ( .Y(n1608), .A0(n1609), .A1(n1611) );
  nor02 U1169 ( .Y(n1612), .A0(n1914), .A1(n1926) );
  inv01 U1170 ( .Y(n1610), .A(n1612) );
  inv02 U1171 ( .Y(v_prod_shl239_37_), .A(n1613) );
  nor02 U1172 ( .Y(n1614), .A0(n1910), .A1(n1615) );
  nor02 U1173 ( .Y(n1616), .A0(n1925), .A1(n1915) );
  nor02 U1174 ( .Y(n1613), .A0(n1614), .A1(n1616) );
  nor02 U1175 ( .Y(n1617), .A0(n1914), .A1(n1646) );
  inv01 U1176 ( .Y(n1615), .A(n1617) );
  buf02 U1177 ( .Y(n1618), .A(n1988) );
  inv02 U1178 ( .Y(v_prod_shl239_38_), .A(n1619) );
  nor02 U1179 ( .Y(n1620), .A0(n1914), .A1(n1621) );
  nor02 U1180 ( .Y(n1622), .A0(n1924), .A1(n1915) );
  nor02 U1181 ( .Y(n1619), .A0(n1620), .A1(n1622) );
  nor02 U1182 ( .Y(n1623), .A0(n1921), .A1(n1910) );
  inv01 U1183 ( .Y(n1621), .A(n1623) );
  buf02 U1184 ( .Y(n1624), .A(n1991) );
  buf02 U1185 ( .Y(n1625), .A(n1986) );
  buf02 U1186 ( .Y(n1627), .A(n1986) );
  buf02 U1187 ( .Y(n1626), .A(n1986) );
  buf02 U1188 ( .Y(n1628), .A(n1979) );
  buf02 U1189 ( .Y(n1630), .A(n1979) );
  buf02 U1190 ( .Y(n1629), .A(n1979) );
  buf02 U1191 ( .Y(n1631), .A(n1994) );
  buf02 U1192 ( .Y(n1632), .A(n1993) );
  ao22 U1193 ( .Y(n1633), .A0(n1903), .A1(n717), .B0(n1907), .B1(n718) );
  inv02 U1194 ( .Y(n1634), .A(n1633) );
  nand02 U1195 ( .Y(n1635), .A0(n1955), .A1(n1913) );
  inv02 U1196 ( .Y(n1636), .A(n1635) );
  nand02 U1197 ( .Y(n1637), .A0(n1157), .A1(n1894) );
  nand02 U1198 ( .Y(n1639), .A0(n1159), .A1(n1894) );
  or02 U1199 ( .Y(n1641), .A0(n1752), .A1(n1762) );
  inv02 U1200 ( .Y(n1642), .A(n1641) );
  buf02 U1201 ( .Y(n1643), .A(n1940) );
  buf02 U1202 ( .Y(n1645), .A(n1940) );
  buf02 U1203 ( .Y(n1644), .A(n1940) );
  buf02 U1204 ( .Y(n1646), .A(n1046) );
  ao22 U1205 ( .Y(n1647), .A0(n1903), .A1(n705), .B0(n1907), .B1(n706) );
  inv02 U1206 ( .Y(n1648), .A(n1647) );
  buf02 U1207 ( .Y(n1649), .A(v_prod_shl239_16_) );
  buf02 U1208 ( .Y(n1650), .A(v_prod_shl239_16_) );
  inv01 U1209 ( .Y(n1651), .A(n1053) );
  inv01 U1210 ( .Y(n1652), .A(n1651) );
  inv02 U1211 ( .Y(n1653), .A(n1651) );
  inv02 U1212 ( .Y(v_prod_shl239_11_), .A(n1654) );
  nor02 U1213 ( .Y(n1655), .A0(n1873), .A1(n1911) );
  nor02 U1214 ( .Y(n1656), .A0(n1238), .A1(n1914) );
  nor02 U1215 ( .Y(n1654), .A0(n1655), .A1(n1656) );
  inv02 U1216 ( .Y(v_prod_shl239_13_), .A(n1657) );
  nor02 U1217 ( .Y(n1658), .A0(n1866), .A1(n1911) );
  nor02 U1218 ( .Y(n1659), .A0(n1968), .A1(n1914) );
  nor02 U1219 ( .Y(n1657), .A0(n1658), .A1(n1659) );
  ao22 U1220 ( .Y(n1660), .A0(n1939), .A1(n1904), .B0(n1644), .B1(n1896) );
  inv02 U1221 ( .Y(n1661), .A(n1660) );
  inv02 U1222 ( .Y(v_prod_shl239_14_), .A(n1662) );
  nor02 U1223 ( .Y(n1663), .A0(n1970), .A1(n1914) );
  nor02 U1224 ( .Y(n1664), .A0(n1930), .A1(n1911) );
  nor02 U1225 ( .Y(n1662), .A0(n1663), .A1(n1664) );
  inv02 U1226 ( .Y(v_prod_shl239_12_), .A(n1665) );
  nor02 U1227 ( .Y(n1666), .A0(n1935), .A1(n1911) );
  nor02 U1228 ( .Y(n1667), .A0(n1966), .A1(n1914) );
  nor02 U1229 ( .Y(n1665), .A0(n1666), .A1(n1667) );
  or02 U1230 ( .Y(n1668), .A0(n1895), .A1(n1759) );
  inv02 U1231 ( .Y(n1669), .A(n1668) );
  buf02 U1232 ( .Y(n1670), .A(n1044) );
  nand02 U1233 ( .Y(n1926), .A0(n1671), .A1(n1672) );
  inv01 U1234 ( .Y(n1673), .A(n1951) );
  inv01 U1235 ( .Y(n1674), .A(n1365) );
  inv01 U1236 ( .Y(n1675), .A(n1946) );
  inv01 U1237 ( .Y(n1676), .A(n1945) );
  nand02 U1238 ( .Y(n1677), .A0(n1673), .A1(n1674) );
  nand02 U1239 ( .Y(n1678), .A0(n1673), .A1(n1675) );
  nand02 U1240 ( .Y(n1679), .A0(n1674), .A1(n1676) );
  nand02 U1241 ( .Y(n1680), .A0(n1675), .A1(n1676) );
  nand02 U1242 ( .Y(n1681), .A0(n1677), .A1(n1678) );
  inv02 U1243 ( .Y(n1671), .A(n1681) );
  nand02 U1244 ( .Y(n1682), .A0(n1679), .A1(n1680) );
  inv02 U1245 ( .Y(n1672), .A(n1682) );
  inv02 U1246 ( .Y(n1951), .A(n1364) );
  inv02 U1247 ( .Y(v_prod_shl239_19_), .A(n1683) );
  nor02 U1248 ( .Y(n1684), .A0(n1238), .A1(n1915) );
  nor02 U1249 ( .Y(n1685), .A0(n1873), .A1(n1914) );
  nor02 U1250 ( .Y(n1686), .A0(n1864), .A1(n1911) );
  nor02 U1251 ( .Y(n1683), .A0(n1686), .A1(n1687) );
  nor02 U1252 ( .Y(n1688), .A0(n1684), .A1(n1685) );
  inv01 U1253 ( .Y(n1687), .A(n1688) );
  inv02 U1254 ( .Y(v_prod_shl239_17_), .A(n1689) );
  nor02 U1255 ( .Y(n1690), .A0(n1860), .A1(n1914) );
  nor02 U1256 ( .Y(n1691), .A0(n1915), .A1(n1252) );
  nor02 U1257 ( .Y(n1692), .A0(n1858), .A1(n1911) );
  nor02 U1258 ( .Y(n1689), .A0(n1692), .A1(n1693) );
  nor02 U1259 ( .Y(n1694), .A0(n1690), .A1(n1691) );
  inv01 U1260 ( .Y(n1693), .A(n1694) );
  inv02 U1261 ( .Y(v_prod_shl239_23_), .A(n1695) );
  nor02 U1262 ( .Y(n1696), .A0(n1764), .A1(n1915) );
  nor02 U1263 ( .Y(n1697), .A0(n1850), .A1(n1911) );
  nor02 U1264 ( .Y(n1698), .A0(n1856), .A1(n1914) );
  nor02 U1265 ( .Y(n1695), .A0(n1698), .A1(n1699) );
  nor02 U1266 ( .Y(n1700), .A0(n1696), .A1(n1697) );
  inv01 U1267 ( .Y(n1699), .A(n1700) );
  inv02 U1268 ( .Y(v_prod_shl239_20_), .A(n1701) );
  nor02 U1269 ( .Y(n1702), .A0(n1966), .A1(n1915) );
  nor02 U1270 ( .Y(n1703), .A0(n1935), .A1(n1914) );
  nor02 U1271 ( .Y(n1704), .A0(n1928), .A1(n1911) );
  nor02 U1272 ( .Y(n1701), .A0(n1704), .A1(n1705) );
  nor02 U1273 ( .Y(n1706), .A0(n1702), .A1(n1703) );
  inv01 U1274 ( .Y(n1705), .A(n1706) );
  inv02 U1275 ( .Y(v_prod_shl239_22_), .A(n1707) );
  nor02 U1276 ( .Y(n1708), .A0(n1930), .A1(n1914) );
  nor02 U1277 ( .Y(n1709), .A0(n1970), .A1(n1915) );
  nor02 U1278 ( .Y(n1710), .A0(n1924), .A1(n1911) );
  nor02 U1279 ( .Y(n1707), .A0(n1710), .A1(n1711) );
  nor02 U1280 ( .Y(n1712), .A0(n1708), .A1(n1709) );
  inv01 U1281 ( .Y(n1711), .A(n1712) );
  inv02 U1282 ( .Y(v_prod_shl239_21_), .A(n1713) );
  nor02 U1283 ( .Y(n1714), .A0(n1968), .A1(n1915) );
  nor02 U1284 ( .Y(n1715), .A0(n1866), .A1(n1914) );
  nor02 U1285 ( .Y(n1716), .A0(n1925), .A1(n1911) );
  nor02 U1286 ( .Y(n1713), .A0(n1716), .A1(n1717) );
  nor02 U1287 ( .Y(n1718), .A0(n1714), .A1(n1715) );
  inv01 U1288 ( .Y(n1717), .A(n1718) );
  inv02 U1289 ( .Y(n1935), .A(n2004) );
  inv02 U1290 ( .Y(n1966), .A(n2003) );
  inv02 U1291 ( .Y(n1970), .A(n2012) );
  inv02 U1292 ( .Y(n1930), .A(n2009) );
  inv02 U1293 ( .Y(n1968), .A(n2006) );
  inv02 U1294 ( .Y(v_prod_shl239_18_), .A(n1719) );
  nor02 U1295 ( .Y(n1720), .A0(n1871), .A1(n1911) );
  nor02 U1296 ( .Y(n1721), .A0(n1915), .A1(n1964) );
  nor02 U1297 ( .Y(n1722), .A0(n1942), .A1(n1914) );
  nor02 U1298 ( .Y(n1719), .A0(n1722), .A1(n1723) );
  nor02 U1299 ( .Y(n1724), .A0(n1720), .A1(n1721) );
  inv01 U1300 ( .Y(n1723), .A(n1724) );
  inv02 U1301 ( .Y(n1942), .A(n1997) );
  buf02 U1302 ( .Y(n1725), .A(v_prod_shl239_7_) );
  or02 U1303 ( .Y(n1726), .A0(n1927), .A1(n1364) );
  inv02 U1304 ( .Y(n1727), .A(n1726) );
  or02 U1305 ( .Y(n1728), .A0(n1964), .A1(n1911) );
  inv01 U1306 ( .Y(n1729), .A(n1728) );
  inv02 U1307 ( .Y(n1730), .A(n1728) );
  or02 U1308 ( .Y(n1731), .A0(n1252), .A1(n1911) );
  inv01 U1309 ( .Y(n1732), .A(n1731) );
  inv02 U1310 ( .Y(n1733), .A(n1731) );
  or02 U1311 ( .Y(n1734), .A0(n1348), .A1(n1752) );
  inv01 U1312 ( .Y(n1735), .A(n1734) );
  inv02 U1313 ( .Y(n1736), .A(n1734) );
  or02 U1314 ( .Y(n1737), .A0(n1911), .A1(n1238) );
  inv01 U1315 ( .Y(n1738), .A(n1737) );
  inv02 U1316 ( .Y(n1739), .A(n1737) );
  or02 U1317 ( .Y(n1740), .A0(n1911), .A1(n1970) );
  inv01 U1318 ( .Y(n1741), .A(n1740) );
  inv02 U1319 ( .Y(n1742), .A(n1740) );
  or02 U1320 ( .Y(n1743), .A0(n1911), .A1(n1966) );
  inv01 U1321 ( .Y(n1744), .A(n1743) );
  inv02 U1322 ( .Y(n1745), .A(n1743) );
  or02 U1323 ( .Y(n1746), .A0(n1911), .A1(n1968) );
  inv01 U1324 ( .Y(n1747), .A(n1746) );
  inv02 U1325 ( .Y(n1748), .A(n1746) );
  inv02 U1326 ( .Y(n1954), .A(n1956) );
  inv02 U1327 ( .Y(n1749), .A(s_count[4]) );
  inv02 U1328 ( .Y(n1750), .A(n1749) );
  inv02 U1329 ( .Y(n1752), .A(n1749) );
  inv02 U1330 ( .Y(n1751), .A(n1749) );
  inv02 U1331 ( .Y(n1754), .A(n1753) );
  inv02 U1332 ( .Y(n1755), .A(n1974) );
  inv02 U1333 ( .Y(n1756), .A(n1755) );
  inv02 U1334 ( .Y(n1758), .A(n1755) );
  inv01 U1335 ( .Y(n1757), .A(n1755) );
  inv02 U1336 ( .Y(n1927), .A(s_count[2]) );
  buf02 U1337 ( .Y(n1759), .A(s_count[3]) );
  buf02 U1338 ( .Y(n1762), .A(s_count[3]) );
  buf02 U1339 ( .Y(n1760), .A(s_count[3]) );
  buf02 U1340 ( .Y(n1761), .A(s_count[3]) );
  ao221 U1341 ( .Y(n1763), .A0(n1987), .A1(n1901), .B0(n1618), .B1(n1897), 
        .C0(n2014) );
  inv02 U1342 ( .Y(n1764), .A(n1763) );
  nand02 U1343 ( .Y(n1918), .A0(n1765), .A1(n1766) );
  inv02 U1344 ( .Y(n1767), .A(n1904) );
  inv02 U1345 ( .Y(n1768), .A(n1945) );
  inv02 U1346 ( .Y(n1769), .A(n1896) );
  inv02 U1347 ( .Y(n1770), .A(n1943) );
  inv02 U1348 ( .Y(n1771), .A(n1901) );
  inv02 U1349 ( .Y(n1772), .A(n1512) );
  nand02 U1350 ( .Y(n1773), .A0(n1769), .A1(n1774) );
  nand02 U1351 ( .Y(n1775), .A0(n1770), .A1(n1776) );
  nand02 U1352 ( .Y(n1777), .A0(n1771), .A1(n1778) );
  nand02 U1353 ( .Y(n1779), .A0(n1771), .A1(n1780) );
  nand02 U1354 ( .Y(n1781), .A0(n1772), .A1(n1782) );
  nand02 U1355 ( .Y(n1783), .A0(n1772), .A1(n1784) );
  nand02 U1356 ( .Y(n1785), .A0(n1772), .A1(n1786) );
  nand02 U1357 ( .Y(n1787), .A0(n1772), .A1(n1788) );
  nand02 U1358 ( .Y(n1789), .A0(n1767), .A1(n1768) );
  inv01 U1359 ( .Y(n1774), .A(n1789) );
  nand02 U1360 ( .Y(n1790), .A0(n1767), .A1(n1768) );
  inv01 U1361 ( .Y(n1776), .A(n1790) );
  nand02 U1362 ( .Y(n1791), .A0(n1767), .A1(n1769) );
  inv01 U1363 ( .Y(n1778), .A(n1791) );
  nand02 U1364 ( .Y(n1792), .A0(n1767), .A1(n1770) );
  inv01 U1365 ( .Y(n1780), .A(n1792) );
  nand02 U1366 ( .Y(n1793), .A0(n1768), .A1(n1769) );
  inv01 U1367 ( .Y(n1782), .A(n1793) );
  nand02 U1368 ( .Y(n1794), .A0(n1768), .A1(n1770) );
  inv01 U1369 ( .Y(n1784), .A(n1794) );
  nand02 U1370 ( .Y(n1795), .A0(n1769), .A1(n1771) );
  inv01 U1371 ( .Y(n1786), .A(n1795) );
  nand02 U1372 ( .Y(n1796), .A0(n1770), .A1(n1771) );
  inv01 U1373 ( .Y(n1788), .A(n1796) );
  nand02 U1374 ( .Y(n1797), .A0(n1773), .A1(n1775) );
  inv02 U1375 ( .Y(n1798), .A(n1797) );
  nand02 U1376 ( .Y(n1799), .A0(n1777), .A1(n1779) );
  inv02 U1377 ( .Y(n1800), .A(n1799) );
  nand02 U1378 ( .Y(n1801), .A0(n1798), .A1(n1800) );
  inv02 U1379 ( .Y(n1765), .A(n1801) );
  nand02 U1380 ( .Y(n1802), .A0(n1781), .A1(n1783) );
  inv02 U1381 ( .Y(n1803), .A(n1802) );
  nand02 U1382 ( .Y(n1804), .A0(n1785), .A1(n1787) );
  inv02 U1383 ( .Y(n1805), .A(n1804) );
  nand02 U1384 ( .Y(n1806), .A0(n1803), .A1(n1805) );
  inv02 U1385 ( .Y(n1766), .A(n1806) );
  inv02 U1386 ( .Y(n1943), .A(n1538) );
  nand02 U1387 ( .Y(n1919), .A0(n1807), .A1(n1808) );
  inv02 U1388 ( .Y(n1809), .A(n1896) );
  inv02 U1389 ( .Y(n1810), .A(n1904) );
  inv02 U1390 ( .Y(n1811), .A(n1901) );
  inv02 U1391 ( .Y(n1812), .A(n1939) );
  inv02 U1392 ( .Y(n1813), .A(n1644) );
  inv02 U1393 ( .Y(n1814), .A(n1947) );
  nand02 U1394 ( .Y(n1815), .A0(n1811), .A1(n1816) );
  nand02 U1395 ( .Y(n1817), .A0(n1812), .A1(n1818) );
  nand02 U1396 ( .Y(n1819), .A0(n1813), .A1(n1820) );
  nand02 U1397 ( .Y(n1821), .A0(n1813), .A1(n1822) );
  nand02 U1398 ( .Y(n1823), .A0(n1814), .A1(n1824) );
  nand02 U1399 ( .Y(n1825), .A0(n1814), .A1(n1826) );
  nand02 U1400 ( .Y(n1827), .A0(n1814), .A1(n1828) );
  nand02 U1401 ( .Y(n1829), .A0(n1814), .A1(n1830) );
  nand02 U1402 ( .Y(n1831), .A0(n1809), .A1(n1810) );
  inv01 U1403 ( .Y(n1816), .A(n1831) );
  nand02 U1404 ( .Y(n1832), .A0(n1809), .A1(n1810) );
  inv01 U1405 ( .Y(n1818), .A(n1832) );
  nand02 U1406 ( .Y(n1833), .A0(n1809), .A1(n1811) );
  inv01 U1407 ( .Y(n1820), .A(n1833) );
  nand02 U1408 ( .Y(n1834), .A0(n1809), .A1(n1812) );
  inv01 U1409 ( .Y(n1822), .A(n1834) );
  nand02 U1410 ( .Y(n1835), .A0(n1810), .A1(n1811) );
  inv01 U1411 ( .Y(n1824), .A(n1835) );
  nand02 U1412 ( .Y(n1836), .A0(n1810), .A1(n1812) );
  inv01 U1413 ( .Y(n1826), .A(n1836) );
  nand02 U1414 ( .Y(n1837), .A0(n1811), .A1(n1813) );
  inv01 U1415 ( .Y(n1828), .A(n1837) );
  nand02 U1416 ( .Y(n1838), .A0(n1812), .A1(n1813) );
  inv01 U1417 ( .Y(n1830), .A(n1838) );
  nand02 U1418 ( .Y(n1839), .A0(n1815), .A1(n1817) );
  inv02 U1419 ( .Y(n1840), .A(n1839) );
  nand02 U1420 ( .Y(n1841), .A0(n1819), .A1(n1821) );
  inv02 U1421 ( .Y(n1842), .A(n1841) );
  nand02 U1422 ( .Y(n1843), .A0(n1840), .A1(n1842) );
  inv02 U1423 ( .Y(n1807), .A(n1843) );
  nand02 U1424 ( .Y(n1844), .A0(n1823), .A1(n1825) );
  inv02 U1425 ( .Y(n1845), .A(n1844) );
  nand02 U1426 ( .Y(n1846), .A0(n1827), .A1(n1829) );
  inv01 U1427 ( .Y(n1847), .A(n1846) );
  nand02 U1428 ( .Y(n1848), .A0(n1845), .A1(n1847) );
  inv02 U1429 ( .Y(n1808), .A(n1848) );
  inv02 U1430 ( .Y(n1939), .A(n1646) );
  buf08 U1431 ( .Y(n1901), .A(n1944) );
  inv02 U1432 ( .Y(n1947), .A(n1424) );
  ao221 U1433 ( .Y(n1849), .A0(n1632), .A1(n1896), .B0(n1947), .B1(n1904), 
        .C0(n2015) );
  inv02 U1434 ( .Y(n1850), .A(n1849) );
  inv01 U1435 ( .Y(n1851), .A(n1056) );
  inv01 U1436 ( .Y(n1852), .A(n1851) );
  inv01 U1437 ( .Y(n1854), .A(n1851) );
  inv01 U1438 ( .Y(n1853), .A(n1851) );
  ao221 U1439 ( .Y(n1855), .A0(n1624), .A1(n1904), .B0(n2001), .B1(n1896), 
        .C0(n2017) );
  inv02 U1440 ( .Y(n1856), .A(n1855) );
  ao221 U1441 ( .Y(n1857), .A0(n1990), .A1(n1901), .B0(n1624), .B1(n1896), 
        .C0(n1992) );
  inv02 U1442 ( .Y(n1858), .A(n1857) );
  ao221 U1443 ( .Y(n1859), .A0(n1987), .A1(n1904), .B0(n1618), .B1(n1901), 
        .C0(n1989) );
  inv02 U1444 ( .Y(n1860), .A(n1859) );
  ao22 U1445 ( .Y(n1861), .A0(n1903), .A1(n703), .B0(n1906), .B1(n704) );
  inv02 U1446 ( .Y(n1862), .A(n1861) );
  ao221 U1447 ( .Y(n1863), .A0(n1631), .A1(n1896), .B0(n1990), .B1(n1904), 
        .C0(n2002) );
  inv02 U1448 ( .Y(n1864), .A(n1863) );
  ao221 U1449 ( .Y(n1865), .A0(n2001), .A1(n1727), .B0(n1618), .B1(n1896), 
        .C0(n2007) );
  inv02 U1450 ( .Y(n1866), .A(n1865) );
  ao22 U1451 ( .Y(n1867), .A0(n1903), .A1(n704), .B0(n1907), .B1(n705) );
  inv01 U1452 ( .Y(n1869), .A(n1867) );
  ao221 U1453 ( .Y(n1870), .A0(n1626), .A1(n1896), .B0(n1995), .B1(n1904), 
        .C0(n1996) );
  inv02 U1454 ( .Y(n1871), .A(n1870) );
  ao221 U1455 ( .Y(n1872), .A0(n1987), .A1(n1896), .B0(n1618), .B1(n1904), 
        .C0(n2000) );
  inv02 U1456 ( .Y(n1873), .A(n1872) );
  ao22 U1457 ( .Y(n1874), .A0(n1903), .A1(n709), .B0(n1906), .B1(n710) );
  inv02 U1458 ( .Y(n1875), .A(n1874) );
  inv02 U1459 ( .Y(n1960), .A(n1876) );
  inv01 U1460 ( .Y(n1877), .A(n1898) );
  inv01 U1461 ( .Y(n1878), .A(s_count[0]) );
  inv01 U1462 ( .Y(n1879), .A(n1911) );
  nand02 U1463 ( .Y(n1876), .A0(n1879), .A1(n1880) );
  nand02 U1464 ( .Y(n1881), .A0(n1877), .A1(n1878) );
  inv01 U1465 ( .Y(n1880), .A(n1881) );
  buf02 U1466 ( .Y(n1882), .A(n1042) );
  inv02 U1467 ( .Y(n1984), .A(n1883) );
  nor02 U1468 ( .Y(n1884), .A0(n1903), .A1(n712) );
  nor02 U1469 ( .Y(n1885), .A0(n711), .A1(n712) );
  nor02 U1470 ( .Y(n1886), .A0(n1903), .A1(n1909) );
  nor02 U1471 ( .Y(n1887), .A0(n711), .A1(n1909) );
  nor02 U1472 ( .Y(n1883), .A0(n1888), .A1(n1889) );
  nor02 U1473 ( .Y(n1890), .A0(n1884), .A1(n1885) );
  inv02 U1474 ( .Y(n1888), .A(n1890) );
  nor02 U1475 ( .Y(n1891), .A0(n1886), .A1(n1887) );
  inv01 U1476 ( .Y(n1889), .A(n1891) );
  inv02 U1477 ( .Y(n1909), .A(n1905) );
  buf02 U1478 ( .Y(n1893), .A(n1752) );
  inv02 U1479 ( .Y(n1894), .A(n1893) );
  inv02 U1480 ( .Y(n1895), .A(n1893) );
  buf12 U1481 ( .Y(n1896), .A(n1941) );
  buf08 U1482 ( .Y(n1897), .A(n1981) );
  inv04 U1483 ( .Y(n1899), .A(n313_0_) );
  inv12 U1484 ( .Y(n1900), .A(n1899) );
  buf16 U1485 ( .Y(n1902), .A(n1962) );
  buf08 U1486 ( .Y(n1903), .A(n1952) );
  inv08 U1487 ( .Y(n1904), .A(n1950) );
  inv02 U1488 ( .Y(n1905), .A(n2011) );
  inv02 U1489 ( .Y(n1906), .A(n1905) );
  inv02 U1490 ( .Y(n1907), .A(n1905) );
  inv02 U1491 ( .Y(n1908), .A(n1905) );
  buf12 U1492 ( .Y(n1911), .A(n1938) );
  buf02 U1493 ( .Y(n1912), .A(n1900) );
  buf16 U1494 ( .Y(n1915), .A(n1917) );
  buf16 U1495 ( .Y(n1916), .A(n1254) );
  oai22 U1496 ( .Y(v_prod_shl239_35_), .A0(n1864), .A1(n1915), .B0(n1661), 
        .B1(n1914) );
  nor02 U1497 ( .Y(n1932), .A0(n1910), .A1(n1921) );
  nor02 U1498 ( .Y(n1934), .A0(n1646), .A1(n1910) );
  nor02 U1499 ( .Y(n1937), .A0(n1926), .A1(n1927) );
  inv01 U1500 ( .Y(n1945), .A(n1921) );
  nand02 U1501 ( .Y(n1921), .A0(s_fracta_i_23_), .A1(n1903) );
  xor2 U1502 ( .Y(s_sign_o), .A0(signb_i), .A1(signa_i) );
  ao22 U1503 ( .Y(n999), .A0(s_fract_o[38]), .A1(n1913), .B0(
        n____return527_38_), .B1(n1916) );
  ao22 U1504 ( .Y(n998), .A0(s_fract_o[39]), .A1(n1913), .B0(
        n____return527_39_), .B1(n1916) );
  ao22 U1505 ( .Y(n997), .A0(s_fract_o[40]), .A1(n1913), .B0(
        n____return527_40_), .B1(n1916) );
  ao22 U1506 ( .Y(n996), .A0(s_fract_o[41]), .A1(n1913), .B0(
        n____return527_41_), .B1(n1916) );
  ao22 U1507 ( .Y(n995), .A0(s_fract_o[42]), .A1(n1913), .B0(
        n____return527_42_), .B1(n1916) );
  ao22 U1508 ( .Y(n994), .A0(s_fract_o[43]), .A1(n1913), .B0(
        n____return527_43_), .B1(n1916) );
  ao22 U1509 ( .Y(n993), .A0(s_fract_o[44]), .A1(n1913), .B0(
        n____return527_44_), .B1(n1916) );
  ao22 U1510 ( .Y(n992), .A0(s_fract_o[45]), .A1(n1913), .B0(
        n____return527_45_), .B1(n1916) );
  ao22 U1511 ( .Y(n991), .A0(s_fract_o[46]), .A1(n1913), .B0(
        n____return527_46_), .B1(n1916) );
  ao22 U1512 ( .Y(n990), .A0(s_fract_o[47]), .A1(n1913), .B0(
        n____return527_47_), .B1(n1916) );
  ao22 U1513 ( .Y(n989), .A0(sum218_4_), .A1(n1954), .B0(n1636), .B1(n1750) );
  ao22 U1514 ( .Y(n988), .A0(sum218_3_), .A1(n1954), .B0(n1636), .B1(n1759) );
  ao22 U1515 ( .Y(n987), .A0(sum218_2_), .A1(n1954), .B0(n1636), .B1(n1362) );
  ao22 U1516 ( .Y(n986), .A0(sum218_1_), .A1(n1954), .B0(n1636), .B1(n1363) );
  ao22 U1517 ( .Y(n985), .A0(sum218_0_), .A1(n1954), .B0(n1636), .B1(
        s_count[0]) );
  ao21 U1518 ( .Y(n1958), .A0(n1959), .A1(n1913), .B0(n2031) );
  nand02 U1519 ( .Y(n1038), .A0(n1959), .A1(n1956) );
  nand02 U1520 ( .Y(n1956), .A0(n1955), .A1(n1900) );
  and02 U1521 ( .Y(n1955), .A0(n1959), .A1(n1957) );
  nand03 U1522 ( .Y(n1957), .A0(n1669), .A1(n1896), .A2(s_count[0]) );
  inv01 U1523 ( .Y(n1959), .A(s_state132) );
  ao21 U1524 ( .Y(n1037), .A0(n____return527_0_), .A1(n1916), .B0(n1214) );
  nand03 U1525 ( .Y(n1953), .A0(n1960), .A1(n1050), .A2(s_fracta_i_0_) );
  nor02 U1526 ( .Y(v_prod_shl239_7_), .A0(n1911), .A1(n1764) );
  inv01 U1527 ( .Y(n1973), .A(n1607) );
  nor02 U1528 ( .Y(n1972), .A0(n1898), .A1(n1756) );
  oai22 U1529 ( .Y(v_prod_shl239_15_), .A0(n1764), .A1(n1914), .B0(n1856), 
        .B1(n1911) );
  aoi22 U1530 ( .Y(n1977), .A0(n1902), .A1(n1649), .B0(n____return527_16_), 
        .B1(n1916) );
  ao21 U1531 ( .Y(v_prod_shl239_16_), .A0(n1642), .A1(n1948), .B0(n1978) );
  inv01 U1532 ( .Y(n1980), .A(n1875) );
  ao22 U1533 ( .Y(n1992), .A0(n1897), .A1(n1632), .B0(n1904), .B1(n1631) );
  nand02 U1534 ( .Y(n1964), .A0(n1153), .A1(n1927) );
  ao22 U1535 ( .Y(n2000), .A0(n1897), .A1(n1624), .B0(n1901), .B1(n2001) );
  ao22 U1536 ( .Y(n2002), .A0(n1901), .A1(n1632), .B0(n1897), .B1(n1947) );
  aoi22 U1537 ( .Y(n2005), .A0(n1896), .A1(n1630), .B0(n1897), .B1(n1625) );
  inv01 U1538 ( .Y(n1928), .A(n1936) );
  inv01 U1539 ( .Y(n1985), .A(n1634) );
  ao22 U1540 ( .Y(n2007), .A0(n1897), .A1(n1631), .B0(n1901), .B1(n1624) );
  inv01 U1541 ( .Y(n1925), .A(n1933) );
  aoi22 U1542 ( .Y(n2008), .A0(n1897), .A1(n1645), .B0(n1904), .B1(n1632) );
  aoi22 U1543 ( .Y(n2010), .A0(n1901), .A1(n1627), .B0(n1897), .B1(n1995) );
  inv01 U1544 ( .Y(n1995), .A(n1670) );
  ao22 U1545 ( .Y(n1986), .A0(n1903), .A1(n713), .B0(n1906), .B1(n714) );
  ao22 U1546 ( .Y(n1979), .A0(n1903), .A1(n707), .B0(n1909), .B1(n708) );
  nand02 U1547 ( .Y(n1974), .A0(s_fracta_i_0_), .A1(n1907) );
  inv01 U1548 ( .Y(n1924), .A(n1931) );
  ao22 U1549 ( .Y(n1946), .A0(n1903), .A1(n723), .B0(n1908), .B1(n724) );
  inv01 U1550 ( .Y(n1917), .A(n1669) );
  ao22 U1551 ( .Y(n1988), .A0(n1903), .A1(n708), .B0(n1908), .B1(n709) );
  ao22 U1552 ( .Y(n2015), .A0(n1901), .A1(n1643), .B0(n1897), .B1(n1939) );
  ao22 U1553 ( .Y(n1940), .A0(n1903), .A1(n722), .B0(n1906), .B1(n723) );
  ao22 U1554 ( .Y(n1993), .A0(n1903), .A1(n718), .B0(n1908), .B1(n719) );
  ao22 U1555 ( .Y(n2017), .A0(n1901), .A1(n1631), .B0(n1897), .B1(n1990) );
  ao22 U1556 ( .Y(n1994), .A0(n1903), .A1(n714), .B0(n1909), .B1(n715) );
  ao22 U1557 ( .Y(n1991), .A0(n1903), .A1(n712), .B0(n1906), .B1(n713) );
  nor02 U1558 ( .Y(n2011), .A0(s_count[0]), .A1(n2018) );
  inv01 U1559 ( .Y(n2018), .A(n1961) );
  and02 U1560 ( .Y(n1952), .A0(s_count[0]), .A1(n1961) );
  ao21 U1561 ( .Y(n1961), .A0(n2056), .A1(n1960), .B0(n2019) );
  mux21 U1562 ( .Y(n2019), .A0(n2020), .A1(n2021), .S0(s_count[0]) );
  nor02 U1563 ( .Y(n1944), .A0(n1951), .A1(n1362) );
  inv01 U1564 ( .Y(n1922), .A(n1896) );
  nor02 U1565 ( .Y(n1941), .A0(n1951), .A1(n1927) );
  nor02 U1566 ( .Y(n2016), .A0(n1539), .A1(n1752) );
  and02 U1567 ( .Y(n1962), .A0(n1900), .A1(n1960) );
  ao22 U1568 ( .Y(n1013), .A0(s_fract_o[24]), .A1(n1913), .B0(
        n____return527_24_), .B1(n1916) );
  ao22 U1569 ( .Y(n1012), .A0(s_fract_o[25]), .A1(n1913), .B0(
        n____return527_25_), .B1(n1916) );
  ao22 U1570 ( .Y(n1011), .A0(s_fract_o[26]), .A1(n1913), .B0(
        n____return527_26_), .B1(n1916) );
  ao22 U1571 ( .Y(n1010), .A0(s_fract_o[27]), .A1(n1913), .B0(
        n____return527_27_), .B1(n1916) );
  ao22 U1572 ( .Y(n1009), .A0(s_fract_o[28]), .A1(n1913), .B0(
        n____return527_28_), .B1(n1916) );
  ao22 U1573 ( .Y(n1008), .A0(s_fract_o[29]), .A1(n1913), .B0(
        n____return527_29_), .B1(n1916) );
  ao22 U1574 ( .Y(n1007), .A0(s_fract_o[30]), .A1(n1913), .B0(
        n____return527_30_), .B1(n1916) );
  ao22 U1575 ( .Y(n1006), .A0(s_fract_o[31]), .A1(n1913), .B0(
        n____return527_31_), .B1(n1916) );
  ao22 U1576 ( .Y(n1005), .A0(s_fract_o[32]), .A1(n1913), .B0(
        n____return527_32_), .B1(n1916) );
  ao22 U1577 ( .Y(n1004), .A0(s_fract_o[33]), .A1(n1913), .B0(
        n____return527_33_), .B1(n1916) );
  ao22 U1578 ( .Y(n1003), .A0(s_fract_o[34]), .A1(n1913), .B0(
        n____return527_34_), .B1(n1916) );
  ao22 U1579 ( .Y(n1002), .A0(s_fract_o[35]), .A1(n1913), .B0(
        n____return527_35_), .B1(n1916) );
  ao22 U1580 ( .Y(n1001), .A0(s_fract_o[36]), .A1(n1913), .B0(
        n____return527_36_), .B1(n1916) );
  ao22 U1581 ( .Y(n1000), .A0(s_fract_o[37]), .A1(n1913), .B0(
        n____return527_37_), .B1(n1916) );
  nor02 U1582 ( .Y(n1981), .A0(n1362), .A1(n1366) );
  inv01 U1583 ( .Y(n1938), .A(n1642) );
  serial_mul_DW01_add_48_0 add_137_plus_plus ( .A({1'b0, n1591, n1593, n1571, 
        n1543, n1549, n1547, n1541, n1545, v_prod_shl239_38_, 
        v_prod_shl239_37_, v_prod_shl239_36_, n1518, v_prod_shl239_34_, 
        v_prod_shl239_33_, v_prod_shl239_32_, v_prod_shl239_31_, 
        v_prod_shl239_30_, v_prod_shl239_29_, v_prod_shl239_28_, 
        v_prod_shl239_27_, v_prod_shl239_26_, v_prod_shl239_25_, 
        v_prod_shl239_24_, v_prod_shl239_23_, v_prod_shl239_22_, 
        v_prod_shl239_21_, v_prod_shl239_20_, v_prod_shl239_19_, 
        v_prod_shl239_18_, v_prod_shl239_17_, n1650, n1653, v_prod_shl239_14_, 
        v_prod_shl239_13_, v_prod_shl239_12_, v_prod_shl239_11_, n1640, n1638, 
        n1736, n1725, n1742, n1748, n1745, n1739, n1730, n1733, 
        v_prod_shl239_0_}), .B(s_fract_o), .CI(1'b0), .SUM({n____return527_47_, 
        n____return527_46_, n____return527_45_, n____return527_44_, 
        n____return527_43_, n____return527_42_, n____return527_41_, 
        n____return527_40_, n____return527_39_, n____return527_38_, 
        n____return527_37_, n____return527_36_, n____return527_35_, 
        n____return527_34_, n____return527_33_, n____return527_32_, 
        n____return527_31_, n____return527_30_, n____return527_29_, 
        n____return527_28_, n____return527_27_, n____return527_26_, 
        n____return527_25_, n____return527_24_, n____return527_23_, 
        n____return527_22_, n____return527_21_, n____return527_20_, 
        n____return527_19_, n____return527_18_, n____return527_17_, 
        n____return527_16_, n____return527_15_, n____return527_14_, 
        n____return527_13_, n____return527_12_, n____return527_11_, 
        n____return527_10_, n____return527_9_, n____return527_8_, 
        n____return527_7_, n____return527_6_, n____return527_5_, 
        n____return527_4_, n____return527_3_, n____return527_2_, 
        n____return527_1_, n____return527_0_}) );
  serial_mul_DW01_inc_5_0 add_118 ( .A({n1750, n1761, n1362, n1363, n1754}), 
        .SUM({sum218_4_, sum218_3_, sum218_2_, sum218_1_, sum218_0_}) );
endmodule


module serial_div_DW01_sub_27_0 ( A, B, CI, DIFF, CO );
  input [26:0] A;
  input [26:0] B;
  output [26:0] DIFF;
  input CI;
  output CO;
  wire   carry_26_, carry_25_, carry_24_, carry_23_, carry_22_, carry_21_,
         carry_20_, carry_19_, carry_18_, carry_17_, carry_16_, carry_15_,
         carry_14_, carry_13_, carry_12_, carry_11_, carry_10_, carry_9_,
         carry_8_, carry_7_, carry_6_, carry_5_, carry_4_, carry_3_, carry_2_,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531;
  wire   [26:0] B_not;

  nor02 U6 ( .Y(n5), .A0(B_not[0]), .A1(A[0]) );
  inv02 U7 ( .Y(n6), .A(n5) );
  buf02 U8 ( .Y(n7), .A(carry_26_) );
  inv01 U9 ( .Y(DIFF[24]), .A(n8) );
  inv02 U10 ( .Y(carry_25_), .A(n9) );
  inv02 U11 ( .Y(n10), .A(B_not[24]) );
  inv02 U12 ( .Y(n11), .A(A[24]) );
  inv02 U13 ( .Y(n12), .A(n34) );
  nor02 U14 ( .Y(n13), .A0(n10), .A1(n14) );
  nor02 U15 ( .Y(n15), .A0(n11), .A1(n16) );
  nor02 U16 ( .Y(n17), .A0(n12), .A1(n18) );
  nor02 U17 ( .Y(n19), .A0(n12), .A1(n20) );
  nor02 U18 ( .Y(n8), .A0(n21), .A1(n22) );
  nor02 U19 ( .Y(n23), .A0(n11), .A1(n12) );
  nor02 U20 ( .Y(n24), .A0(n10), .A1(n12) );
  nor02 U21 ( .Y(n25), .A0(n10), .A1(n11) );
  nor02 U22 ( .Y(n9), .A0(n25), .A1(n26) );
  nor02 U23 ( .Y(n27), .A0(A[24]), .A1(n34) );
  inv01 U24 ( .Y(n14), .A(n27) );
  nor02 U25 ( .Y(n28), .A0(B_not[24]), .A1(n34) );
  inv01 U26 ( .Y(n16), .A(n28) );
  nor02 U27 ( .Y(n29), .A0(B_not[24]), .A1(A[24]) );
  inv01 U28 ( .Y(n18), .A(n29) );
  nor02 U29 ( .Y(n30), .A0(n10), .A1(n11) );
  inv01 U30 ( .Y(n20), .A(n30) );
  nor02 U31 ( .Y(n31), .A0(n13), .A1(n15) );
  inv01 U32 ( .Y(n21), .A(n31) );
  nor02 U33 ( .Y(n32), .A0(n17), .A1(n19) );
  inv01 U34 ( .Y(n22), .A(n32) );
  nor02 U35 ( .Y(n33), .A0(n23), .A1(n24) );
  inv01 U36 ( .Y(n26), .A(n33) );
  inv02 U37 ( .Y(B_not[24]), .A(B[24]) );
  buf02 U38 ( .Y(n34), .A(carry_24_) );
  buf02 U39 ( .Y(n35), .A(carry_23_) );
  buf02 U40 ( .Y(n36), .A(carry_22_) );
  inv01 U41 ( .Y(DIFF[20]), .A(n37) );
  inv02 U42 ( .Y(carry_21_), .A(n38) );
  inv02 U43 ( .Y(n39), .A(B_not[20]) );
  inv02 U44 ( .Y(n40), .A(A[20]) );
  inv02 U45 ( .Y(n41), .A(carry_20_) );
  nor02 U46 ( .Y(n42), .A0(n39), .A1(n43) );
  nor02 U47 ( .Y(n44), .A0(n40), .A1(n45) );
  nor02 U48 ( .Y(n46), .A0(n41), .A1(n47) );
  nor02 U49 ( .Y(n48), .A0(n41), .A1(n49) );
  nor02 U50 ( .Y(n37), .A0(n50), .A1(n51) );
  nor02 U51 ( .Y(n52), .A0(n40), .A1(n41) );
  nor02 U52 ( .Y(n53), .A0(n39), .A1(n41) );
  nor02 U53 ( .Y(n54), .A0(n39), .A1(n40) );
  nor02 U54 ( .Y(n38), .A0(n54), .A1(n55) );
  nor02 U55 ( .Y(n56), .A0(A[20]), .A1(carry_20_) );
  inv01 U56 ( .Y(n43), .A(n56) );
  nor02 U57 ( .Y(n57), .A0(B_not[20]), .A1(carry_20_) );
  inv01 U58 ( .Y(n45), .A(n57) );
  nor02 U59 ( .Y(n58), .A0(B_not[20]), .A1(A[20]) );
  inv01 U60 ( .Y(n47), .A(n58) );
  nor02 U61 ( .Y(n59), .A0(n39), .A1(n40) );
  inv01 U62 ( .Y(n49), .A(n59) );
  nor02 U63 ( .Y(n60), .A0(n42), .A1(n44) );
  inv01 U64 ( .Y(n50), .A(n60) );
  nor02 U65 ( .Y(n61), .A0(n46), .A1(n48) );
  inv01 U66 ( .Y(n51), .A(n61) );
  nor02 U67 ( .Y(n62), .A0(n52), .A1(n53) );
  inv01 U68 ( .Y(n55), .A(n62) );
  inv02 U69 ( .Y(B_not[20]), .A(B[20]) );
  inv01 U70 ( .Y(DIFF[19]), .A(n63) );
  inv02 U71 ( .Y(carry_20_), .A(n64) );
  inv02 U72 ( .Y(n65), .A(B_not[19]) );
  inv02 U73 ( .Y(n66), .A(A[19]) );
  inv02 U74 ( .Y(n67), .A(carry_19_) );
  nor02 U75 ( .Y(n68), .A0(n65), .A1(n69) );
  nor02 U76 ( .Y(n70), .A0(n66), .A1(n71) );
  nor02 U77 ( .Y(n72), .A0(n67), .A1(n73) );
  nor02 U78 ( .Y(n74), .A0(n67), .A1(n75) );
  nor02 U79 ( .Y(n63), .A0(n76), .A1(n77) );
  nor02 U80 ( .Y(n78), .A0(n66), .A1(n67) );
  nor02 U81 ( .Y(n79), .A0(n65), .A1(n67) );
  nor02 U82 ( .Y(n80), .A0(n65), .A1(n66) );
  nor02 U83 ( .Y(n64), .A0(n80), .A1(n81) );
  nor02 U84 ( .Y(n82), .A0(A[19]), .A1(carry_19_) );
  inv01 U85 ( .Y(n69), .A(n82) );
  nor02 U86 ( .Y(n83), .A0(B_not[19]), .A1(carry_19_) );
  inv01 U87 ( .Y(n71), .A(n83) );
  nor02 U88 ( .Y(n84), .A0(B_not[19]), .A1(A[19]) );
  inv01 U89 ( .Y(n73), .A(n84) );
  nor02 U90 ( .Y(n85), .A0(n65), .A1(n66) );
  inv01 U91 ( .Y(n75), .A(n85) );
  nor02 U92 ( .Y(n86), .A0(n68), .A1(n70) );
  inv01 U93 ( .Y(n76), .A(n86) );
  nor02 U94 ( .Y(n87), .A0(n72), .A1(n74) );
  inv01 U95 ( .Y(n77), .A(n87) );
  nor02 U96 ( .Y(n88), .A0(n78), .A1(n79) );
  inv01 U97 ( .Y(n81), .A(n88) );
  inv02 U98 ( .Y(B_not[19]), .A(B[19]) );
  inv01 U99 ( .Y(DIFF[18]), .A(n89) );
  inv02 U100 ( .Y(carry_19_), .A(n90) );
  inv02 U101 ( .Y(n91), .A(B_not[18]) );
  inv02 U102 ( .Y(n92), .A(A[18]) );
  inv02 U103 ( .Y(n93), .A(carry_18_) );
  nor02 U104 ( .Y(n94), .A0(n91), .A1(n95) );
  nor02 U105 ( .Y(n96), .A0(n92), .A1(n97) );
  nor02 U106 ( .Y(n98), .A0(n93), .A1(n99) );
  nor02 U107 ( .Y(n100), .A0(n93), .A1(n101) );
  nor02 U108 ( .Y(n89), .A0(n102), .A1(n103) );
  nor02 U109 ( .Y(n104), .A0(n92), .A1(n93) );
  nor02 U110 ( .Y(n105), .A0(n91), .A1(n93) );
  nor02 U111 ( .Y(n106), .A0(n91), .A1(n92) );
  nor02 U112 ( .Y(n90), .A0(n106), .A1(n107) );
  nor02 U113 ( .Y(n108), .A0(A[18]), .A1(carry_18_) );
  inv01 U114 ( .Y(n95), .A(n108) );
  nor02 U115 ( .Y(n109), .A0(B_not[18]), .A1(carry_18_) );
  inv01 U116 ( .Y(n97), .A(n109) );
  nor02 U117 ( .Y(n110), .A0(B_not[18]), .A1(A[18]) );
  inv01 U118 ( .Y(n99), .A(n110) );
  nor02 U119 ( .Y(n111), .A0(n91), .A1(n92) );
  inv01 U120 ( .Y(n101), .A(n111) );
  nor02 U121 ( .Y(n112), .A0(n94), .A1(n96) );
  inv01 U122 ( .Y(n102), .A(n112) );
  nor02 U123 ( .Y(n113), .A0(n98), .A1(n100) );
  inv01 U124 ( .Y(n103), .A(n113) );
  nor02 U125 ( .Y(n114), .A0(n104), .A1(n105) );
  inv01 U126 ( .Y(n107), .A(n114) );
  inv02 U127 ( .Y(B_not[18]), .A(B[18]) );
  inv01 U128 ( .Y(DIFF[17]), .A(n115) );
  inv02 U129 ( .Y(carry_18_), .A(n116) );
  inv02 U130 ( .Y(n117), .A(B_not[17]) );
  inv02 U131 ( .Y(n118), .A(A[17]) );
  inv02 U132 ( .Y(n119), .A(carry_17_) );
  nor02 U133 ( .Y(n120), .A0(n117), .A1(n121) );
  nor02 U134 ( .Y(n122), .A0(n118), .A1(n123) );
  nor02 U135 ( .Y(n124), .A0(n119), .A1(n125) );
  nor02 U136 ( .Y(n126), .A0(n119), .A1(n127) );
  nor02 U137 ( .Y(n115), .A0(n128), .A1(n129) );
  nor02 U138 ( .Y(n130), .A0(n118), .A1(n119) );
  nor02 U139 ( .Y(n131), .A0(n117), .A1(n119) );
  nor02 U140 ( .Y(n132), .A0(n117), .A1(n118) );
  nor02 U141 ( .Y(n116), .A0(n132), .A1(n133) );
  nor02 U142 ( .Y(n134), .A0(A[17]), .A1(carry_17_) );
  inv01 U143 ( .Y(n121), .A(n134) );
  nor02 U144 ( .Y(n135), .A0(B_not[17]), .A1(carry_17_) );
  inv01 U145 ( .Y(n123), .A(n135) );
  nor02 U146 ( .Y(n136), .A0(B_not[17]), .A1(A[17]) );
  inv01 U147 ( .Y(n125), .A(n136) );
  nor02 U148 ( .Y(n137), .A0(n117), .A1(n118) );
  inv01 U149 ( .Y(n127), .A(n137) );
  nor02 U150 ( .Y(n138), .A0(n120), .A1(n122) );
  inv01 U151 ( .Y(n128), .A(n138) );
  nor02 U152 ( .Y(n139), .A0(n124), .A1(n126) );
  inv01 U153 ( .Y(n129), .A(n139) );
  nor02 U154 ( .Y(n140), .A0(n130), .A1(n131) );
  inv01 U155 ( .Y(n133), .A(n140) );
  inv02 U156 ( .Y(B_not[17]), .A(B[17]) );
  inv01 U157 ( .Y(DIFF[16]), .A(n141) );
  inv02 U158 ( .Y(carry_17_), .A(n142) );
  inv02 U159 ( .Y(n143), .A(B_not[16]) );
  inv02 U160 ( .Y(n144), .A(A[16]) );
  inv02 U161 ( .Y(n145), .A(carry_16_) );
  nor02 U162 ( .Y(n146), .A0(n143), .A1(n147) );
  nor02 U163 ( .Y(n148), .A0(n144), .A1(n149) );
  nor02 U164 ( .Y(n150), .A0(n145), .A1(n151) );
  nor02 U165 ( .Y(n152), .A0(n145), .A1(n153) );
  nor02 U166 ( .Y(n141), .A0(n154), .A1(n155) );
  nor02 U167 ( .Y(n156), .A0(n144), .A1(n145) );
  nor02 U168 ( .Y(n157), .A0(n143), .A1(n145) );
  nor02 U169 ( .Y(n158), .A0(n143), .A1(n144) );
  nor02 U170 ( .Y(n142), .A0(n158), .A1(n159) );
  nor02 U171 ( .Y(n160), .A0(A[16]), .A1(carry_16_) );
  inv01 U172 ( .Y(n147), .A(n160) );
  nor02 U173 ( .Y(n161), .A0(B_not[16]), .A1(carry_16_) );
  inv01 U174 ( .Y(n149), .A(n161) );
  nor02 U175 ( .Y(n162), .A0(B_not[16]), .A1(A[16]) );
  inv01 U176 ( .Y(n151), .A(n162) );
  nor02 U177 ( .Y(n163), .A0(n143), .A1(n144) );
  inv01 U178 ( .Y(n153), .A(n163) );
  nor02 U179 ( .Y(n164), .A0(n146), .A1(n148) );
  inv01 U180 ( .Y(n154), .A(n164) );
  nor02 U181 ( .Y(n165), .A0(n150), .A1(n152) );
  inv01 U182 ( .Y(n155), .A(n165) );
  nor02 U183 ( .Y(n166), .A0(n156), .A1(n157) );
  inv01 U184 ( .Y(n159), .A(n166) );
  inv02 U185 ( .Y(B_not[16]), .A(B[16]) );
  inv01 U186 ( .Y(DIFF[15]), .A(n167) );
  inv02 U187 ( .Y(carry_16_), .A(n168) );
  inv02 U188 ( .Y(n169), .A(B_not[15]) );
  inv02 U189 ( .Y(n170), .A(A[15]) );
  inv02 U190 ( .Y(n171), .A(carry_15_) );
  nor02 U191 ( .Y(n172), .A0(n169), .A1(n173) );
  nor02 U192 ( .Y(n174), .A0(n170), .A1(n175) );
  nor02 U193 ( .Y(n176), .A0(n171), .A1(n177) );
  nor02 U194 ( .Y(n178), .A0(n171), .A1(n179) );
  nor02 U195 ( .Y(n167), .A0(n180), .A1(n181) );
  nor02 U196 ( .Y(n182), .A0(n170), .A1(n171) );
  nor02 U197 ( .Y(n183), .A0(n169), .A1(n171) );
  nor02 U198 ( .Y(n184), .A0(n169), .A1(n170) );
  nor02 U199 ( .Y(n168), .A0(n184), .A1(n185) );
  nor02 U200 ( .Y(n186), .A0(A[15]), .A1(carry_15_) );
  inv01 U201 ( .Y(n173), .A(n186) );
  nor02 U202 ( .Y(n187), .A0(B_not[15]), .A1(carry_15_) );
  inv01 U203 ( .Y(n175), .A(n187) );
  nor02 U204 ( .Y(n188), .A0(B_not[15]), .A1(A[15]) );
  inv01 U205 ( .Y(n177), .A(n188) );
  nor02 U206 ( .Y(n189), .A0(n169), .A1(n170) );
  inv01 U207 ( .Y(n179), .A(n189) );
  nor02 U208 ( .Y(n190), .A0(n172), .A1(n174) );
  inv01 U209 ( .Y(n180), .A(n190) );
  nor02 U210 ( .Y(n191), .A0(n176), .A1(n178) );
  inv01 U211 ( .Y(n181), .A(n191) );
  nor02 U212 ( .Y(n192), .A0(n182), .A1(n183) );
  inv01 U213 ( .Y(n185), .A(n192) );
  inv02 U214 ( .Y(B_not[15]), .A(B[15]) );
  inv01 U215 ( .Y(DIFF[14]), .A(n193) );
  inv02 U216 ( .Y(carry_15_), .A(n194) );
  inv02 U217 ( .Y(n195), .A(B_not[14]) );
  inv02 U218 ( .Y(n196), .A(A[14]) );
  inv02 U219 ( .Y(n197), .A(carry_14_) );
  nor02 U220 ( .Y(n198), .A0(n195), .A1(n199) );
  nor02 U221 ( .Y(n200), .A0(n196), .A1(n201) );
  nor02 U222 ( .Y(n202), .A0(n197), .A1(n203) );
  nor02 U223 ( .Y(n204), .A0(n197), .A1(n205) );
  nor02 U224 ( .Y(n193), .A0(n206), .A1(n207) );
  nor02 U225 ( .Y(n208), .A0(n196), .A1(n197) );
  nor02 U226 ( .Y(n209), .A0(n195), .A1(n197) );
  nor02 U227 ( .Y(n210), .A0(n195), .A1(n196) );
  nor02 U228 ( .Y(n194), .A0(n210), .A1(n211) );
  nor02 U229 ( .Y(n212), .A0(A[14]), .A1(carry_14_) );
  inv01 U230 ( .Y(n199), .A(n212) );
  nor02 U231 ( .Y(n213), .A0(B_not[14]), .A1(carry_14_) );
  inv01 U232 ( .Y(n201), .A(n213) );
  nor02 U233 ( .Y(n214), .A0(B_not[14]), .A1(A[14]) );
  inv01 U234 ( .Y(n203), .A(n214) );
  nor02 U235 ( .Y(n215), .A0(n195), .A1(n196) );
  inv01 U236 ( .Y(n205), .A(n215) );
  nor02 U237 ( .Y(n216), .A0(n198), .A1(n200) );
  inv01 U238 ( .Y(n206), .A(n216) );
  nor02 U239 ( .Y(n217), .A0(n202), .A1(n204) );
  inv01 U240 ( .Y(n207), .A(n217) );
  nor02 U241 ( .Y(n218), .A0(n208), .A1(n209) );
  inv01 U242 ( .Y(n211), .A(n218) );
  inv02 U243 ( .Y(B_not[14]), .A(B[14]) );
  inv01 U244 ( .Y(DIFF[13]), .A(n219) );
  inv02 U245 ( .Y(carry_14_), .A(n220) );
  inv02 U246 ( .Y(n221), .A(B_not[13]) );
  inv02 U247 ( .Y(n222), .A(A[13]) );
  inv02 U248 ( .Y(n223), .A(carry_13_) );
  nor02 U249 ( .Y(n224), .A0(n221), .A1(n225) );
  nor02 U250 ( .Y(n226), .A0(n222), .A1(n227) );
  nor02 U251 ( .Y(n228), .A0(n223), .A1(n229) );
  nor02 U252 ( .Y(n230), .A0(n223), .A1(n231) );
  nor02 U253 ( .Y(n219), .A0(n232), .A1(n233) );
  nor02 U254 ( .Y(n234), .A0(n222), .A1(n223) );
  nor02 U255 ( .Y(n235), .A0(n221), .A1(n223) );
  nor02 U256 ( .Y(n236), .A0(n221), .A1(n222) );
  nor02 U257 ( .Y(n220), .A0(n236), .A1(n237) );
  nor02 U258 ( .Y(n238), .A0(A[13]), .A1(carry_13_) );
  inv01 U259 ( .Y(n225), .A(n238) );
  nor02 U260 ( .Y(n239), .A0(B_not[13]), .A1(carry_13_) );
  inv01 U261 ( .Y(n227), .A(n239) );
  nor02 U262 ( .Y(n240), .A0(B_not[13]), .A1(A[13]) );
  inv01 U263 ( .Y(n229), .A(n240) );
  nor02 U264 ( .Y(n241), .A0(n221), .A1(n222) );
  inv01 U265 ( .Y(n231), .A(n241) );
  nor02 U266 ( .Y(n242), .A0(n224), .A1(n226) );
  inv01 U267 ( .Y(n232), .A(n242) );
  nor02 U268 ( .Y(n243), .A0(n228), .A1(n230) );
  inv01 U269 ( .Y(n233), .A(n243) );
  nor02 U270 ( .Y(n244), .A0(n234), .A1(n235) );
  inv01 U271 ( .Y(n237), .A(n244) );
  inv02 U272 ( .Y(B_not[13]), .A(B[13]) );
  inv01 U273 ( .Y(DIFF[12]), .A(n245) );
  inv02 U274 ( .Y(carry_13_), .A(n246) );
  inv02 U275 ( .Y(n247), .A(B_not[12]) );
  inv02 U276 ( .Y(n248), .A(A[12]) );
  inv02 U277 ( .Y(n249), .A(carry_12_) );
  nor02 U278 ( .Y(n250), .A0(n247), .A1(n251) );
  nor02 U279 ( .Y(n252), .A0(n248), .A1(n253) );
  nor02 U280 ( .Y(n254), .A0(n249), .A1(n255) );
  nor02 U281 ( .Y(n256), .A0(n249), .A1(n257) );
  nor02 U282 ( .Y(n245), .A0(n258), .A1(n259) );
  nor02 U283 ( .Y(n260), .A0(n248), .A1(n249) );
  nor02 U284 ( .Y(n261), .A0(n247), .A1(n249) );
  nor02 U285 ( .Y(n262), .A0(n247), .A1(n248) );
  nor02 U286 ( .Y(n246), .A0(n262), .A1(n263) );
  nor02 U287 ( .Y(n264), .A0(A[12]), .A1(carry_12_) );
  inv01 U288 ( .Y(n251), .A(n264) );
  nor02 U289 ( .Y(n265), .A0(B_not[12]), .A1(carry_12_) );
  inv01 U290 ( .Y(n253), .A(n265) );
  nor02 U291 ( .Y(n266), .A0(B_not[12]), .A1(A[12]) );
  inv01 U292 ( .Y(n255), .A(n266) );
  nor02 U293 ( .Y(n267), .A0(n247), .A1(n248) );
  inv01 U294 ( .Y(n257), .A(n267) );
  nor02 U295 ( .Y(n268), .A0(n250), .A1(n252) );
  inv01 U296 ( .Y(n258), .A(n268) );
  nor02 U297 ( .Y(n269), .A0(n254), .A1(n256) );
  inv01 U298 ( .Y(n259), .A(n269) );
  nor02 U299 ( .Y(n270), .A0(n260), .A1(n261) );
  inv01 U300 ( .Y(n263), .A(n270) );
  inv02 U301 ( .Y(B_not[12]), .A(B[12]) );
  inv01 U302 ( .Y(DIFF[11]), .A(n271) );
  inv02 U303 ( .Y(carry_12_), .A(n272) );
  inv02 U304 ( .Y(n273), .A(B_not[11]) );
  inv02 U305 ( .Y(n274), .A(A[11]) );
  inv02 U306 ( .Y(n275), .A(carry_11_) );
  nor02 U307 ( .Y(n276), .A0(n273), .A1(n277) );
  nor02 U308 ( .Y(n278), .A0(n274), .A1(n279) );
  nor02 U309 ( .Y(n280), .A0(n275), .A1(n281) );
  nor02 U310 ( .Y(n282), .A0(n275), .A1(n283) );
  nor02 U311 ( .Y(n271), .A0(n284), .A1(n285) );
  nor02 U312 ( .Y(n286), .A0(n274), .A1(n275) );
  nor02 U313 ( .Y(n287), .A0(n273), .A1(n275) );
  nor02 U314 ( .Y(n288), .A0(n273), .A1(n274) );
  nor02 U315 ( .Y(n272), .A0(n288), .A1(n289) );
  nor02 U316 ( .Y(n290), .A0(A[11]), .A1(carry_11_) );
  inv01 U317 ( .Y(n277), .A(n290) );
  nor02 U318 ( .Y(n291), .A0(B_not[11]), .A1(carry_11_) );
  inv01 U319 ( .Y(n279), .A(n291) );
  nor02 U320 ( .Y(n292), .A0(B_not[11]), .A1(A[11]) );
  inv01 U321 ( .Y(n281), .A(n292) );
  nor02 U322 ( .Y(n293), .A0(n273), .A1(n274) );
  inv01 U323 ( .Y(n283), .A(n293) );
  nor02 U324 ( .Y(n294), .A0(n276), .A1(n278) );
  inv01 U325 ( .Y(n284), .A(n294) );
  nor02 U326 ( .Y(n295), .A0(n280), .A1(n282) );
  inv01 U327 ( .Y(n285), .A(n295) );
  nor02 U328 ( .Y(n296), .A0(n286), .A1(n287) );
  inv01 U329 ( .Y(n289), .A(n296) );
  inv02 U330 ( .Y(B_not[11]), .A(B[11]) );
  inv01 U331 ( .Y(DIFF[10]), .A(n297) );
  inv02 U332 ( .Y(carry_11_), .A(n298) );
  inv02 U333 ( .Y(n299), .A(B_not[10]) );
  inv02 U334 ( .Y(n300), .A(A[10]) );
  inv02 U335 ( .Y(n301), .A(carry_10_) );
  nor02 U336 ( .Y(n302), .A0(n299), .A1(n303) );
  nor02 U337 ( .Y(n304), .A0(n300), .A1(n305) );
  nor02 U338 ( .Y(n306), .A0(n301), .A1(n307) );
  nor02 U339 ( .Y(n308), .A0(n301), .A1(n309) );
  nor02 U340 ( .Y(n297), .A0(n310), .A1(n311) );
  nor02 U341 ( .Y(n312), .A0(n300), .A1(n301) );
  nor02 U342 ( .Y(n313), .A0(n299), .A1(n301) );
  nor02 U343 ( .Y(n314), .A0(n299), .A1(n300) );
  nor02 U344 ( .Y(n298), .A0(n314), .A1(n315) );
  nor02 U345 ( .Y(n316), .A0(A[10]), .A1(carry_10_) );
  inv01 U346 ( .Y(n303), .A(n316) );
  nor02 U347 ( .Y(n317), .A0(B_not[10]), .A1(carry_10_) );
  inv01 U348 ( .Y(n305), .A(n317) );
  nor02 U349 ( .Y(n318), .A0(B_not[10]), .A1(A[10]) );
  inv01 U350 ( .Y(n307), .A(n318) );
  nor02 U351 ( .Y(n319), .A0(n299), .A1(n300) );
  inv01 U352 ( .Y(n309), .A(n319) );
  nor02 U353 ( .Y(n320), .A0(n302), .A1(n304) );
  inv01 U354 ( .Y(n310), .A(n320) );
  nor02 U355 ( .Y(n321), .A0(n306), .A1(n308) );
  inv01 U356 ( .Y(n311), .A(n321) );
  nor02 U357 ( .Y(n322), .A0(n312), .A1(n313) );
  inv01 U358 ( .Y(n315), .A(n322) );
  inv02 U359 ( .Y(B_not[10]), .A(B[10]) );
  inv01 U360 ( .Y(DIFF[9]), .A(n323) );
  inv02 U361 ( .Y(carry_10_), .A(n324) );
  inv02 U362 ( .Y(n325), .A(B_not[9]) );
  inv02 U363 ( .Y(n326), .A(A[9]) );
  inv02 U364 ( .Y(n327), .A(carry_9_) );
  nor02 U365 ( .Y(n328), .A0(n325), .A1(n329) );
  nor02 U366 ( .Y(n330), .A0(n326), .A1(n331) );
  nor02 U367 ( .Y(n332), .A0(n327), .A1(n333) );
  nor02 U368 ( .Y(n334), .A0(n327), .A1(n335) );
  nor02 U369 ( .Y(n323), .A0(n336), .A1(n337) );
  nor02 U370 ( .Y(n338), .A0(n326), .A1(n327) );
  nor02 U371 ( .Y(n339), .A0(n325), .A1(n327) );
  nor02 U372 ( .Y(n340), .A0(n325), .A1(n326) );
  nor02 U373 ( .Y(n324), .A0(n340), .A1(n341) );
  nor02 U374 ( .Y(n342), .A0(A[9]), .A1(carry_9_) );
  inv01 U375 ( .Y(n329), .A(n342) );
  nor02 U376 ( .Y(n343), .A0(B_not[9]), .A1(carry_9_) );
  inv01 U377 ( .Y(n331), .A(n343) );
  nor02 U378 ( .Y(n344), .A0(B_not[9]), .A1(A[9]) );
  inv01 U379 ( .Y(n333), .A(n344) );
  nor02 U380 ( .Y(n345), .A0(n325), .A1(n326) );
  inv01 U381 ( .Y(n335), .A(n345) );
  nor02 U382 ( .Y(n346), .A0(n328), .A1(n330) );
  inv01 U383 ( .Y(n336), .A(n346) );
  nor02 U384 ( .Y(n347), .A0(n332), .A1(n334) );
  inv01 U385 ( .Y(n337), .A(n347) );
  nor02 U386 ( .Y(n348), .A0(n338), .A1(n339) );
  inv01 U387 ( .Y(n341), .A(n348) );
  inv02 U388 ( .Y(B_not[9]), .A(B[9]) );
  inv01 U389 ( .Y(DIFF[8]), .A(n349) );
  inv02 U390 ( .Y(carry_9_), .A(n350) );
  inv02 U391 ( .Y(n351), .A(B_not[8]) );
  inv02 U392 ( .Y(n352), .A(A[8]) );
  inv02 U393 ( .Y(n353), .A(carry_8_) );
  nor02 U394 ( .Y(n354), .A0(n351), .A1(n355) );
  nor02 U395 ( .Y(n356), .A0(n352), .A1(n357) );
  nor02 U396 ( .Y(n358), .A0(n353), .A1(n359) );
  nor02 U397 ( .Y(n360), .A0(n353), .A1(n361) );
  nor02 U398 ( .Y(n349), .A0(n362), .A1(n363) );
  nor02 U399 ( .Y(n364), .A0(n352), .A1(n353) );
  nor02 U400 ( .Y(n365), .A0(n351), .A1(n353) );
  nor02 U401 ( .Y(n366), .A0(n351), .A1(n352) );
  nor02 U402 ( .Y(n350), .A0(n366), .A1(n367) );
  nor02 U403 ( .Y(n368), .A0(A[8]), .A1(carry_8_) );
  inv01 U404 ( .Y(n355), .A(n368) );
  nor02 U405 ( .Y(n369), .A0(B_not[8]), .A1(carry_8_) );
  inv01 U406 ( .Y(n357), .A(n369) );
  nor02 U407 ( .Y(n370), .A0(B_not[8]), .A1(A[8]) );
  inv01 U408 ( .Y(n359), .A(n370) );
  nor02 U409 ( .Y(n371), .A0(n351), .A1(n352) );
  inv01 U410 ( .Y(n361), .A(n371) );
  nor02 U411 ( .Y(n372), .A0(n354), .A1(n356) );
  inv01 U412 ( .Y(n362), .A(n372) );
  nor02 U413 ( .Y(n373), .A0(n358), .A1(n360) );
  inv01 U414 ( .Y(n363), .A(n373) );
  nor02 U415 ( .Y(n374), .A0(n364), .A1(n365) );
  inv01 U416 ( .Y(n367), .A(n374) );
  inv02 U417 ( .Y(B_not[8]), .A(B[8]) );
  inv01 U418 ( .Y(DIFF[7]), .A(n375) );
  inv02 U419 ( .Y(carry_8_), .A(n376) );
  inv02 U420 ( .Y(n377), .A(B_not[7]) );
  inv02 U421 ( .Y(n378), .A(A[7]) );
  inv02 U422 ( .Y(n379), .A(carry_7_) );
  nor02 U423 ( .Y(n380), .A0(n377), .A1(n381) );
  nor02 U424 ( .Y(n382), .A0(n378), .A1(n383) );
  nor02 U425 ( .Y(n384), .A0(n379), .A1(n385) );
  nor02 U426 ( .Y(n386), .A0(n379), .A1(n387) );
  nor02 U427 ( .Y(n375), .A0(n388), .A1(n389) );
  nor02 U428 ( .Y(n390), .A0(n378), .A1(n379) );
  nor02 U429 ( .Y(n391), .A0(n377), .A1(n379) );
  nor02 U430 ( .Y(n392), .A0(n377), .A1(n378) );
  nor02 U431 ( .Y(n376), .A0(n392), .A1(n393) );
  nor02 U432 ( .Y(n394), .A0(A[7]), .A1(carry_7_) );
  inv01 U433 ( .Y(n381), .A(n394) );
  nor02 U434 ( .Y(n395), .A0(B_not[7]), .A1(carry_7_) );
  inv01 U435 ( .Y(n383), .A(n395) );
  nor02 U436 ( .Y(n396), .A0(B_not[7]), .A1(A[7]) );
  inv01 U437 ( .Y(n385), .A(n396) );
  nor02 U438 ( .Y(n397), .A0(n377), .A1(n378) );
  inv01 U439 ( .Y(n387), .A(n397) );
  nor02 U440 ( .Y(n398), .A0(n380), .A1(n382) );
  inv01 U441 ( .Y(n388), .A(n398) );
  nor02 U442 ( .Y(n399), .A0(n384), .A1(n386) );
  inv01 U443 ( .Y(n389), .A(n399) );
  nor02 U444 ( .Y(n400), .A0(n390), .A1(n391) );
  inv01 U445 ( .Y(n393), .A(n400) );
  inv02 U446 ( .Y(B_not[7]), .A(B[7]) );
  inv01 U447 ( .Y(DIFF[6]), .A(n401) );
  inv02 U448 ( .Y(carry_7_), .A(n402) );
  inv02 U449 ( .Y(n403), .A(B_not[6]) );
  inv02 U450 ( .Y(n404), .A(A[6]) );
  inv02 U451 ( .Y(n405), .A(carry_6_) );
  nor02 U452 ( .Y(n406), .A0(n403), .A1(n407) );
  nor02 U453 ( .Y(n408), .A0(n404), .A1(n409) );
  nor02 U454 ( .Y(n410), .A0(n405), .A1(n411) );
  nor02 U455 ( .Y(n412), .A0(n405), .A1(n413) );
  nor02 U456 ( .Y(n401), .A0(n414), .A1(n415) );
  nor02 U457 ( .Y(n416), .A0(n404), .A1(n405) );
  nor02 U458 ( .Y(n417), .A0(n403), .A1(n405) );
  nor02 U459 ( .Y(n418), .A0(n403), .A1(n404) );
  nor02 U460 ( .Y(n402), .A0(n418), .A1(n419) );
  nor02 U461 ( .Y(n420), .A0(A[6]), .A1(carry_6_) );
  inv01 U462 ( .Y(n407), .A(n420) );
  nor02 U463 ( .Y(n421), .A0(B_not[6]), .A1(carry_6_) );
  inv01 U464 ( .Y(n409), .A(n421) );
  nor02 U465 ( .Y(n422), .A0(B_not[6]), .A1(A[6]) );
  inv01 U466 ( .Y(n411), .A(n422) );
  nor02 U467 ( .Y(n423), .A0(n403), .A1(n404) );
  inv01 U468 ( .Y(n413), .A(n423) );
  nor02 U469 ( .Y(n424), .A0(n406), .A1(n408) );
  inv01 U470 ( .Y(n414), .A(n424) );
  nor02 U471 ( .Y(n425), .A0(n410), .A1(n412) );
  inv01 U472 ( .Y(n415), .A(n425) );
  nor02 U473 ( .Y(n426), .A0(n416), .A1(n417) );
  inv01 U474 ( .Y(n419), .A(n426) );
  inv02 U475 ( .Y(B_not[6]), .A(B[6]) );
  inv01 U476 ( .Y(DIFF[5]), .A(n427) );
  inv02 U477 ( .Y(carry_6_), .A(n428) );
  inv02 U478 ( .Y(n429), .A(B_not[5]) );
  inv02 U479 ( .Y(n430), .A(A[5]) );
  inv02 U480 ( .Y(n431), .A(carry_5_) );
  nor02 U481 ( .Y(n432), .A0(n429), .A1(n433) );
  nor02 U482 ( .Y(n434), .A0(n430), .A1(n435) );
  nor02 U483 ( .Y(n436), .A0(n431), .A1(n437) );
  nor02 U484 ( .Y(n438), .A0(n431), .A1(n439) );
  nor02 U485 ( .Y(n427), .A0(n440), .A1(n441) );
  nor02 U486 ( .Y(n442), .A0(n430), .A1(n431) );
  nor02 U487 ( .Y(n443), .A0(n429), .A1(n431) );
  nor02 U488 ( .Y(n444), .A0(n429), .A1(n430) );
  nor02 U489 ( .Y(n428), .A0(n444), .A1(n445) );
  nor02 U490 ( .Y(n446), .A0(A[5]), .A1(carry_5_) );
  inv01 U491 ( .Y(n433), .A(n446) );
  nor02 U492 ( .Y(n447), .A0(B_not[5]), .A1(carry_5_) );
  inv01 U493 ( .Y(n435), .A(n447) );
  nor02 U494 ( .Y(n448), .A0(B_not[5]), .A1(A[5]) );
  inv01 U495 ( .Y(n437), .A(n448) );
  nor02 U496 ( .Y(n449), .A0(n429), .A1(n430) );
  inv01 U497 ( .Y(n439), .A(n449) );
  nor02 U498 ( .Y(n450), .A0(n432), .A1(n434) );
  inv01 U499 ( .Y(n440), .A(n450) );
  nor02 U500 ( .Y(n451), .A0(n436), .A1(n438) );
  inv01 U501 ( .Y(n441), .A(n451) );
  nor02 U502 ( .Y(n452), .A0(n442), .A1(n443) );
  inv01 U503 ( .Y(n445), .A(n452) );
  inv02 U504 ( .Y(B_not[5]), .A(B[5]) );
  inv01 U505 ( .Y(DIFF[4]), .A(n453) );
  inv02 U506 ( .Y(carry_5_), .A(n454) );
  inv02 U507 ( .Y(n455), .A(B_not[4]) );
  inv02 U508 ( .Y(n456), .A(A[4]) );
  inv02 U509 ( .Y(n457), .A(carry_4_) );
  nor02 U510 ( .Y(n458), .A0(n455), .A1(n459) );
  nor02 U511 ( .Y(n460), .A0(n456), .A1(n461) );
  nor02 U512 ( .Y(n462), .A0(n457), .A1(n463) );
  nor02 U513 ( .Y(n464), .A0(n457), .A1(n465) );
  nor02 U514 ( .Y(n453), .A0(n466), .A1(n467) );
  nor02 U515 ( .Y(n468), .A0(n456), .A1(n457) );
  nor02 U516 ( .Y(n469), .A0(n455), .A1(n457) );
  nor02 U517 ( .Y(n470), .A0(n455), .A1(n456) );
  nor02 U518 ( .Y(n454), .A0(n470), .A1(n471) );
  nor02 U519 ( .Y(n472), .A0(A[4]), .A1(carry_4_) );
  inv01 U520 ( .Y(n459), .A(n472) );
  nor02 U521 ( .Y(n473), .A0(B_not[4]), .A1(carry_4_) );
  inv01 U522 ( .Y(n461), .A(n473) );
  nor02 U523 ( .Y(n474), .A0(B_not[4]), .A1(A[4]) );
  inv01 U524 ( .Y(n463), .A(n474) );
  nor02 U525 ( .Y(n475), .A0(n455), .A1(n456) );
  inv01 U526 ( .Y(n465), .A(n475) );
  nor02 U527 ( .Y(n476), .A0(n458), .A1(n460) );
  inv01 U528 ( .Y(n466), .A(n476) );
  nor02 U529 ( .Y(n477), .A0(n462), .A1(n464) );
  inv01 U530 ( .Y(n467), .A(n477) );
  nor02 U531 ( .Y(n478), .A0(n468), .A1(n469) );
  inv01 U532 ( .Y(n471), .A(n478) );
  inv02 U533 ( .Y(B_not[4]), .A(B[4]) );
  inv01 U534 ( .Y(DIFF[3]), .A(n479) );
  inv02 U535 ( .Y(carry_4_), .A(n480) );
  inv02 U536 ( .Y(n481), .A(B_not[3]) );
  inv02 U537 ( .Y(n482), .A(A[3]) );
  inv02 U538 ( .Y(n483), .A(carry_3_) );
  nor02 U539 ( .Y(n484), .A0(n481), .A1(n485) );
  nor02 U540 ( .Y(n486), .A0(n482), .A1(n487) );
  nor02 U541 ( .Y(n488), .A0(n483), .A1(n489) );
  nor02 U542 ( .Y(n490), .A0(n483), .A1(n491) );
  nor02 U543 ( .Y(n479), .A0(n492), .A1(n493) );
  nor02 U544 ( .Y(n494), .A0(n482), .A1(n483) );
  nor02 U545 ( .Y(n495), .A0(n481), .A1(n483) );
  nor02 U546 ( .Y(n496), .A0(n481), .A1(n482) );
  nor02 U547 ( .Y(n480), .A0(n496), .A1(n497) );
  nor02 U548 ( .Y(n498), .A0(A[3]), .A1(carry_3_) );
  inv01 U549 ( .Y(n485), .A(n498) );
  nor02 U550 ( .Y(n499), .A0(B_not[3]), .A1(carry_3_) );
  inv01 U551 ( .Y(n487), .A(n499) );
  nor02 U552 ( .Y(n500), .A0(B_not[3]), .A1(A[3]) );
  inv01 U553 ( .Y(n489), .A(n500) );
  nor02 U554 ( .Y(n501), .A0(n481), .A1(n482) );
  inv01 U555 ( .Y(n491), .A(n501) );
  nor02 U556 ( .Y(n502), .A0(n484), .A1(n486) );
  inv01 U557 ( .Y(n492), .A(n502) );
  nor02 U558 ( .Y(n503), .A0(n488), .A1(n490) );
  inv01 U559 ( .Y(n493), .A(n503) );
  nor02 U560 ( .Y(n504), .A0(n494), .A1(n495) );
  inv01 U561 ( .Y(n497), .A(n504) );
  inv02 U562 ( .Y(B_not[3]), .A(B[3]) );
  inv01 U563 ( .Y(DIFF[2]), .A(n505) );
  inv02 U564 ( .Y(carry_3_), .A(n506) );
  inv02 U565 ( .Y(n507), .A(B_not[2]) );
  inv02 U566 ( .Y(n508), .A(A[2]) );
  inv02 U567 ( .Y(n509), .A(n531) );
  nor02 U568 ( .Y(n510), .A0(n507), .A1(n511) );
  nor02 U569 ( .Y(n512), .A0(n508), .A1(n513) );
  nor02 U570 ( .Y(n514), .A0(n509), .A1(n515) );
  nor02 U571 ( .Y(n516), .A0(n509), .A1(n517) );
  nor02 U572 ( .Y(n505), .A0(n518), .A1(n519) );
  nor02 U573 ( .Y(n520), .A0(n508), .A1(n509) );
  nor02 U574 ( .Y(n521), .A0(n507), .A1(n509) );
  nor02 U575 ( .Y(n522), .A0(n507), .A1(n508) );
  nor02 U576 ( .Y(n506), .A0(n522), .A1(n523) );
  nor02 U577 ( .Y(n524), .A0(A[2]), .A1(n531) );
  inv01 U578 ( .Y(n511), .A(n524) );
  nor02 U579 ( .Y(n525), .A0(B_not[2]), .A1(n531) );
  inv01 U580 ( .Y(n513), .A(n525) );
  nor02 U581 ( .Y(n526), .A0(B_not[2]), .A1(A[2]) );
  inv01 U582 ( .Y(n515), .A(n526) );
  nor02 U583 ( .Y(n527), .A0(n507), .A1(n508) );
  inv01 U584 ( .Y(n517), .A(n527) );
  nor02 U585 ( .Y(n528), .A0(n510), .A1(n512) );
  inv01 U586 ( .Y(n518), .A(n528) );
  nor02 U587 ( .Y(n529), .A0(n514), .A1(n516) );
  inv01 U588 ( .Y(n519), .A(n529) );
  nor02 U589 ( .Y(n530), .A0(n520), .A1(n521) );
  inv01 U590 ( .Y(n523), .A(n530) );
  inv02 U591 ( .Y(B_not[2]), .A(B[2]) );
  buf02 U592 ( .Y(n531), .A(carry_2_) );
  xnor2 U593 ( .Y(DIFF[0]), .A0(B_not[0]), .A1(A[0]) );
  inv04 U594 ( .Y(B_not[26]), .A(B[26]) );
  inv04 U595 ( .Y(B_not[25]), .A(B[25]) );
  inv04 U596 ( .Y(B_not[23]), .A(B[23]) );
  inv04 U597 ( .Y(B_not[22]), .A(B[22]) );
  inv04 U598 ( .Y(B_not[21]), .A(B[21]) );
  inv04 U599 ( .Y(B_not[1]), .A(B[1]) );
  inv04 U600 ( .Y(B_not[0]), .A(B[0]) );
  fadd1 U2_1 ( .S(DIFF[1]), .CO(carry_2_), .A(A[1]), .B(B_not[1]), .CI(n6) );
  fadd1 U2_21 ( .S(DIFF[21]), .CO(carry_22_), .A(A[21]), .B(B_not[21]), .CI(
        carry_21_) );
  fadd1 U2_22 ( .S(DIFF[22]), .CO(carry_23_), .A(A[22]), .B(B_not[22]), .CI(
        n36) );
  fadd1 U2_23 ( .S(DIFF[23]), .CO(carry_24_), .A(A[23]), .B(B_not[23]), .CI(
        n35) );
  fadd1 U2_25 ( .S(DIFF[25]), .CO(carry_26_), .A(A[25]), .B(B_not[25]), .CI(
        carry_25_) );
  fadd1 U2_26 ( .S(DIFF[26]), .A(A[26]), .B(B_not[26]), .CI(n7) );
endmodule


module serial_div_DW01_cmp2_27_0 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [26:0] A;
  input [26:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163;

  aoi21 U6 ( .Y(n15), .A0(B[26]), .A1(n97), .B0(n98) );
  inv01 U7 ( .Y(LT_LE), .A(n15) );
  nand02 U8 ( .Y(n159), .A0(n162), .A1(n17) );
  inv01 U9 ( .Y(n18), .A(n161) );
  inv01 U10 ( .Y(n19), .A(n160) );
  inv01 U11 ( .Y(n20), .A(B[2]) );
  inv01 U12 ( .Y(n21), .A(n157) );
  nand02 U13 ( .Y(n22), .A0(n18), .A1(n19) );
  nand02 U14 ( .Y(n23), .A0(n20), .A1(n21) );
  nand02 U15 ( .Y(n24), .A0(n22), .A1(n23) );
  inv01 U16 ( .Y(n17), .A(n24) );
  inv01 U17 ( .Y(n158), .A(n159) );
  inv01 U18 ( .Y(n114), .A(n25) );
  nor02 U19 ( .Y(n26), .A0(n115), .A1(B[19]) );
  nor02 U20 ( .Y(n27), .A0(n112), .A1(B[20]) );
  inv01 U21 ( .Y(n28), .A(n116) );
  nor02 U22 ( .Y(n25), .A0(n28), .A1(n29) );
  nor02 U23 ( .Y(n30), .A0(n26), .A1(n27) );
  inv01 U24 ( .Y(n29), .A(n30) );
  inv01 U25 ( .Y(n124), .A(n31) );
  nor02 U26 ( .Y(n32), .A0(n125), .A1(B[15]) );
  nor02 U27 ( .Y(n33), .A0(n122), .A1(B[16]) );
  inv01 U28 ( .Y(n34), .A(n126) );
  nor02 U29 ( .Y(n31), .A0(n34), .A1(n35) );
  nor02 U30 ( .Y(n36), .A0(n32), .A1(n33) );
  inv01 U31 ( .Y(n35), .A(n36) );
  inv01 U32 ( .Y(n113), .A(n114) );
  inv01 U33 ( .Y(n123), .A(n124) );
  inv01 U34 ( .Y(n104), .A(n37) );
  nor02 U35 ( .Y(n38), .A0(n105), .A1(B[23]) );
  nor02 U36 ( .Y(n39), .A0(n102), .A1(B[24]) );
  inv01 U37 ( .Y(n40), .A(n106) );
  nor02 U38 ( .Y(n37), .A0(n40), .A1(n41) );
  nor02 U39 ( .Y(n42), .A0(n38), .A1(n39) );
  inv01 U40 ( .Y(n41), .A(n42) );
  inv01 U41 ( .Y(n109), .A(n43) );
  nor02 U42 ( .Y(n44), .A0(n110), .A1(B[21]) );
  nor02 U43 ( .Y(n45), .A0(n107), .A1(B[22]) );
  inv01 U44 ( .Y(n46), .A(n111) );
  nor02 U45 ( .Y(n43), .A0(n46), .A1(n47) );
  nor02 U46 ( .Y(n48), .A0(n44), .A1(n45) );
  inv01 U47 ( .Y(n47), .A(n48) );
  inv01 U48 ( .Y(n103), .A(n104) );
  inv01 U49 ( .Y(n108), .A(n109) );
  inv01 U50 ( .Y(n139), .A(n49) );
  nor02 U51 ( .Y(n50), .A0(n137), .A1(B[10]) );
  nor02 U52 ( .Y(n51), .A0(n140), .A1(B[9]) );
  inv01 U53 ( .Y(n52), .A(n141) );
  nor02 U54 ( .Y(n49), .A0(n52), .A1(n53) );
  nor02 U55 ( .Y(n54), .A0(n50), .A1(n51) );
  inv01 U56 ( .Y(n53), .A(n54) );
  inv01 U57 ( .Y(n138), .A(n139) );
  inv01 U58 ( .Y(n119), .A(n55) );
  nor02 U59 ( .Y(n56), .A0(n120), .A1(B[17]) );
  nor02 U60 ( .Y(n57), .A0(n117), .A1(B[18]) );
  inv01 U61 ( .Y(n58), .A(n121) );
  nor02 U62 ( .Y(n55), .A0(n58), .A1(n59) );
  nor02 U63 ( .Y(n60), .A0(n56), .A1(n57) );
  inv01 U64 ( .Y(n59), .A(n60) );
  inv01 U65 ( .Y(n144), .A(n61) );
  nor02 U66 ( .Y(n62), .A0(n145), .A1(B[7]) );
  nor02 U67 ( .Y(n63), .A0(n142), .A1(B[8]) );
  inv01 U68 ( .Y(n64), .A(n146) );
  nor02 U69 ( .Y(n61), .A0(n64), .A1(n65) );
  nor02 U70 ( .Y(n66), .A0(n62), .A1(n63) );
  inv01 U71 ( .Y(n65), .A(n66) );
  inv01 U72 ( .Y(n118), .A(n119) );
  inv01 U73 ( .Y(n143), .A(n144) );
  inv01 U74 ( .Y(n149), .A(n67) );
  nor02 U75 ( .Y(n68), .A0(n150), .A1(B[5]) );
  nor02 U76 ( .Y(n69), .A0(n147), .A1(B[6]) );
  inv01 U77 ( .Y(n70), .A(n151) );
  nor02 U78 ( .Y(n67), .A0(n70), .A1(n71) );
  nor02 U79 ( .Y(n72), .A0(n68), .A1(n69) );
  inv01 U80 ( .Y(n71), .A(n72) );
  inv01 U81 ( .Y(n134), .A(n73) );
  nor02 U82 ( .Y(n74), .A0(n135), .A1(B[11]) );
  nor02 U83 ( .Y(n75), .A0(n132), .A1(B[12]) );
  inv01 U84 ( .Y(n76), .A(n136) );
  nor02 U85 ( .Y(n73), .A0(n76), .A1(n77) );
  nor02 U86 ( .Y(n78), .A0(n74), .A1(n75) );
  inv01 U87 ( .Y(n77), .A(n78) );
  inv01 U88 ( .Y(n148), .A(n149) );
  inv01 U89 ( .Y(n133), .A(n134) );
  inv01 U90 ( .Y(n154), .A(n79) );
  nor02 U91 ( .Y(n80), .A0(n155), .A1(B[3]) );
  nor02 U92 ( .Y(n81), .A0(n152), .A1(B[4]) );
  inv01 U93 ( .Y(n82), .A(n156) );
  nor02 U94 ( .Y(n79), .A0(n82), .A1(n83) );
  nor02 U95 ( .Y(n84), .A0(n80), .A1(n81) );
  inv01 U96 ( .Y(n83), .A(n84) );
  inv01 U97 ( .Y(n129), .A(n85) );
  nor02 U98 ( .Y(n86), .A0(n130), .A1(B[13]) );
  nor02 U99 ( .Y(n87), .A0(n127), .A1(B[14]) );
  inv01 U100 ( .Y(n88), .A(n131) );
  nor02 U101 ( .Y(n85), .A0(n88), .A1(n89) );
  nor02 U102 ( .Y(n90), .A0(n86), .A1(n87) );
  inv01 U103 ( .Y(n89), .A(n90) );
  inv01 U104 ( .Y(n153), .A(n154) );
  inv01 U105 ( .Y(n128), .A(n129) );
  inv01 U106 ( .Y(n99), .A(n91) );
  nor02 U107 ( .Y(n92), .A0(n100), .A1(B[25]) );
  nor02 U108 ( .Y(n93), .A0(n97), .A1(B[26]) );
  inv01 U109 ( .Y(n94), .A(n101) );
  nor02 U110 ( .Y(n91), .A0(n94), .A1(n95) );
  nor02 U111 ( .Y(n96), .A0(n92), .A1(n93) );
  inv01 U112 ( .Y(n95), .A(n96) );
  inv01 U113 ( .Y(n98), .A(n99) );
  inv02 U114 ( .Y(n100), .A(A[25]) );
  inv02 U115 ( .Y(n102), .A(A[24]) );
  inv02 U116 ( .Y(n155), .A(A[3]) );
  inv02 U117 ( .Y(n125), .A(A[15]) );
  inv02 U118 ( .Y(n130), .A(A[13]) );
  inv02 U119 ( .Y(n142), .A(A[8]) );
  inv02 U120 ( .Y(n117), .A(A[18]) );
  inv02 U121 ( .Y(n157), .A(A[2]) );
  inv02 U122 ( .Y(n135), .A(A[11]) );
  inv02 U123 ( .Y(n107), .A(A[22]) );
  inv02 U124 ( .Y(n160), .A(A[1]) );
  inv02 U125 ( .Y(n147), .A(A[6]) );
  inv02 U126 ( .Y(n112), .A(A[20]) );
  inv02 U127 ( .Y(n110), .A(A[21]) );
  inv02 U128 ( .Y(n115), .A(A[19]) );
  inv02 U129 ( .Y(n120), .A(A[17]) );
  inv02 U130 ( .Y(n140), .A(A[9]) );
  inv02 U131 ( .Y(n105), .A(A[23]) );
  inv02 U132 ( .Y(n145), .A(A[7]) );
  inv02 U133 ( .Y(n132), .A(A[12]) );
  inv02 U134 ( .Y(n122), .A(A[16]) );
  inv02 U135 ( .Y(n127), .A(A[14]) );
  inv02 U136 ( .Y(n150), .A(A[5]) );
  inv02 U137 ( .Y(n152), .A(A[4]) );
  inv02 U138 ( .Y(n137), .A(A[10]) );
  inv02 U139 ( .Y(n97), .A(A[26]) );
  inv04 U140 ( .Y(n163), .A(B[0]) );
  ao221 U141 ( .Y(n101), .A0(B[25]), .A1(n100), .B0(B[24]), .B1(n102), .C0(
        n103) );
  ao221 U142 ( .Y(n106), .A0(B[23]), .A1(n105), .B0(B[22]), .B1(n107), .C0(
        n108) );
  ao221 U143 ( .Y(n111), .A0(B[21]), .A1(n110), .B0(B[20]), .B1(n112), .C0(
        n113) );
  ao221 U144 ( .Y(n116), .A0(B[19]), .A1(n115), .B0(B[18]), .B1(n117), .C0(
        n118) );
  ao221 U145 ( .Y(n121), .A0(B[17]), .A1(n120), .B0(B[16]), .B1(n122), .C0(
        n123) );
  ao221 U146 ( .Y(n126), .A0(B[15]), .A1(n125), .B0(B[14]), .B1(n127), .C0(
        n128) );
  ao221 U147 ( .Y(n131), .A0(B[13]), .A1(n130), .B0(B[12]), .B1(n132), .C0(
        n133) );
  ao221 U148 ( .Y(n136), .A0(B[11]), .A1(n135), .B0(B[10]), .B1(n137), .C0(
        n138) );
  ao221 U149 ( .Y(n141), .A0(B[9]), .A1(n140), .B0(B[8]), .B1(n142), .C0(n143)
         );
  ao221 U150 ( .Y(n146), .A0(B[7]), .A1(n145), .B0(B[6]), .B1(n147), .C0(n148)
         );
  ao221 U151 ( .Y(n151), .A0(B[5]), .A1(n150), .B0(B[4]), .B1(n152), .C0(n153)
         );
  ao221 U152 ( .Y(n156), .A0(B[3]), .A1(n155), .B0(B[2]), .B1(n157), .C0(n158)
         );
  ao21 U153 ( .Y(n162), .A0(n161), .A1(n160), .B0(B[1]) );
  nor02 U154 ( .Y(n161), .A0(n163), .A1(A[0]) );
endmodule


module serial_div_DW01_dec_5_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   carry_4_, carry_3_, n5, n7, n9, n11, n13, n14, n15;

  xor2 U6 ( .Y(n5), .A0(carry_4_), .A1(A[4]) );
  inv01 U7 ( .Y(SUM[4]), .A(n5) );
  xor2 U8 ( .Y(n7), .A0(A[3]), .A1(n15) );
  inv01 U9 ( .Y(SUM[3]), .A(n7) );
  xor2 U10 ( .Y(n9), .A0(A[1]), .A1(A[0]) );
  inv01 U11 ( .Y(SUM[1]), .A(n9) );
  xor2 U12 ( .Y(n11), .A0(A[2]), .A1(n14) );
  inv01 U13 ( .Y(SUM[2]), .A(n11) );
  nor02 U14 ( .Y(n13), .A0(A[1]), .A1(A[0]) );
  inv02 U15 ( .Y(n14), .A(n13) );
  buf02 U16 ( .Y(n15), .A(carry_3_) );
  inv01 U17 ( .Y(SUM[0]), .A(A[0]) );
  or02 U1_B_2 ( .Y(carry_3_), .A0(A[2]), .A1(n14) );
  or02 U1_B_3 ( .Y(carry_4_), .A0(A[3]), .A1(n15) );
endmodule


module serial_div ( clk_i, dvdnd_i, dvsor_i, sign_dvd_i, sign_div_i, start_i, 
        ready_o, qutnt_o, rmndr_o, sign_o, div_zero_o );
  input [49:0] dvdnd_i;
  input [26:0] dvsor_i;
  output [26:0] qutnt_o;
  output [26:0] rmndr_o;
  input clk_i, sign_dvd_i, sign_div_i, start_i;
  output ready_o, sign_o, div_zero_o;
  wire   s_dvdnd_i_49_, s_dvdnd_i_48_, s_dvdnd_i_47_, s_dvdnd_i_46_,
         s_dvdnd_i_45_, s_dvdnd_i_44_, s_dvdnd_i_43_, s_dvdnd_i_42_,
         s_dvdnd_i_41_, s_dvdnd_i_40_, s_dvdnd_i_39_, s_dvdnd_i_38_,
         s_dvdnd_i_37_, s_dvdnd_i_36_, s_dvdnd_i_35_, s_dvdnd_i_34_,
         s_dvdnd_i_33_, s_dvdnd_i_32_, s_dvdnd_i_31_, s_dvdnd_i_30_,
         s_dvdnd_i_29_, s_dvdnd_i_28_, s_dvdnd_i_27_, s_dvdnd_i_26_,
         s_dvdnd_i_25_, s_dvdnd_i_14_, s_dvdnd_i_5_, s_dvdnd_i_4_,
         s_dvsor_i_26_, s_dvsor_i_25_, s_dvsor_i_24_, s_dvsor_i_23_,
         s_dvsor_i_22_, s_dvsor_i_21_, s_dvsor_i_20_, s_dvsor_i_19_,
         s_dvsor_i_18_, s_dvsor_i_17_, s_dvsor_i_16_, s_dvsor_i_15_,
         s_dvsor_i_14_, s_dvsor_i_13_, s_dvsor_i_12_, s_dvsor_i_11_,
         s_dvsor_i_10_, s_dvsor_i_9_, s_dvsor_i_8_, s_dvsor_i_7_, s_dvsor_i_6_,
         s_dvsor_i_5_, s_dvsor_i_4_, s_dvsor_i_3_, s_dvsor_i_2_, s_dvsor_i_1_,
         s_dvsor_i_0_, s_state, s_state355, sum426_4_, sum426_3_, sum426_2_,
         sum426_1_, sum426_0_, n____return556, n____return927_26_,
         n____return927_25_, n____return927_24_, n____return927_23_,
         n____return927_22_, n____return927_21_, n____return927_20_,
         n____return927_19_, n____return927_18_, n____return927_17_,
         n____return927_16_, n____return927_15_, n____return927_14_,
         n____return927_13_, n____return927_12_, n____return927_11_,
         n____return927_10_, n____return927_9_, n____return927_8_,
         n____return927_7_, n____return927_6_, n____return927_5_,
         n____return927_4_, n____return927_3_, n____return927_2_,
         n____return927_1_, n____return927_0_, L546_26_, L546_25_, L546_24_,
         L546_23_, L546_22_, L546_21_, L546_20_, L546_19_, L546_18_, L546_17_,
         L546_16_, L546_15_, L546_14_, L546_13_, L546_12_, L546_11_, L546_10_,
         L546_9_, L546_8_, L546_7_, L546_6_, L546_5_, L546_4_, L546_3_,
         L546_2_, L546_1_, L546_0_, n1385, n1387, n1388, n1389, n1390, n1394,
         n1395, n1396, n1397, n1401, n1405, n1406, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589;
  wire   [4:0] s_count;
  wire   [26:0] s_dvd;

  dff s_count_reg_0_ ( .Q(s_count[0]), .QB(n2286), .D(n1681), .CLK(clk_i) );
  dff s_count_reg_1_ ( .Q(s_count[1]), .D(n1682), .CLK(clk_i) );
  dff s_count_reg_2_ ( .Q(s_count[2]), .D(n1683), .CLK(clk_i) );
  dff s_count_reg_3_ ( .Q(s_count[3]), .D(n1684), .CLK(clk_i) );
  dff s_count_reg_4_ ( .Q(s_count[4]), .D(n1685), .CLK(clk_i) );
  dff s_qutnt_o_reg_26_ ( .Q(qutnt_o[26]), .QB(n2550), .D(n1686), .CLK(clk_i)
         );
  dff s_qutnt_o_reg_25_ ( .Q(qutnt_o[25]), .QB(n2551), .D(n1687), .CLK(clk_i)
         );
  dff s_qutnt_o_reg_24_ ( .Q(qutnt_o[24]), .QB(n2552), .D(n1688), .CLK(clk_i)
         );
  dff s_qutnt_o_reg_23_ ( .Q(qutnt_o[23]), .QB(n2553), .D(n1689), .CLK(clk_i)
         );
  dff s_qutnt_o_reg_22_ ( .Q(qutnt_o[22]), .QB(n2554), .D(n1690), .CLK(clk_i)
         );
  dff s_qutnt_o_reg_21_ ( .Q(qutnt_o[21]), .QB(n2555), .D(n1691), .CLK(clk_i)
         );
  dff s_qutnt_o_reg_20_ ( .Q(qutnt_o[20]), .QB(n2556), .D(n1692), .CLK(clk_i)
         );
  dff s_qutnt_o_reg_19_ ( .Q(qutnt_o[19]), .QB(n2558), .D(n1693), .CLK(clk_i)
         );
  dff s_qutnt_o_reg_18_ ( .Q(qutnt_o[18]), .QB(n2559), .D(n1694), .CLK(clk_i)
         );
  dff s_qutnt_o_reg_17_ ( .Q(qutnt_o[17]), .QB(n2560), .D(n1695), .CLK(clk_i)
         );
  dff s_qutnt_o_reg_16_ ( .Q(qutnt_o[16]), .QB(n2561), .D(n1696), .CLK(clk_i)
         );
  dff s_qutnt_o_reg_15_ ( .Q(qutnt_o[15]), .QB(n2562), .D(n1697), .CLK(clk_i)
         );
  dff s_qutnt_o_reg_14_ ( .Q(qutnt_o[14]), .QB(n2563), .D(n1698), .CLK(clk_i)
         );
  dff s_qutnt_o_reg_13_ ( .Q(qutnt_o[13]), .QB(n2564), .D(n1699), .CLK(clk_i)
         );
  dff s_qutnt_o_reg_12_ ( .Q(qutnt_o[12]), .QB(n2565), .D(n1700), .CLK(clk_i)
         );
  dff s_qutnt_o_reg_11_ ( .Q(qutnt_o[11]), .QB(n2566), .D(n1701), .CLK(clk_i)
         );
  dff s_qutnt_o_reg_10_ ( .Q(qutnt_o[10]), .QB(n2567), .D(n1702), .CLK(clk_i)
         );
  dff s_qutnt_o_reg_9_ ( .Q(qutnt_o[9]), .QB(n2542), .D(n1703), .CLK(clk_i) );
  dff s_qutnt_o_reg_8_ ( .Q(qutnt_o[8]), .QB(n2543), .D(n1704), .CLK(clk_i) );
  dff s_qutnt_o_reg_7_ ( .Q(qutnt_o[7]), .QB(n2544), .D(n1705), .CLK(clk_i) );
  dff s_qutnt_o_reg_6_ ( .Q(qutnt_o[6]), .QB(n2545), .D(n1706), .CLK(clk_i) );
  dff s_qutnt_o_reg_5_ ( .Q(qutnt_o[5]), .QB(n2546), .D(n1707), .CLK(clk_i) );
  dff s_qutnt_o_reg_4_ ( .Q(qutnt_o[4]), .QB(n2547), .D(n1708), .CLK(clk_i) );
  dff s_qutnt_o_reg_3_ ( .Q(qutnt_o[3]), .QB(n2548), .D(n1709), .CLK(clk_i) );
  dff s_qutnt_o_reg_2_ ( .Q(qutnt_o[2]), .QB(n2549), .D(n1710), .CLK(clk_i) );
  dff s_qutnt_o_reg_1_ ( .Q(qutnt_o[1]), .QB(n2557), .D(n1711), .CLK(clk_i) );
  dff s_qutnt_o_reg_0_ ( .Q(qutnt_o[0]), .QB(n2568), .D(n1712), .CLK(clk_i) );
  dff s_rmndr_o_reg_26_ ( .Q(rmndr_o[26]), .QB(n2541), .D(n1713), .CLK(clk_i)
         );
  dff s_rmndr_o_reg_25_ ( .Q(rmndr_o[25]), .QB(n1672), .D(n1714), .CLK(clk_i)
         );
  dff s_rmndr_o_reg_24_ ( .Q(rmndr_o[24]), .QB(n1671), .D(n1715), .CLK(clk_i)
         );
  dff s_rmndr_o_reg_23_ ( .Q(rmndr_o[23]), .QB(n1670), .D(n1716), .CLK(clk_i)
         );
  dff s_rmndr_o_reg_22_ ( .Q(rmndr_o[22]), .QB(n1669), .D(n1717), .CLK(clk_i)
         );
  dff s_rmndr_o_reg_21_ ( .Q(rmndr_o[21]), .QB(n1668), .D(n1718), .CLK(clk_i)
         );
  dff s_rmndr_o_reg_20_ ( .Q(rmndr_o[20]), .QB(n1667), .D(n1719), .CLK(clk_i)
         );
  dff s_rmndr_o_reg_19_ ( .Q(rmndr_o[19]), .QB(n1665), .D(n1720), .CLK(clk_i)
         );
  dff s_rmndr_o_reg_18_ ( .Q(rmndr_o[18]), .QB(n1664), .D(n1721), .CLK(clk_i)
         );
  dff s_rmndr_o_reg_17_ ( .Q(rmndr_o[17]), .QB(n1663), .D(n1722), .CLK(clk_i)
         );
  dff s_rmndr_o_reg_16_ ( .Q(rmndr_o[16]), .QB(n1662), .D(n1723), .CLK(clk_i)
         );
  dff s_rmndr_o_reg_15_ ( .Q(rmndr_o[15]), .QB(n1661), .D(n1724), .CLK(clk_i)
         );
  dff s_rmndr_o_reg_14_ ( .Q(rmndr_o[14]), .QB(n1660), .D(n1725), .CLK(clk_i)
         );
  dff s_rmndr_o_reg_13_ ( .Q(rmndr_o[13]), .QB(n1659), .D(n1726), .CLK(clk_i)
         );
  dff s_rmndr_o_reg_12_ ( .Q(rmndr_o[12]), .QB(n1658), .D(n1727), .CLK(clk_i)
         );
  dff s_rmndr_o_reg_11_ ( .Q(rmndr_o[11]), .QB(n1657), .D(n1728), .CLK(clk_i)
         );
  dff s_rmndr_o_reg_10_ ( .Q(rmndr_o[10]), .QB(n1656), .D(n1729), .CLK(clk_i)
         );
  dff s_rmndr_o_reg_9_ ( .Q(rmndr_o[9]), .QB(n1680), .D(n1730), .CLK(clk_i) );
  dff s_rmndr_o_reg_8_ ( .Q(rmndr_o[8]), .QB(n1679), .D(n1731), .CLK(clk_i) );
  dff s_rmndr_o_reg_7_ ( .Q(rmndr_o[7]), .QB(n1678), .D(n1732), .CLK(clk_i) );
  dff s_rmndr_o_reg_6_ ( .Q(rmndr_o[6]), .QB(n1677), .D(n1733), .CLK(clk_i) );
  dff s_rmndr_o_reg_5_ ( .Q(rmndr_o[5]), .QB(n1676), .D(n1734), .CLK(clk_i) );
  dff s_rmndr_o_reg_4_ ( .Q(rmndr_o[4]), .QB(n1675), .D(n1735), .CLK(clk_i) );
  dff s_rmndr_o_reg_3_ ( .Q(rmndr_o[3]), .QB(n1674), .D(n1736), .CLK(clk_i) );
  dff s_rmndr_o_reg_2_ ( .Q(rmndr_o[2]), .QB(n1673), .D(n1737), .CLK(clk_i) );
  dff s_rmndr_o_reg_1_ ( .Q(rmndr_o[1]), .QB(n1666), .D(n1738), .CLK(clk_i) );
  dff s_rmndr_o_reg_0_ ( .Q(rmndr_o[0]), .QB(n1655), .D(n1739), .CLK(clk_i) );
  dff s_dvd_reg_26_ ( .Q(s_dvd[26]), .D(n1740), .CLK(clk_i) );
  dff s_dvd_reg_25_ ( .Q(s_dvd[25]), .D(n1741), .CLK(clk_i) );
  dff s_dvd_reg_24_ ( .Q(s_dvd[24]), .D(n1742), .CLK(clk_i) );
  dff s_dvd_reg_23_ ( .Q(s_dvd[23]), .D(n1743), .CLK(clk_i) );
  dff s_dvd_reg_22_ ( .Q(s_dvd[22]), .D(n1744), .CLK(clk_i) );
  dff s_dvd_reg_21_ ( .Q(s_dvd[21]), .D(n1745), .CLK(clk_i) );
  dff s_dvd_reg_20_ ( .Q(s_dvd[20]), .D(n1746), .CLK(clk_i) );
  dff s_dvd_reg_19_ ( .Q(s_dvd[19]), .D(n1747), .CLK(clk_i) );
  dff s_dvd_reg_18_ ( .Q(s_dvd[18]), .D(n1748), .CLK(clk_i) );
  dff s_dvd_reg_17_ ( .Q(s_dvd[17]), .D(n1749), .CLK(clk_i) );
  dff s_dvd_reg_16_ ( .Q(s_dvd[16]), .D(n1750), .CLK(clk_i) );
  dff s_dvd_reg_15_ ( .Q(s_dvd[15]), .D(n1751), .CLK(clk_i) );
  dff s_dvd_reg_14_ ( .Q(s_dvd[14]), .D(n1752), .CLK(clk_i) );
  dff s_dvd_reg_13_ ( .Q(s_dvd[13]), .D(n1753), .CLK(clk_i) );
  dff s_dvd_reg_12_ ( .Q(s_dvd[12]), .D(n1754), .CLK(clk_i) );
  dff s_dvd_reg_11_ ( .Q(s_dvd[11]), .D(n1755), .CLK(clk_i) );
  dff s_dvd_reg_10_ ( .Q(s_dvd[10]), .D(n1756), .CLK(clk_i) );
  dff s_dvd_reg_9_ ( .Q(s_dvd[9]), .D(n1757), .CLK(clk_i) );
  dff s_dvd_reg_8_ ( .Q(s_dvd[8]), .D(n1758), .CLK(clk_i) );
  dff s_dvd_reg_7_ ( .Q(s_dvd[7]), .D(n1759), .CLK(clk_i) );
  dff s_dvd_reg_6_ ( .Q(s_dvd[6]), .D(n1760), .CLK(clk_i) );
  dff s_dvd_reg_5_ ( .Q(s_dvd[5]), .D(n1761), .CLK(clk_i) );
  dff s_dvd_reg_4_ ( .Q(s_dvd[4]), .D(n1762), .CLK(clk_i) );
  dff s_dvd_reg_3_ ( .Q(s_dvd[3]), .D(n1763), .CLK(clk_i) );
  dff s_dvd_reg_2_ ( .Q(s_dvd[2]), .D(n1764), .CLK(clk_i) );
  dff s_dvd_reg_1_ ( .Q(s_dvd[1]), .D(n1765), .CLK(clk_i) );
  dff s_dvd_reg_0_ ( .Q(s_dvd[0]), .D(n1766), .CLK(clk_i) );
  dff s_state_reg ( .Q(s_state), .D(n1767), .CLK(clk_i) );
  dff s_ready_o_reg ( .Q(ready_o), .QB(n1654), .D(n1768), .CLK(clk_i) );
  dff s_dvdnd_i_reg_49_ ( .Q(s_dvdnd_i_49_), .D(dvdnd_i[49]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_48_ ( .Q(s_dvdnd_i_48_), .D(dvdnd_i[48]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_47_ ( .Q(s_dvdnd_i_47_), .D(dvdnd_i[47]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_46_ ( .Q(s_dvdnd_i_46_), .D(dvdnd_i[46]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_45_ ( .Q(s_dvdnd_i_45_), .D(dvdnd_i[45]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_44_ ( .Q(s_dvdnd_i_44_), .D(dvdnd_i[44]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_43_ ( .Q(s_dvdnd_i_43_), .D(dvdnd_i[43]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_42_ ( .Q(s_dvdnd_i_42_), .D(dvdnd_i[42]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_41_ ( .Q(s_dvdnd_i_41_), .D(dvdnd_i[41]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_40_ ( .Q(s_dvdnd_i_40_), .D(dvdnd_i[40]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_39_ ( .Q(s_dvdnd_i_39_), .D(dvdnd_i[39]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_38_ ( .Q(s_dvdnd_i_38_), .D(dvdnd_i[38]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_37_ ( .Q(s_dvdnd_i_37_), .D(dvdnd_i[37]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_36_ ( .Q(s_dvdnd_i_36_), .D(dvdnd_i[36]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_35_ ( .Q(s_dvdnd_i_35_), .D(dvdnd_i[35]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_34_ ( .Q(s_dvdnd_i_34_), .D(dvdnd_i[34]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_33_ ( .Q(s_dvdnd_i_33_), .D(dvdnd_i[33]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_32_ ( .Q(s_dvdnd_i_32_), .D(dvdnd_i[32]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_31_ ( .Q(s_dvdnd_i_31_), .D(dvdnd_i[31]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_30_ ( .Q(s_dvdnd_i_30_), .D(dvdnd_i[30]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_29_ ( .Q(s_dvdnd_i_29_), .D(dvdnd_i[29]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_28_ ( .Q(s_dvdnd_i_28_), .D(dvdnd_i[28]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_27_ ( .Q(s_dvdnd_i_27_), .D(dvdnd_i[27]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_26_ ( .Q(s_dvdnd_i_26_), .D(dvdnd_i[26]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_25_ ( .Q(s_dvdnd_i_25_), .D(dvdnd_i[25]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_24_ ( .QB(n2581), .D(dvdnd_i[24]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_23_ ( .QB(n2582), .D(dvdnd_i[23]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_22_ ( .QB(n2584), .D(dvdnd_i[22]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_21_ ( .QB(n2583), .D(dvdnd_i[21]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_20_ ( .QB(n2585), .D(dvdnd_i[20]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_19_ ( .QB(n2577), .D(dvdnd_i[19]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_18_ ( .QB(n2579), .D(dvdnd_i[18]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_17_ ( .QB(n1406), .D(dvdnd_i[17]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_16_ ( .QB(n1405), .D(dvdnd_i[16]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_15_ ( .Q(n2576), .D(dvdnd_i[15]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_14_ ( .Q(s_dvdnd_i_14_), .D(dvdnd_i[14]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_13_ ( .QB(n2574), .D(dvdnd_i[13]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_12_ ( .QB(n2575), .D(dvdnd_i[12]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_11_ ( .Q(n2572), .D(dvdnd_i[11]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_10_ ( .Q(n2573), .D(dvdnd_i[10]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_9_ ( .QB(n1401), .D(dvdnd_i[9]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_8_ ( .Q(n2586), .D(dvdnd_i[8]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_7_ ( .Q(n2587), .D(dvdnd_i[7]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_6_ ( .Q(n2588), .D(dvdnd_i[6]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_5_ ( .Q(s_dvdnd_i_5_), .D(dvdnd_i[5]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_4_ ( .Q(s_dvdnd_i_4_), .D(dvdnd_i[4]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_3_ ( .QB(n2589), .D(dvdnd_i[3]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_2_ ( .QB(n2580), .D(dvdnd_i[2]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_1_ ( .QB(n2578), .D(dvdnd_i[1]), .CLK(clk_i) );
  dff s_dvdnd_i_reg_0_ ( .QB(n1397), .D(dvdnd_i[0]), .CLK(clk_i) );
  dff s_dvsor_i_reg_26_ ( .Q(s_dvsor_i_26_), .D(dvsor_i[26]), .CLK(clk_i) );
  dff s_dvsor_i_reg_25_ ( .Q(s_dvsor_i_25_), .D(dvsor_i[25]), .CLK(clk_i) );
  dff s_dvsor_i_reg_24_ ( .Q(s_dvsor_i_24_), .D(dvsor_i[24]), .CLK(clk_i) );
  dff s_dvsor_i_reg_23_ ( .Q(s_dvsor_i_23_), .QB(n1396), .D(dvsor_i[23]), 
        .CLK(clk_i) );
  dff s_dvsor_i_reg_22_ ( .Q(s_dvsor_i_22_), .QB(n1395), .D(dvsor_i[22]), 
        .CLK(clk_i) );
  dff s_dvsor_i_reg_21_ ( .Q(s_dvsor_i_21_), .QB(n1394), .D(dvsor_i[21]), 
        .CLK(clk_i) );
  dff s_dvsor_i_reg_20_ ( .Q(s_dvsor_i_20_), .D(dvsor_i[20]), .CLK(clk_i) );
  dff s_dvsor_i_reg_19_ ( .Q(s_dvsor_i_19_), .D(dvsor_i[19]), .CLK(clk_i) );
  dff s_dvsor_i_reg_18_ ( .Q(s_dvsor_i_18_), .D(dvsor_i[18]), .CLK(clk_i) );
  dff s_dvsor_i_reg_17_ ( .Q(s_dvsor_i_17_), .QB(n2570), .D(dvsor_i[17]), 
        .CLK(clk_i) );
  dff s_dvsor_i_reg_16_ ( .Q(s_dvsor_i_16_), .QB(n2569), .D(dvsor_i[16]), 
        .CLK(clk_i) );
  dff s_dvsor_i_reg_15_ ( .Q(s_dvsor_i_15_), .QB(n2571), .D(dvsor_i[15]), 
        .CLK(clk_i) );
  dff s_dvsor_i_reg_14_ ( .Q(s_dvsor_i_14_), .D(dvsor_i[14]), .CLK(clk_i) );
  dff s_dvsor_i_reg_13_ ( .Q(s_dvsor_i_13_), .D(dvsor_i[13]), .CLK(clk_i) );
  dff s_dvsor_i_reg_12_ ( .Q(s_dvsor_i_12_), .D(dvsor_i[12]), .CLK(clk_i) );
  dff s_dvsor_i_reg_11_ ( .Q(s_dvsor_i_11_), .D(dvsor_i[11]), .CLK(clk_i) );
  dff s_dvsor_i_reg_10_ ( .Q(s_dvsor_i_10_), .QB(n1390), .D(dvsor_i[10]), 
        .CLK(clk_i) );
  dff s_dvsor_i_reg_9_ ( .Q(s_dvsor_i_9_), .D(dvsor_i[9]), .CLK(clk_i) );
  dff s_dvsor_i_reg_8_ ( .Q(s_dvsor_i_8_), .D(dvsor_i[8]), .CLK(clk_i) );
  dff s_dvsor_i_reg_7_ ( .Q(s_dvsor_i_7_), .D(dvsor_i[7]), .CLK(clk_i) );
  dff s_dvsor_i_reg_6_ ( .Q(s_dvsor_i_6_), .D(dvsor_i[6]), .CLK(clk_i) );
  dff s_dvsor_i_reg_5_ ( .Q(s_dvsor_i_5_), .QB(n1389), .D(dvsor_i[5]), .CLK(
        clk_i) );
  dff s_dvsor_i_reg_4_ ( .Q(s_dvsor_i_4_), .QB(n1388), .D(dvsor_i[4]), .CLK(
        clk_i) );
  dff s_dvsor_i_reg_3_ ( .Q(s_dvsor_i_3_), .QB(n1387), .D(dvsor_i[3]), .CLK(
        clk_i) );
  dff s_dvsor_i_reg_2_ ( .Q(s_dvsor_i_2_), .D(dvsor_i[2]), .CLK(clk_i) );
  dff s_dvsor_i_reg_1_ ( .Q(s_dvsor_i_1_), .D(dvsor_i[1]), .CLK(clk_i) );
  dff s_dvsor_i_reg_0_ ( .Q(s_dvsor_i_0_), .QB(n1385), .D(dvsor_i[0]), .CLK(
        clk_i) );
  dff s_start_i_reg ( .Q(s_state355), .D(start_i), .CLK(clk_i) );
  ao22 U587 ( .Y(n1769), .A0(L546_26_), .A1(n2269), .B0(n____return927_26_), 
        .B1(n2455) );
  inv01 U588 ( .Y(n1770), .A(n1769) );
  nand02 U589 ( .Y(n2515), .A0(n1771), .A1(n1772) );
  inv01 U590 ( .Y(n1773), .A(s_state) );
  inv01 U591 ( .Y(n1774), .A(n2389) );
  inv01 U592 ( .Y(n1775), .A(s_count[3]) );
  inv01 U593 ( .Y(n1776), .A(sum426_3_) );
  nand02 U594 ( .Y(n1777), .A0(n1773), .A1(n1774) );
  nand02 U595 ( .Y(n1778), .A0(n1773), .A1(n1775) );
  nand02 U596 ( .Y(n1779), .A0(n1774), .A1(n1776) );
  nand02 U597 ( .Y(n1780), .A0(n1775), .A1(n1776) );
  nand02 U598 ( .Y(n1781), .A0(n1777), .A1(n1778) );
  inv01 U599 ( .Y(n1771), .A(n1781) );
  nand02 U600 ( .Y(n1782), .A0(n1779), .A1(n1780) );
  inv01 U601 ( .Y(n1772), .A(n1782) );
  nand02 U602 ( .Y(n2514), .A0(n1783), .A1(n1784) );
  inv01 U603 ( .Y(n1785), .A(s_state) );
  inv01 U604 ( .Y(n1786), .A(n2389) );
  inv01 U605 ( .Y(n1787), .A(s_count[4]) );
  inv01 U606 ( .Y(n1788), .A(sum426_4_) );
  nand02 U607 ( .Y(n1789), .A0(n1785), .A1(n1786) );
  nand02 U608 ( .Y(n1790), .A0(n1785), .A1(n1787) );
  nand02 U609 ( .Y(n1791), .A0(n1786), .A1(n1788) );
  nand02 U610 ( .Y(n1792), .A0(n1787), .A1(n1788) );
  nand02 U611 ( .Y(n1793), .A0(n1789), .A1(n1790) );
  inv01 U612 ( .Y(n1783), .A(n1793) );
  nand02 U613 ( .Y(n1794), .A0(n1791), .A1(n1792) );
  inv01 U614 ( .Y(n1784), .A(n1794) );
  nand02 U615 ( .Y(n2517), .A0(n1795), .A1(n1796) );
  inv01 U616 ( .Y(n1797), .A(s_state) );
  inv01 U617 ( .Y(n1798), .A(n2389) );
  inv01 U618 ( .Y(n1799), .A(s_count[1]) );
  inv01 U619 ( .Y(n1800), .A(sum426_1_) );
  nand02 U620 ( .Y(n1801), .A0(n1797), .A1(n1798) );
  nand02 U621 ( .Y(n1802), .A0(n1797), .A1(n1799) );
  nand02 U622 ( .Y(n1803), .A0(n1798), .A1(n1800) );
  nand02 U623 ( .Y(n1804), .A0(n1799), .A1(n1800) );
  nand02 U624 ( .Y(n1805), .A0(n1801), .A1(n1802) );
  inv01 U625 ( .Y(n1795), .A(n1805) );
  nand02 U626 ( .Y(n1806), .A0(n1803), .A1(n1804) );
  inv01 U627 ( .Y(n1796), .A(n1806) );
  buf02 U628 ( .Y(n1807), .A(n2524) );
  inv01 U629 ( .Y(n2516), .A(n1808) );
  nor02 U630 ( .Y(n1809), .A0(n1904), .A1(n2393) );
  nor02 U631 ( .Y(n1810), .A0(s_state355), .A1(n2499) );
  nor02 U632 ( .Y(n1808), .A0(n1809), .A1(n1810) );
  inv01 U633 ( .Y(n1709), .A(n1811) );
  nor02 U634 ( .Y(n1812), .A0(n2381), .A1(n1905) );
  inv01 U635 ( .Y(n1813), .A(n2466) );
  nor02 U636 ( .Y(n1811), .A0(n1812), .A1(n1813) );
  inv01 U637 ( .Y(n1707), .A(n1814) );
  nor02 U638 ( .Y(n1815), .A0(n2381), .A1(n2469) );
  inv01 U639 ( .Y(n1816), .A(n2470) );
  nor02 U640 ( .Y(n1814), .A0(n1815), .A1(n1816) );
  inv01 U641 ( .Y(n1705), .A(n1817) );
  nor02 U642 ( .Y(n1818), .A0(n2381), .A1(n2235) );
  inv01 U643 ( .Y(n1819), .A(n2476) );
  nor02 U644 ( .Y(n1817), .A0(n1818), .A1(n1819) );
  inv01 U645 ( .Y(n1708), .A(n1820) );
  nor02 U646 ( .Y(n1821), .A0(n2381), .A1(n2467) );
  inv01 U647 ( .Y(n1822), .A(n2468) );
  nor02 U648 ( .Y(n1820), .A0(n1821), .A1(n1822) );
  inv01 U649 ( .Y(n1712), .A(n1823) );
  nor02 U650 ( .Y(n1824), .A0(n2381), .A1(n2285) );
  inv01 U651 ( .Y(n1825), .A(n2458) );
  nor02 U652 ( .Y(n1823), .A0(n1824), .A1(n1825) );
  inv01 U653 ( .Y(n1710), .A(n1826) );
  nor02 U654 ( .Y(n1827), .A0(n2381), .A1(n1902) );
  inv01 U655 ( .Y(n1828), .A(n2464) );
  nor02 U656 ( .Y(n1826), .A0(n1827), .A1(n1828) );
  inv01 U657 ( .Y(n1706), .A(n1829) );
  nor02 U658 ( .Y(n1830), .A0(n2381), .A1(n2236) );
  inv01 U659 ( .Y(n1831), .A(n2472) );
  nor02 U660 ( .Y(n1829), .A0(n1830), .A1(n1831) );
  inv01 U661 ( .Y(n1687), .A(n1832) );
  nor02 U662 ( .Y(n1833), .A0(n2280), .A1(n2284) );
  inv01 U663 ( .Y(n1834), .A(n2510) );
  nor02 U664 ( .Y(n1832), .A0(n1833), .A1(n1834) );
  inv01 U665 ( .Y(n1697), .A(n1835) );
  nor02 U666 ( .Y(n1836), .A0(n2235), .A1(n2379) );
  inv01 U667 ( .Y(n1837), .A(n2485) );
  nor02 U668 ( .Y(n1835), .A0(n1836), .A1(n1837) );
  inv01 U669 ( .Y(n1698), .A(n1838) );
  nor02 U670 ( .Y(n1839), .A0(n2236), .A1(n2379) );
  inv01 U671 ( .Y(n1840), .A(n2484) );
  nor02 U672 ( .Y(n1838), .A0(n1839), .A1(n1840) );
  inv01 U673 ( .Y(n1690), .A(n1841) );
  nor02 U674 ( .Y(n1842), .A0(n2236), .A1(n2380) );
  inv01 U675 ( .Y(n1843), .A(n2500) );
  nor02 U676 ( .Y(n1841), .A0(n1842), .A1(n1843) );
  inv01 U677 ( .Y(n1689), .A(n1844) );
  nor02 U678 ( .Y(n1845), .A0(n2235), .A1(n2380) );
  inv01 U679 ( .Y(n1846), .A(n2502) );
  nor02 U680 ( .Y(n1844), .A0(n1845), .A1(n1846) );
  inv01 U681 ( .Y(n1693), .A(n1847) );
  nor02 U682 ( .Y(n1848), .A0(n1905), .A1(n2380) );
  inv01 U683 ( .Y(n1849), .A(n2493) );
  nor02 U684 ( .Y(n1847), .A0(n1848), .A1(n1849) );
  inv01 U685 ( .Y(n1694), .A(n1850) );
  nor02 U686 ( .Y(n1851), .A0(n1902), .A1(n2380) );
  inv01 U687 ( .Y(n1852), .A(n2491) );
  nor02 U688 ( .Y(n1850), .A0(n1851), .A1(n1852) );
  inv01 U689 ( .Y(n1700), .A(n1853) );
  nor02 U690 ( .Y(n1854), .A0(n1901), .A1(n2379) );
  inv01 U691 ( .Y(n1855), .A(n2482) );
  nor02 U692 ( .Y(n1853), .A0(n1854), .A1(n1855) );
  inv01 U693 ( .Y(n1692), .A(n1856) );
  nor02 U694 ( .Y(n1857), .A0(n1901), .A1(n2380) );
  inv01 U695 ( .Y(n1858), .A(n2495) );
  nor02 U696 ( .Y(n1856), .A0(n1857), .A1(n1858) );
  inv01 U697 ( .Y(n1701), .A(n1859) );
  nor02 U698 ( .Y(n1860), .A0(n1905), .A1(n2379) );
  inv01 U699 ( .Y(n1861), .A(n2481) );
  nor02 U700 ( .Y(n1859), .A0(n1860), .A1(n1861) );
  inv01 U701 ( .Y(n1702), .A(n1862) );
  nor02 U702 ( .Y(n1863), .A0(n1902), .A1(n2379) );
  inv01 U703 ( .Y(n1864), .A(n2480) );
  nor02 U704 ( .Y(n1862), .A0(n1863), .A1(n1864) );
  inv01 U705 ( .Y(n1691), .A(n1865) );
  nor02 U706 ( .Y(n1866), .A0(n1900), .A1(n2380) );
  inv01 U707 ( .Y(n1867), .A(n2497) );
  nor02 U708 ( .Y(n1865), .A0(n1866), .A1(n1867) );
  inv01 U709 ( .Y(n1699), .A(n1868) );
  nor02 U710 ( .Y(n1869), .A0(n2469), .A1(n2379) );
  inv01 U711 ( .Y(n1870), .A(n2483) );
  nor02 U712 ( .Y(n1868), .A0(n1869), .A1(n1870) );
  inv01 U713 ( .Y(n1703), .A(n1871) );
  nor02 U714 ( .Y(n1872), .A0(n2284), .A1(n2379) );
  inv01 U715 ( .Y(n1873), .A(n2479) );
  nor02 U716 ( .Y(n1871), .A0(n1872), .A1(n1873) );
  inv01 U717 ( .Y(n1704), .A(n1874) );
  nor02 U718 ( .Y(n1875), .A0(n2285), .A1(n2379) );
  inv01 U719 ( .Y(n1876), .A(n2478) );
  nor02 U720 ( .Y(n1874), .A0(n1875), .A1(n1876) );
  inv01 U721 ( .Y(n1695), .A(n1877) );
  nor02 U722 ( .Y(n1878), .A0(n2284), .A1(n2380) );
  inv01 U723 ( .Y(n1879), .A(n2489) );
  nor02 U724 ( .Y(n1877), .A0(n1878), .A1(n1879) );
  inv01 U725 ( .Y(n1711), .A(n1880) );
  nor02 U726 ( .Y(n1881), .A0(n2381), .A1(n2284) );
  inv01 U727 ( .Y(n1882), .A(n2462) );
  nor02 U728 ( .Y(n1880), .A0(n1881), .A1(n1882) );
  inv01 U729 ( .Y(n1696), .A(n1883) );
  nor02 U730 ( .Y(n1884), .A0(n2285), .A1(n2380) );
  inv01 U731 ( .Y(n1885), .A(n2488) );
  nor02 U732 ( .Y(n1883), .A0(n1884), .A1(n1885) );
  inv01 U733 ( .Y(n1688), .A(n1886) );
  nor02 U734 ( .Y(n1887), .A0(n2280), .A1(n2285) );
  inv01 U735 ( .Y(n1888), .A(n2507) );
  nor02 U736 ( .Y(n1886), .A0(n1887), .A1(n1888) );
  nand02 U737 ( .Y(n1686), .A0(n1889), .A1(n1890) );
  inv01 U738 ( .Y(n1891), .A(n2550) );
  inv01 U739 ( .Y(n1892), .A(n2513) );
  inv01 U740 ( .Y(n1893), .A(n2385) );
  inv01 U741 ( .Y(n1894), .A(n2512) );
  nand02 U742 ( .Y(n1889), .A0(n1891), .A1(n1892) );
  nand02 U743 ( .Y(n1890), .A0(n1893), .A1(n1894) );
  inv01 U744 ( .Y(n1713), .A(n1895) );
  nor02 U745 ( .Y(n1896), .A0(n2386), .A1(n2541) );
  inv01 U746 ( .Y(n1897), .A(n1770) );
  nor02 U747 ( .Y(n1895), .A0(n1896), .A1(n1897) );
  or03 U748 ( .Y(n1898), .A0(n2280), .A1(s_count[0]), .A2(n2494) );
  inv01 U749 ( .Y(n1899), .A(n1898) );
  nand02 U750 ( .Y(n1900), .A0(n2238), .A1(n2248) );
  nand02 U751 ( .Y(n1901), .A0(n2237), .A1(n2245) );
  inv02 U752 ( .Y(n2245), .A(n2243) );
  buf02 U753 ( .Y(n1902), .A(n2463) );
  or03 U754 ( .Y(n1903), .A0(n2381), .A1(s_count[1]), .A2(s_count[0]) );
  inv01 U755 ( .Y(n1904), .A(n1903) );
  buf02 U756 ( .Y(n1905), .A(n2465) );
  or03 U757 ( .Y(n1906), .A0(s_dvdnd_i_42_), .A1(s_dvdnd_i_44_), .A2(
        s_dvdnd_i_43_) );
  inv01 U758 ( .Y(n1907), .A(n1906) );
  or03 U759 ( .Y(n1908), .A0(s_dvdnd_i_31_), .A1(s_dvdnd_i_33_), .A2(
        s_dvdnd_i_32_) );
  inv01 U760 ( .Y(n1909), .A(n1908) );
  ao21 U761 ( .Y(n1910), .A0(n2280), .A1(n2282), .B0(n2490) );
  inv01 U762 ( .Y(n1911), .A(n1910) );
  inv01 U763 ( .Y(n1765), .A(n1912) );
  nor02 U764 ( .Y(n1913), .A0(n2387), .A1(n2398) );
  nor02 U765 ( .Y(n1914), .A0(n2296), .A1(n2383) );
  nor02 U766 ( .Y(n1915), .A0(n2382), .A1(n2395) );
  nor02 U767 ( .Y(n1912), .A0(n1915), .A1(n1916) );
  nor02 U768 ( .Y(n1917), .A0(n1913), .A1(n1914) );
  inv01 U769 ( .Y(n1916), .A(n1917) );
  inv01 U770 ( .Y(n1762), .A(n1918) );
  nor02 U771 ( .Y(n1919), .A0(n2387), .A1(n2404) );
  nor02 U772 ( .Y(n1920), .A0(n2309), .A1(n2383) );
  nor02 U773 ( .Y(n1921), .A0(n2382), .A1(n2403) );
  nor02 U774 ( .Y(n1918), .A0(n1921), .A1(n1922) );
  nor02 U775 ( .Y(n1923), .A0(n1919), .A1(n1920) );
  inv01 U776 ( .Y(n1922), .A(n1923) );
  inv01 U777 ( .Y(n1749), .A(n1924) );
  nor02 U778 ( .Y(n1925), .A0(n2387), .A1(n2430) );
  nor02 U779 ( .Y(n1926), .A0(n2346), .A1(n2383) );
  nor02 U780 ( .Y(n1927), .A0(n2382), .A1(n2429) );
  nor02 U781 ( .Y(n1924), .A0(n1927), .A1(n1928) );
  nor02 U782 ( .Y(n1929), .A0(n1925), .A1(n1926) );
  inv01 U783 ( .Y(n1928), .A(n1929) );
  inv01 U784 ( .Y(n1763), .A(n1930) );
  nor02 U785 ( .Y(n1931), .A0(n2387), .A1(n2402) );
  nor02 U786 ( .Y(n1932), .A0(n2316), .A1(n2383) );
  nor02 U787 ( .Y(n1933), .A0(n2382), .A1(n2401) );
  nor02 U788 ( .Y(n1930), .A0(n1933), .A1(n1934) );
  nor02 U789 ( .Y(n1935), .A0(n1931), .A1(n1932) );
  inv01 U790 ( .Y(n1934), .A(n1935) );
  inv01 U791 ( .Y(n1757), .A(n1936) );
  nor02 U792 ( .Y(n1937), .A0(n2387), .A1(n2414) );
  nor02 U793 ( .Y(n1938), .A0(n2314), .A1(n2383) );
  nor02 U794 ( .Y(n1939), .A0(n2382), .A1(n2413) );
  nor02 U795 ( .Y(n1936), .A0(n1939), .A1(n1940) );
  nor02 U796 ( .Y(n1941), .A0(n1937), .A1(n1938) );
  inv01 U797 ( .Y(n1940), .A(n1941) );
  inv01 U798 ( .Y(n1745), .A(n1942) );
  nor02 U799 ( .Y(n1943), .A0(n2387), .A1(n2438) );
  nor02 U800 ( .Y(n1944), .A0(n2326), .A1(n2383) );
  nor02 U801 ( .Y(n1945), .A0(n2382), .A1(n2437) );
  nor02 U802 ( .Y(n1942), .A0(n1945), .A1(n1946) );
  nor02 U803 ( .Y(n1947), .A0(n1943), .A1(n1944) );
  inv01 U804 ( .Y(n1946), .A(n1947) );
  inv01 U805 ( .Y(n1746), .A(n1948) );
  nor02 U806 ( .Y(n1949), .A0(n2387), .A1(n2436) );
  nor02 U807 ( .Y(n1950), .A0(n2336), .A1(n2383) );
  nor02 U808 ( .Y(n1951), .A0(n2382), .A1(n2435) );
  nor02 U809 ( .Y(n1948), .A0(n1951), .A1(n1952) );
  nor02 U810 ( .Y(n1953), .A0(n1949), .A1(n1950) );
  inv01 U811 ( .Y(n1952), .A(n1953) );
  inv01 U812 ( .Y(n1751), .A(n1954) );
  nor02 U813 ( .Y(n1955), .A0(n2387), .A1(n2426) );
  nor02 U814 ( .Y(n1956), .A0(n2354), .A1(n2383) );
  nor02 U815 ( .Y(n1957), .A0(n2382), .A1(n2425) );
  nor02 U816 ( .Y(n1954), .A0(n1957), .A1(n1958) );
  nor02 U817 ( .Y(n1959), .A0(n1955), .A1(n1956) );
  inv01 U818 ( .Y(n1958), .A(n1959) );
  inv01 U819 ( .Y(n1750), .A(n1960) );
  nor02 U820 ( .Y(n1961), .A0(n2387), .A1(n2428) );
  nor02 U821 ( .Y(n1962), .A0(n2306), .A1(n2383) );
  nor02 U822 ( .Y(n1963), .A0(n2382), .A1(n2427) );
  nor02 U823 ( .Y(n1960), .A0(n1963), .A1(n1964) );
  nor02 U824 ( .Y(n1965), .A0(n1961), .A1(n1962) );
  inv01 U825 ( .Y(n1964), .A(n1965) );
  inv01 U826 ( .Y(n1761), .A(n1966) );
  nor02 U827 ( .Y(n1967), .A0(n2387), .A1(n2406) );
  nor02 U828 ( .Y(n1968), .A0(n2356), .A1(n2383) );
  nor02 U829 ( .Y(n1969), .A0(n2382), .A1(n2405) );
  nor02 U830 ( .Y(n1966), .A0(n1969), .A1(n1970) );
  nor02 U831 ( .Y(n1971), .A0(n1967), .A1(n1968) );
  inv01 U832 ( .Y(n1970), .A(n1971) );
  inv01 U833 ( .Y(n1756), .A(n1972) );
  nor02 U834 ( .Y(n1973), .A0(n2387), .A1(n2416) );
  nor02 U835 ( .Y(n1974), .A0(n2338), .A1(n2383) );
  nor02 U836 ( .Y(n1975), .A0(n2382), .A1(n2415) );
  nor02 U837 ( .Y(n1972), .A0(n1975), .A1(n1976) );
  nor02 U838 ( .Y(n1977), .A0(n1973), .A1(n1974) );
  inv01 U839 ( .Y(n1976), .A(n1977) );
  inv01 U840 ( .Y(n1747), .A(n1978) );
  nor02 U841 ( .Y(n1979), .A0(n2387), .A1(n2434) );
  nor02 U842 ( .Y(n1980), .A0(n2321), .A1(n2383) );
  nor02 U843 ( .Y(n1981), .A0(n2382), .A1(n2433) );
  nor02 U844 ( .Y(n1978), .A0(n1981), .A1(n1982) );
  nor02 U845 ( .Y(n1983), .A0(n1979), .A1(n1980) );
  inv01 U846 ( .Y(n1982), .A(n1983) );
  inv01 U847 ( .Y(n1759), .A(n1984) );
  nor02 U848 ( .Y(n1985), .A0(n2387), .A1(n2410) );
  nor02 U849 ( .Y(n1986), .A0(n2328), .A1(n2383) );
  nor02 U850 ( .Y(n1987), .A0(n2382), .A1(n2409) );
  nor02 U851 ( .Y(n1984), .A0(n1987), .A1(n1988) );
  nor02 U852 ( .Y(n1989), .A0(n1985), .A1(n1986) );
  inv01 U853 ( .Y(n1988), .A(n1989) );
  inv01 U854 ( .Y(n1758), .A(n1990) );
  nor02 U855 ( .Y(n1991), .A0(n2387), .A1(n2412) );
  nor02 U856 ( .Y(n1992), .A0(n2348), .A1(n2383) );
  nor02 U857 ( .Y(n1993), .A0(n2382), .A1(n2411) );
  nor02 U858 ( .Y(n1990), .A0(n1993), .A1(n1994) );
  nor02 U859 ( .Y(n1995), .A0(n1991), .A1(n1992) );
  inv01 U860 ( .Y(n1994), .A(n1995) );
  inv01 U861 ( .Y(n1760), .A(n1996) );
  nor02 U862 ( .Y(n1997), .A0(n2387), .A1(n2408) );
  nor02 U863 ( .Y(n1998), .A0(n2358), .A1(n2383) );
  nor02 U864 ( .Y(n1999), .A0(n2382), .A1(n2407) );
  nor02 U865 ( .Y(n1996), .A0(n1999), .A1(n2000) );
  nor02 U866 ( .Y(n2001), .A0(n1997), .A1(n1998) );
  inv01 U867 ( .Y(n2000), .A(n2001) );
  inv01 U868 ( .Y(n1748), .A(n2002) );
  nor02 U869 ( .Y(n2003), .A0(n2387), .A1(n2432) );
  nor02 U870 ( .Y(n2004), .A0(n2341), .A1(n2383) );
  nor02 U871 ( .Y(n2005), .A0(n2382), .A1(n2431) );
  nor02 U872 ( .Y(n2002), .A0(n2005), .A1(n2006) );
  nor02 U873 ( .Y(n2007), .A0(n2003), .A1(n2004) );
  inv01 U874 ( .Y(n2006), .A(n2007) );
  inv01 U875 ( .Y(n1755), .A(n2008) );
  nor02 U876 ( .Y(n2009), .A0(n2387), .A1(n2418) );
  nor02 U877 ( .Y(n2010), .A0(n2361), .A1(n2383) );
  nor02 U878 ( .Y(n2011), .A0(n2382), .A1(n2417) );
  nor02 U879 ( .Y(n2008), .A0(n2011), .A1(n2012) );
  nor02 U880 ( .Y(n2013), .A0(n2009), .A1(n2010) );
  inv01 U881 ( .Y(n2012), .A(n2013) );
  inv01 U882 ( .Y(n1754), .A(n2014) );
  nor02 U883 ( .Y(n2015), .A0(n2387), .A1(n2420) );
  nor02 U884 ( .Y(n2016), .A0(n2318), .A1(n2383) );
  nor02 U885 ( .Y(n2017), .A0(n2382), .A1(n2419) );
  nor02 U886 ( .Y(n2014), .A0(n2017), .A1(n2018) );
  nor02 U887 ( .Y(n2019), .A0(n2015), .A1(n2016) );
  inv01 U888 ( .Y(n2018), .A(n2019) );
  inv01 U889 ( .Y(n1753), .A(n2020) );
  nor02 U890 ( .Y(n2021), .A0(n2387), .A1(n2422) );
  nor02 U891 ( .Y(n2022), .A0(n2351), .A1(n2383) );
  nor02 U892 ( .Y(n2023), .A0(n2382), .A1(n2421) );
  nor02 U893 ( .Y(n2020), .A0(n2023), .A1(n2024) );
  nor02 U894 ( .Y(n2025), .A0(n2021), .A1(n2022) );
  inv01 U895 ( .Y(n2024), .A(n2025) );
  inv01 U896 ( .Y(n1752), .A(n2026) );
  nor02 U897 ( .Y(n2027), .A0(n2387), .A1(n2424) );
  nor02 U898 ( .Y(n2028), .A0(n2311), .A1(n2383) );
  nor02 U899 ( .Y(n2029), .A0(n2382), .A1(n2423) );
  nor02 U900 ( .Y(n2026), .A0(n2029), .A1(n2030) );
  nor02 U901 ( .Y(n2031), .A0(n2027), .A1(n2028) );
  inv01 U902 ( .Y(n2030), .A(n2031) );
  inv01 U903 ( .Y(n1764), .A(n2032) );
  nor02 U904 ( .Y(n2033), .A0(n2387), .A1(n2400) );
  nor02 U905 ( .Y(n2034), .A0(n2331), .A1(n2383) );
  nor02 U906 ( .Y(n2035), .A0(n2382), .A1(n2399) );
  nor02 U907 ( .Y(n2032), .A0(n2035), .A1(n2036) );
  nor02 U908 ( .Y(n2037), .A0(n2033), .A1(n2034) );
  inv01 U909 ( .Y(n2036), .A(n2037) );
  inv01 U910 ( .Y(n1744), .A(n2038) );
  nor02 U911 ( .Y(n2039), .A0(n2387), .A1(n2440) );
  nor02 U912 ( .Y(n2040), .A0(n2334), .A1(n2383) );
  nor02 U913 ( .Y(n2041), .A0(n2382), .A1(n2439) );
  nor02 U914 ( .Y(n2038), .A0(n2041), .A1(n2042) );
  nor02 U915 ( .Y(n2043), .A0(n2039), .A1(n2040) );
  inv01 U916 ( .Y(n2042), .A(n2043) );
  inv01 U917 ( .Y(n1742), .A(n2044) );
  nor02 U918 ( .Y(n2045), .A0(n2387), .A1(n2444) );
  nor02 U919 ( .Y(n2046), .A0(n2344), .A1(n2383) );
  nor02 U920 ( .Y(n2047), .A0(n2382), .A1(n2443) );
  nor02 U921 ( .Y(n2044), .A0(n2047), .A1(n2048) );
  nor02 U922 ( .Y(n2049), .A0(n2045), .A1(n2046) );
  inv01 U923 ( .Y(n2048), .A(n2049) );
  inv01 U924 ( .Y(n1743), .A(n2050) );
  nor02 U925 ( .Y(n2051), .A0(n2387), .A1(n2442) );
  nor02 U926 ( .Y(n2052), .A0(n2324), .A1(n2383) );
  nor02 U927 ( .Y(n2053), .A0(n2382), .A1(n2441) );
  nor02 U928 ( .Y(n2050), .A0(n2053), .A1(n2054) );
  nor02 U929 ( .Y(n2055), .A0(n2051), .A1(n2052) );
  inv01 U930 ( .Y(n2054), .A(n2055) );
  inv01 U931 ( .Y(n1741), .A(n2056) );
  nor02 U932 ( .Y(n2057), .A0(n2387), .A1(n2447) );
  nor02 U933 ( .Y(n2058), .A0(n2383), .A1(n2291) );
  nor02 U934 ( .Y(n2059), .A0(n2382), .A1(n2445) );
  nor02 U935 ( .Y(n2056), .A0(n2059), .A1(n2060) );
  nor02 U936 ( .Y(n2061), .A0(n2057), .A1(n2058) );
  inv01 U937 ( .Y(n2060), .A(n2061) );
  inv01 U938 ( .Y(n1740), .A(n2062) );
  nor02 U939 ( .Y(n2063), .A0(n2387), .A1(n2450) );
  nor02 U940 ( .Y(n2064), .A0(n2383), .A1(n2290) );
  nor02 U941 ( .Y(n2065), .A0(n2382), .A1(n2448) );
  nor02 U942 ( .Y(n2062), .A0(n2065), .A1(n2066) );
  nor02 U943 ( .Y(n2067), .A0(n2063), .A1(n2064) );
  inv01 U944 ( .Y(n2066), .A(n2067) );
  inv02 U945 ( .Y(L546_20_), .A(n2326) );
  inv02 U946 ( .Y(L546_19_), .A(n2336) );
  inv02 U947 ( .Y(L546_16_), .A(n2346) );
  inv02 U948 ( .Y(L546_15_), .A(n2306) );
  inv02 U949 ( .Y(L546_14_), .A(n2354) );
  inv02 U950 ( .Y(L546_8_), .A(n2314) );
  inv02 U951 ( .Y(L546_4_), .A(n2356) );
  inv02 U952 ( .Y(L546_2_), .A(n2316) );
  inv01 U953 ( .Y(n1730), .A(n2068) );
  nor02 U954 ( .Y(n2069), .A0(n2371), .A1(n1680) );
  nor02 U955 ( .Y(n2070), .A0(n2339), .A1(n2388) );
  nor02 U956 ( .Y(n2071), .A0(n2415), .A1(n2385) );
  nor02 U957 ( .Y(n2068), .A0(n2071), .A1(n2072) );
  nor02 U958 ( .Y(n2073), .A0(n2069), .A1(n2070) );
  inv01 U959 ( .Y(n2072), .A(n2073) );
  inv01 U960 ( .Y(n1718), .A(n2074) );
  nor02 U961 ( .Y(n2075), .A0(n2371), .A1(n1668) );
  nor02 U962 ( .Y(n2076), .A0(n2334), .A1(n2388) );
  nor02 U963 ( .Y(n2077), .A0(n2439), .A1(n2385) );
  nor02 U964 ( .Y(n2074), .A0(n2077), .A1(n2078) );
  nor02 U965 ( .Y(n2079), .A0(n2075), .A1(n2076) );
  inv01 U966 ( .Y(n2078), .A(n2079) );
  inv01 U967 ( .Y(n1723), .A(n2080) );
  nor02 U968 ( .Y(n2081), .A0(n2386), .A1(n1662) );
  nor02 U969 ( .Y(n2082), .A0(n2346), .A1(n2388) );
  nor02 U970 ( .Y(n2083), .A0(n2429), .A1(n2385) );
  nor02 U971 ( .Y(n2080), .A0(n2083), .A1(n2084) );
  nor02 U972 ( .Y(n2085), .A0(n2081), .A1(n2082) );
  inv01 U973 ( .Y(n2084), .A(n2085) );
  inv01 U974 ( .Y(n1716), .A(n2086) );
  nor02 U975 ( .Y(n2087), .A0(n2386), .A1(n1670) );
  nor02 U976 ( .Y(n2088), .A0(n2344), .A1(n2388) );
  nor02 U977 ( .Y(n2089), .A0(n2443), .A1(n2385) );
  nor02 U978 ( .Y(n2086), .A0(n2089), .A1(n2090) );
  nor02 U979 ( .Y(n2091), .A0(n2087), .A1(n2088) );
  inv01 U980 ( .Y(n2090), .A(n2091) );
  inv01 U981 ( .Y(n1735), .A(n2092) );
  nor02 U982 ( .Y(n2093), .A0(n2371), .A1(n1675) );
  nor02 U983 ( .Y(n2094), .A0(n2356), .A1(n2388) );
  nor02 U984 ( .Y(n2095), .A0(n2405), .A1(n2385) );
  nor02 U985 ( .Y(n2092), .A0(n2095), .A1(n2096) );
  nor02 U986 ( .Y(n2097), .A0(n2093), .A1(n2094) );
  inv01 U987 ( .Y(n2096), .A(n2097) );
  inv01 U988 ( .Y(n1729), .A(n2098) );
  nor02 U989 ( .Y(n2099), .A0(n2386), .A1(n1656) );
  nor02 U990 ( .Y(n2100), .A0(n2362), .A1(n2388) );
  nor02 U991 ( .Y(n2101), .A0(n2417), .A1(n2385) );
  nor02 U992 ( .Y(n2098), .A0(n2101), .A1(n2102) );
  nor02 U993 ( .Y(n2103), .A0(n2099), .A1(n2100) );
  inv01 U994 ( .Y(n2102), .A(n2103) );
  inv01 U995 ( .Y(n1734), .A(n2104) );
  nor02 U996 ( .Y(n2105), .A0(n2386), .A1(n1676) );
  nor02 U997 ( .Y(n2106), .A0(n2359), .A1(n2388) );
  nor02 U998 ( .Y(n2107), .A0(n2407), .A1(n2385) );
  nor02 U999 ( .Y(n2104), .A0(n2107), .A1(n2108) );
  nor02 U1000 ( .Y(n2109), .A0(n2105), .A1(n2106) );
  inv01 U1001 ( .Y(n2108), .A(n2109) );
  inv01 U1002 ( .Y(n1719), .A(n2110) );
  nor02 U1003 ( .Y(n2111), .A0(n2386), .A1(n1667) );
  nor02 U1004 ( .Y(n2112), .A0(n2326), .A1(n2388) );
  nor02 U1005 ( .Y(n2113), .A0(n2437), .A1(n2385) );
  nor02 U1006 ( .Y(n2110), .A0(n2113), .A1(n2114) );
  nor02 U1007 ( .Y(n2115), .A0(n2111), .A1(n2112) );
  inv01 U1008 ( .Y(n2114), .A(n2115) );
  inv01 U1009 ( .Y(n1731), .A(n2116) );
  nor02 U1010 ( .Y(n2117), .A0(n2386), .A1(n1679) );
  nor02 U1011 ( .Y(n2118), .A0(n2314), .A1(n2388) );
  nor02 U1012 ( .Y(n2119), .A0(n2413), .A1(n2385) );
  nor02 U1013 ( .Y(n2116), .A0(n2119), .A1(n2120) );
  nor02 U1014 ( .Y(n2121), .A0(n2117), .A1(n2118) );
  inv01 U1015 ( .Y(n2120), .A(n2121) );
  inv01 U1016 ( .Y(n1733), .A(n2122) );
  nor02 U1017 ( .Y(n2123), .A0(n2386), .A1(n1677) );
  nor02 U1018 ( .Y(n2124), .A0(n2329), .A1(n2388) );
  nor02 U1019 ( .Y(n2125), .A0(n2409), .A1(n2385) );
  nor02 U1020 ( .Y(n2122), .A0(n2125), .A1(n2126) );
  nor02 U1021 ( .Y(n2127), .A0(n2123), .A1(n2124) );
  inv01 U1022 ( .Y(n2126), .A(n2127) );
  inv01 U1023 ( .Y(n1721), .A(n2128) );
  nor02 U1024 ( .Y(n2129), .A0(n2386), .A1(n1664) );
  nor02 U1025 ( .Y(n2130), .A0(n2322), .A1(n2388) );
  nor02 U1026 ( .Y(n2131), .A0(n2433), .A1(n2385) );
  nor02 U1027 ( .Y(n2128), .A0(n2131), .A1(n2132) );
  nor02 U1028 ( .Y(n2133), .A0(n2129), .A1(n2130) );
  inv01 U1029 ( .Y(n2132), .A(n2133) );
  inv01 U1030 ( .Y(n1724), .A(n2134) );
  nor02 U1031 ( .Y(n2135), .A0(n2386), .A1(n1661) );
  nor02 U1032 ( .Y(n2136), .A0(n2306), .A1(n2388) );
  nor02 U1033 ( .Y(n2137), .A0(n2427), .A1(n2385) );
  nor02 U1034 ( .Y(n2134), .A0(n2137), .A1(n2138) );
  nor02 U1035 ( .Y(n2139), .A0(n2135), .A1(n2136) );
  inv01 U1036 ( .Y(n2138), .A(n2139) );
  inv01 U1037 ( .Y(n1736), .A(n2140) );
  nor02 U1038 ( .Y(n2141), .A0(n2386), .A1(n1674) );
  nor02 U1039 ( .Y(n2142), .A0(n2308), .A1(n2388) );
  nor02 U1040 ( .Y(n2143), .A0(n2403), .A1(n2385) );
  nor02 U1041 ( .Y(n2140), .A0(n2143), .A1(n2144) );
  nor02 U1042 ( .Y(n2145), .A0(n2141), .A1(n2142) );
  inv01 U1043 ( .Y(n2144), .A(n2145) );
  inv01 U1044 ( .Y(n1720), .A(n2146) );
  nor02 U1045 ( .Y(n2147), .A0(n2386), .A1(n1665) );
  nor02 U1046 ( .Y(n2148), .A0(n2336), .A1(n2388) );
  nor02 U1047 ( .Y(n2149), .A0(n2435), .A1(n2385) );
  nor02 U1048 ( .Y(n2146), .A0(n2149), .A1(n2150) );
  nor02 U1049 ( .Y(n2151), .A0(n2147), .A1(n2148) );
  inv01 U1050 ( .Y(n2150), .A(n2151) );
  inv01 U1051 ( .Y(n1717), .A(n2152) );
  nor02 U1052 ( .Y(n2153), .A0(n2386), .A1(n1669) );
  nor02 U1053 ( .Y(n2154), .A0(n2324), .A1(n2388) );
  nor02 U1054 ( .Y(n2155), .A0(n2441), .A1(n2385) );
  nor02 U1055 ( .Y(n2152), .A0(n2155), .A1(n2156) );
  nor02 U1056 ( .Y(n2157), .A0(n2153), .A1(n2154) );
  inv01 U1057 ( .Y(n2156), .A(n2157) );
  inv01 U1058 ( .Y(n1722), .A(n2158) );
  nor02 U1059 ( .Y(n2159), .A0(n2386), .A1(n1663) );
  nor02 U1060 ( .Y(n2160), .A0(n2342), .A1(n2388) );
  nor02 U1061 ( .Y(n2161), .A0(n2431), .A1(n2385) );
  nor02 U1062 ( .Y(n2158), .A0(n2161), .A1(n2162) );
  nor02 U1063 ( .Y(n2163), .A0(n2159), .A1(n2160) );
  inv01 U1064 ( .Y(n2162), .A(n2163) );
  inv01 U1065 ( .Y(n1727), .A(n2164) );
  nor02 U1066 ( .Y(n2165), .A0(n2386), .A1(n1658) );
  nor02 U1067 ( .Y(n2166), .A0(n2352), .A1(n2388) );
  nor02 U1068 ( .Y(n2167), .A0(n2421), .A1(n2385) );
  nor02 U1069 ( .Y(n2164), .A0(n2167), .A1(n2168) );
  nor02 U1070 ( .Y(n2169), .A0(n2165), .A1(n2166) );
  inv01 U1071 ( .Y(n2168), .A(n2169) );
  inv01 U1072 ( .Y(n1714), .A(n2170) );
  nor02 U1073 ( .Y(n2171), .A0(n2386), .A1(n1672) );
  nor02 U1074 ( .Y(n2172), .A0(n2290), .A1(n2388) );
  nor02 U1075 ( .Y(n2173), .A0(n2448), .A1(n2385) );
  nor02 U1076 ( .Y(n2170), .A0(n2173), .A1(n2174) );
  nor02 U1077 ( .Y(n2175), .A0(n2171), .A1(n2172) );
  inv01 U1078 ( .Y(n2174), .A(n2175) );
  inv01 U1079 ( .Y(n1725), .A(n2176) );
  nor02 U1080 ( .Y(n2177), .A0(n2386), .A1(n1660) );
  nor02 U1081 ( .Y(n2178), .A0(n2354), .A1(n2388) );
  nor02 U1082 ( .Y(n2179), .A0(n2425), .A1(n2385) );
  nor02 U1083 ( .Y(n2176), .A0(n2179), .A1(n2180) );
  nor02 U1084 ( .Y(n2181), .A0(n2177), .A1(n2178) );
  inv01 U1085 ( .Y(n2180), .A(n2181) );
  inv01 U1086 ( .Y(n1737), .A(n2182) );
  nor02 U1087 ( .Y(n2183), .A0(n2386), .A1(n1673) );
  nor02 U1088 ( .Y(n2184), .A0(n2316), .A1(n2388) );
  nor02 U1089 ( .Y(n2185), .A0(n2401), .A1(n2385) );
  nor02 U1090 ( .Y(n2182), .A0(n2185), .A1(n2186) );
  nor02 U1091 ( .Y(n2187), .A0(n2183), .A1(n2184) );
  inv01 U1092 ( .Y(n2186), .A(n2187) );
  inv01 U1093 ( .Y(n1732), .A(n2188) );
  nor02 U1094 ( .Y(n2189), .A0(n2386), .A1(n1678) );
  nor02 U1095 ( .Y(n2190), .A0(n2349), .A1(n2388) );
  nor02 U1096 ( .Y(n2191), .A0(n2411), .A1(n2385) );
  nor02 U1097 ( .Y(n2188), .A0(n2191), .A1(n2192) );
  nor02 U1098 ( .Y(n2193), .A0(n2189), .A1(n2190) );
  inv01 U1099 ( .Y(n2192), .A(n2193) );
  inv01 U1100 ( .Y(n1715), .A(n2194) );
  nor02 U1101 ( .Y(n2195), .A0(n2386), .A1(n1671) );
  nor02 U1102 ( .Y(n2196), .A0(n2291), .A1(n2388) );
  nor02 U1103 ( .Y(n2197), .A0(n2445), .A1(n2385) );
  nor02 U1104 ( .Y(n2194), .A0(n2197), .A1(n2198) );
  nor02 U1105 ( .Y(n2199), .A0(n2195), .A1(n2196) );
  inv01 U1106 ( .Y(n2198), .A(n2199) );
  inv01 U1107 ( .Y(n1726), .A(n2200) );
  nor02 U1108 ( .Y(n2201), .A0(n2386), .A1(n1659) );
  nor02 U1109 ( .Y(n2202), .A0(n2312), .A1(n2388) );
  nor02 U1110 ( .Y(n2203), .A0(n2423), .A1(n2385) );
  nor02 U1111 ( .Y(n2200), .A0(n2203), .A1(n2204) );
  nor02 U1112 ( .Y(n2205), .A0(n2201), .A1(n2202) );
  inv01 U1113 ( .Y(n2204), .A(n2205) );
  inv01 U1114 ( .Y(n1728), .A(n2206) );
  nor02 U1115 ( .Y(n2207), .A0(n2386), .A1(n1657) );
  nor02 U1116 ( .Y(n2208), .A0(n2319), .A1(n2388) );
  nor02 U1117 ( .Y(n2209), .A0(n2419), .A1(n2385) );
  nor02 U1118 ( .Y(n2206), .A0(n2209), .A1(n2210) );
  nor02 U1119 ( .Y(n2211), .A0(n2207), .A1(n2208) );
  inv01 U1120 ( .Y(n2210), .A(n2211) );
  inv01 U1121 ( .Y(n1738), .A(n2212) );
  nor02 U1122 ( .Y(n2213), .A0(n2386), .A1(n1666) );
  nor02 U1123 ( .Y(n2214), .A0(n2332), .A1(n2388) );
  nor02 U1124 ( .Y(n2215), .A0(n2399), .A1(n2385) );
  nor02 U1125 ( .Y(n2212), .A0(n2215), .A1(n2216) );
  nor02 U1126 ( .Y(n2217), .A0(n2213), .A1(n2214) );
  inv01 U1127 ( .Y(n2216), .A(n2217) );
  inv01 U1128 ( .Y(n1739), .A(n2218) );
  nor02 U1129 ( .Y(n2219), .A0(n2386), .A1(n1655) );
  nor02 U1130 ( .Y(n2220), .A0(n2295), .A1(n2388) );
  nor02 U1131 ( .Y(n2221), .A0(n2395), .A1(n2385) );
  nor02 U1132 ( .Y(n2218), .A0(n2221), .A1(n2222) );
  nor02 U1133 ( .Y(n2223), .A0(n2219), .A1(n2220) );
  inv01 U1134 ( .Y(n2222), .A(n2223) );
  or04 U1135 ( .Y(n2224), .A0(s_dvdnd_i_5_), .A1(s_dvdnd_i_4_), .A2(
        s_dvdnd_i_49_), .A3(s_dvdnd_i_48_) );
  inv01 U1136 ( .Y(n2225), .A(n2224) );
  or04 U1137 ( .Y(n2226), .A0(s_dvdnd_i_46_), .A1(s_dvdnd_i_47_), .A2(
        s_dvdnd_i_45_), .A3(n2535) );
  inv01 U1138 ( .Y(n2227), .A(n2226) );
  or04 U1139 ( .Y(n2228), .A0(s_dvdnd_i_35_), .A1(s_dvdnd_i_36_), .A2(
        s_dvdnd_i_34_), .A3(n2532) );
  inv01 U1140 ( .Y(n2229), .A(n2228) );
  inv01 U1141 ( .Y(n2230), .A(n2503) );
  nor02 U1142 ( .Y(div_zero_o), .A0(n2231), .A1(n2232) );
  nor02 U1143 ( .Y(n2233), .A0(n2520), .A1(n2521) );
  inv01 U1144 ( .Y(n2231), .A(n2233) );
  nor02 U1145 ( .Y(n2234), .A0(n2522), .A1(n2523) );
  inv01 U1146 ( .Y(n2232), .A(n2234) );
  buf02 U1147 ( .Y(n2235), .A(n2475) );
  buf02 U1148 ( .Y(n2236), .A(n2471) );
  buf02 U1149 ( .Y(n2237), .A(n2496) );
  buf02 U1150 ( .Y(n2238), .A(n2496) );
  or02 U1151 ( .Y(n2239), .A0(n____return556), .A1(n2391) );
  inv01 U1152 ( .Y(n2240), .A(n2239) );
  or04 U1153 ( .Y(n2241), .A0(n2540), .A1(n2588), .A2(n2586), .A3(n2587) );
  inv01 U1154 ( .Y(n2242), .A(n2241) );
  nand02 U1155 ( .Y(n2243), .A0(n2240), .A1(n2369) );
  inv01 U1156 ( .Y(n2244), .A(n2243) );
  inv01 U1157 ( .Y(n2246), .A(n2243) );
  nand02 U1158 ( .Y(n2247), .A0(n2474), .A1(n2240) );
  inv02 U1159 ( .Y(n2248), .A(n2247) );
  or04 U1160 ( .Y(n2249), .A0(n2539), .A1(n2576), .A2(n2572), .A3(n2573) );
  inv01 U1161 ( .Y(n2250), .A(n2249) );
  or04 U1162 ( .Y(n2251), .A0(n2536), .A1(n2537), .A2(s_dvdnd_i_14_), .A3(
        n2538) );
  inv01 U1163 ( .Y(n2252), .A(n2251) );
  or04 U1164 ( .Y(n2253), .A0(s_dvdnd_i_28_), .A1(s_dvdnd_i_27_), .A2(
        s_dvdnd_i_26_), .A3(s_dvdnd_i_25_) );
  inv01 U1165 ( .Y(n2254), .A(n2253) );
  inv01 U1166 ( .Y(n1768), .A(n2255) );
  nor02 U1167 ( .Y(n2256), .A0(n2293), .A1(n2257) );
  nor02 U1168 ( .Y(n2258), .A0(n2391), .A1(n1654) );
  nor02 U1169 ( .Y(n2255), .A0(n2256), .A1(n2258) );
  nor02 U1170 ( .Y(n2259), .A0(n2389), .A1(n2390) );
  inv01 U1171 ( .Y(n2257), .A(n2259) );
  or04 U1172 ( .Y(n2260), .A0(s_dvsor_i_20_), .A1(s_dvsor_i_1_), .A2(
        s_dvsor_i_19_), .A3(s_dvsor_i_18_) );
  inv01 U1173 ( .Y(n2261), .A(n2260) );
  or04 U1174 ( .Y(n2262), .A0(s_dvsor_i_14_), .A1(s_dvsor_i_13_), .A2(
        s_dvsor_i_12_), .A3(s_dvsor_i_11_) );
  inv01 U1175 ( .Y(n2263), .A(n2262) );
  or04 U1176 ( .Y(n2264), .A0(s_dvsor_i_9_), .A1(s_dvsor_i_8_), .A2(
        s_dvsor_i_7_), .A3(s_dvsor_i_6_) );
  inv01 U1177 ( .Y(n2265), .A(n2264) );
  or04 U1178 ( .Y(n2266), .A0(s_dvsor_i_2_), .A1(s_dvsor_i_26_), .A2(
        s_dvsor_i_25_), .A3(s_dvsor_i_24_) );
  inv01 U1179 ( .Y(n2267), .A(n2266) );
  or03 U1180 ( .Y(n2268), .A0(n2391), .A1(s_state355), .A2(n2451) );
  inv01 U1181 ( .Y(n2269), .A(n2268) );
  inv01 U1182 ( .Y(n2270), .A(n2268) );
  inv01 U1183 ( .Y(n2525), .A(n2271) );
  inv01 U1184 ( .Y(n2272), .A(n2529) );
  inv01 U1185 ( .Y(n2273), .A(n2528) );
  inv01 U1186 ( .Y(n2274), .A(n2527) );
  inv01 U1187 ( .Y(n2275), .A(n2526) );
  nand02 U1188 ( .Y(n2271), .A0(n2276), .A1(n2277) );
  nand02 U1189 ( .Y(n2278), .A0(n2272), .A1(n2273) );
  inv01 U1190 ( .Y(n2276), .A(n2278) );
  nand02 U1191 ( .Y(n2279), .A0(n2274), .A1(n2275) );
  inv01 U1192 ( .Y(n2277), .A(n2279) );
  buf02 U1193 ( .Y(n2280), .A(n2506) );
  buf02 U1194 ( .Y(n2281), .A(n2473) );
  buf02 U1195 ( .Y(n2283), .A(n2473) );
  buf04 U1196 ( .Y(n2282), .A(n2473) );
  inv02 U1197 ( .Y(n2473), .A(s_state355) );
  buf02 U1198 ( .Y(n2284), .A(n2461) );
  buf02 U1199 ( .Y(n2285), .A(n2457) );
  inv02 U1200 ( .Y(n2287), .A(n2286) );
  ao21 U1201 ( .Y(n2288), .A0(n2518), .A1(s_state), .B0(s_state355) );
  inv02 U1202 ( .Y(n2289), .A(n2288) );
  buf02 U1203 ( .Y(n2290), .A(n2449) );
  buf02 U1204 ( .Y(n2291), .A(n2446) );
  inv02 U1205 ( .Y(L546_25_), .A(n2290) );
  inv02 U1206 ( .Y(L546_24_), .A(n2291) );
  nor02 U1207 ( .Y(n2292), .A0(n2381), .A1(n2511) );
  inv02 U1208 ( .Y(n2293), .A(n2292) );
  ao22 U1209 ( .Y(n2294), .A0(s_dvd[0]), .A1(n2512), .B0(s_dvdnd_i_26_), .B1(
        n2384) );
  inv01 U1210 ( .Y(n2295), .A(n2294) );
  inv02 U1211 ( .Y(n2296), .A(n2294) );
  inv02 U1212 ( .Y(L546_0_), .A(n2296) );
  inv02 U1213 ( .Y(n2499), .A(s_count[2]) );
  ao21 U1214 ( .Y(n2297), .A0(n2379), .A1(n2282), .B0(n2474) );
  inv02 U1215 ( .Y(n2298), .A(n2297) );
  ao21 U1216 ( .Y(n2299), .A0(n2380), .A1(n2281), .B0(n2370) );
  inv02 U1217 ( .Y(n2300), .A(n2299) );
  ao21 U1218 ( .Y(n2301), .A0(n2379), .A1(n2283), .B0(n2370) );
  inv02 U1219 ( .Y(n2302), .A(n2301) );
  ao21 U1220 ( .Y(n2303), .A0(n2380), .A1(n2281), .B0(n2474) );
  inv02 U1221 ( .Y(n2304), .A(n2303) );
  ao22 U1222 ( .Y(n2305), .A0(s_dvd[15]), .A1(n2512), .B0(s_dvdnd_i_41_), .B1(
        n2384) );
  inv02 U1223 ( .Y(n2306), .A(n2305) );
  ao22 U1224 ( .Y(n2307), .A0(s_dvd[3]), .A1(n2512), .B0(s_dvdnd_i_29_), .B1(
        n2384) );
  inv01 U1225 ( .Y(n2308), .A(n2307) );
  inv02 U1226 ( .Y(n2309), .A(n2307) );
  ao22 U1227 ( .Y(n2310), .A0(s_dvd[13]), .A1(n2512), .B0(s_dvdnd_i_39_), .B1(
        n2384) );
  inv01 U1228 ( .Y(n2311), .A(n2310) );
  inv02 U1229 ( .Y(n2312), .A(n2310) );
  inv02 U1230 ( .Y(L546_3_), .A(n2309) );
  inv02 U1231 ( .Y(L546_13_), .A(n2312) );
  ao22 U1232 ( .Y(n2313), .A0(s_dvd[8]), .A1(n2512), .B0(s_dvdnd_i_34_), .B1(
        n2384) );
  inv02 U1233 ( .Y(n2314), .A(n2313) );
  ao22 U1234 ( .Y(n2315), .A0(s_dvd[2]), .A1(n2512), .B0(s_dvdnd_i_28_), .B1(
        n2384) );
  inv02 U1235 ( .Y(n2316), .A(n2315) );
  ao22 U1236 ( .Y(n2317), .A0(s_dvd[11]), .A1(n2512), .B0(s_dvdnd_i_37_), .B1(
        n2384) );
  inv01 U1237 ( .Y(n2318), .A(n2317) );
  inv02 U1238 ( .Y(n2319), .A(n2317) );
  ao22 U1239 ( .Y(n2320), .A0(s_dvd[18]), .A1(n2512), .B0(s_dvdnd_i_44_), .B1(
        n2384) );
  inv01 U1240 ( .Y(n2321), .A(n2320) );
  inv02 U1241 ( .Y(n2322), .A(n2320) );
  inv02 U1242 ( .Y(L546_11_), .A(n2319) );
  inv02 U1243 ( .Y(L546_18_), .A(n2322) );
  ao22 U1244 ( .Y(n2323), .A0(s_dvd[22]), .A1(n2512), .B0(s_dvdnd_i_48_), .B1(
        n2384) );
  inv02 U1245 ( .Y(n2324), .A(n2323) );
  ao22 U1246 ( .Y(n2325), .A0(s_dvd[20]), .A1(n2512), .B0(s_dvdnd_i_46_), .B1(
        n2384) );
  inv02 U1247 ( .Y(n2326), .A(n2325) );
  ao22 U1248 ( .Y(n2327), .A0(s_dvd[6]), .A1(n2512), .B0(s_dvdnd_i_32_), .B1(
        n2384) );
  inv01 U1249 ( .Y(n2328), .A(n2327) );
  inv02 U1250 ( .Y(n2329), .A(n2327) );
  ao22 U1251 ( .Y(n2330), .A0(s_dvd[1]), .A1(n2512), .B0(s_dvdnd_i_27_), .B1(
        n2384) );
  inv01 U1252 ( .Y(n2331), .A(n2330) );
  inv02 U1253 ( .Y(n2332), .A(n2330) );
  inv02 U1254 ( .Y(L546_6_), .A(n2329) );
  inv02 U1255 ( .Y(L546_1_), .A(n2332) );
  inv04 U1256 ( .Y(L546_22_), .A(n2324) );
  ao22 U1257 ( .Y(n2333), .A0(s_dvd[21]), .A1(n2512), .B0(s_dvdnd_i_47_), .B1(
        n2384) );
  inv02 U1258 ( .Y(n2334), .A(n2333) );
  ao22 U1259 ( .Y(n2335), .A0(s_dvd[19]), .A1(n2512), .B0(s_dvdnd_i_45_), .B1(
        n2384) );
  inv02 U1260 ( .Y(n2336), .A(n2335) );
  ao22 U1261 ( .Y(n2337), .A0(s_dvd[9]), .A1(n2512), .B0(s_dvdnd_i_35_), .B1(
        n2384) );
  inv01 U1262 ( .Y(n2338), .A(n2337) );
  inv02 U1263 ( .Y(n2339), .A(n2337) );
  ao22 U1264 ( .Y(n2340), .A0(s_dvd[17]), .A1(n2512), .B0(s_dvdnd_i_43_), .B1(
        n2384) );
  inv01 U1265 ( .Y(n2341), .A(n2340) );
  inv02 U1266 ( .Y(n2342), .A(n2340) );
  inv02 U1267 ( .Y(L546_9_), .A(n2339) );
  inv02 U1268 ( .Y(L546_17_), .A(n2342) );
  inv04 U1269 ( .Y(L546_21_), .A(n2334) );
  ao22 U1270 ( .Y(n2343), .A0(s_dvd[23]), .A1(n2512), .B0(s_dvdnd_i_49_), .B1(
        n2384) );
  inv02 U1271 ( .Y(n2344), .A(n2343) );
  ao22 U1272 ( .Y(n2345), .A0(s_dvd[16]), .A1(n2512), .B0(s_dvdnd_i_42_), .B1(
        n2384) );
  inv02 U1273 ( .Y(n2346), .A(n2345) );
  ao22 U1274 ( .Y(n2347), .A0(s_dvd[7]), .A1(n2512), .B0(s_dvdnd_i_33_), .B1(
        n2384) );
  inv01 U1275 ( .Y(n2348), .A(n2347) );
  inv02 U1276 ( .Y(n2349), .A(n2347) );
  ao22 U1277 ( .Y(n2350), .A0(s_dvd[12]), .A1(n2512), .B0(s_dvdnd_i_38_), .B1(
        n2384) );
  inv01 U1278 ( .Y(n2351), .A(n2350) );
  inv02 U1279 ( .Y(n2352), .A(n2350) );
  inv02 U1280 ( .Y(L546_7_), .A(n2349) );
  inv02 U1281 ( .Y(L546_12_), .A(n2352) );
  inv04 U1282 ( .Y(L546_23_), .A(n2344) );
  ao22 U1283 ( .Y(n2353), .A0(s_dvd[14]), .A1(n2512), .B0(s_dvdnd_i_40_), .B1(
        n2384) );
  inv02 U1284 ( .Y(n2354), .A(n2353) );
  ao22 U1285 ( .Y(n2355), .A0(s_dvd[4]), .A1(n2512), .B0(s_dvdnd_i_30_), .B1(
        n2384) );
  inv02 U1286 ( .Y(n2356), .A(n2355) );
  ao22 U1287 ( .Y(n2357), .A0(s_dvd[5]), .A1(n2512), .B0(s_dvdnd_i_31_), .B1(
        n2384) );
  inv01 U1288 ( .Y(n2358), .A(n2357) );
  inv02 U1289 ( .Y(n2359), .A(n2357) );
  ao22 U1290 ( .Y(n2360), .A0(s_dvd[10]), .A1(n2512), .B0(s_dvdnd_i_36_), .B1(
        n2384) );
  inv01 U1291 ( .Y(n2361), .A(n2360) );
  inv02 U1292 ( .Y(n2362), .A(n2360) );
  inv02 U1293 ( .Y(L546_5_), .A(n2359) );
  inv02 U1294 ( .Y(L546_10_), .A(n2362) );
  ao21 U1295 ( .Y(n2363), .A0(n2381), .A1(n2283), .B0(n2369) );
  inv02 U1296 ( .Y(n2364), .A(n2363) );
  inv02 U1297 ( .Y(n2460), .A(n2365) );
  nor02 U1298 ( .Y(n2366), .A0(n2283), .A1(n2474) );
  nor02 U1299 ( .Y(n2367), .A0(n2381), .A1(n2474) );
  nor02 U1300 ( .Y(n2365), .A0(n2366), .A1(n2367) );
  inv02 U1301 ( .Y(n2474), .A(n2508) );
  or02 U1302 ( .Y(n2368), .A0(s_state355), .A1(s_count[0]) );
  inv01 U1303 ( .Y(n2369), .A(n2368) );
  inv02 U1304 ( .Y(n2370), .A(n2368) );
  inv02 U1305 ( .Y(n2459), .A(n2490) );
  buf04 U1306 ( .Y(n2371), .A(n2454) );
  buf02 U1307 ( .Y(n2372), .A(L546_26_) );
  inv02 U1308 ( .Y(n2389), .A(s_state) );
  ao21 U1309 ( .Y(n2373), .A0(n2494), .A1(n2282), .B0(n2391) );
  inv02 U1310 ( .Y(n2374), .A(n2373) );
  ao21 U1311 ( .Y(n2375), .A0(n2498), .A1(n2281), .B0(n2391) );
  inv02 U1312 ( .Y(n2376), .A(n2375) );
  ao21 U1313 ( .Y(n2377), .A0(n2503), .A1(n2283), .B0(n2391) );
  inv02 U1314 ( .Y(n2378), .A(n2377) );
  buf04 U1315 ( .Y(n2379), .A(n2477) );
  buf04 U1316 ( .Y(n2380), .A(n2487) );
  buf04 U1317 ( .Y(n2381), .A(n2456) );
  buf16 U1318 ( .Y(n2382), .A(n2394) );
  buf16 U1319 ( .Y(n2383), .A(n2396) );
  buf12 U1320 ( .Y(n2384), .A(n1899) );
  buf16 U1321 ( .Y(n2385), .A(n2452) );
  inv08 U1322 ( .Y(n2512), .A(n2384) );
  inv16 U1323 ( .Y(n2386), .A(n2391) );
  inv08 U1324 ( .Y(n2391), .A(n2371) );
  buf16 U1325 ( .Y(n2387), .A(n2397) );
  buf16 U1326 ( .Y(n2388), .A(n2453) );
  xor2 U1327 ( .Y(sign_o), .A0(sign_dvd_i), .A1(sign_div_i) );
  ao21 U1328 ( .Y(n1767), .A0(s_state), .A1(n2392), .B0(s_state355) );
  or02 U1329 ( .Y(n2392), .A0(n2293), .A1(s_count[0]) );
  and02 U1330 ( .Y(n1766), .A0(n2393), .A1(s_dvd[0]) );
  inv01 U1331 ( .Y(n2398), .A(s_dvd[1]) );
  inv01 U1332 ( .Y(n2400), .A(s_dvd[2]) );
  inv01 U1333 ( .Y(n2402), .A(s_dvd[3]) );
  inv01 U1334 ( .Y(n2404), .A(s_dvd[4]) );
  inv01 U1335 ( .Y(n2406), .A(s_dvd[5]) );
  inv01 U1336 ( .Y(n2408), .A(s_dvd[6]) );
  inv01 U1337 ( .Y(n2410), .A(s_dvd[7]) );
  inv01 U1338 ( .Y(n2412), .A(s_dvd[8]) );
  inv01 U1339 ( .Y(n2414), .A(s_dvd[9]) );
  inv01 U1340 ( .Y(n2416), .A(s_dvd[10]) );
  inv01 U1341 ( .Y(n2418), .A(s_dvd[11]) );
  inv01 U1342 ( .Y(n2420), .A(s_dvd[12]) );
  inv01 U1343 ( .Y(n2422), .A(s_dvd[13]) );
  inv01 U1344 ( .Y(n2424), .A(s_dvd[14]) );
  inv01 U1345 ( .Y(n2426), .A(s_dvd[15]) );
  inv01 U1346 ( .Y(n2428), .A(s_dvd[16]) );
  inv01 U1347 ( .Y(n2430), .A(s_dvd[17]) );
  inv01 U1348 ( .Y(n2432), .A(s_dvd[18]) );
  inv01 U1349 ( .Y(n2434), .A(s_dvd[19]) );
  inv01 U1350 ( .Y(n2436), .A(s_dvd[20]) );
  inv01 U1351 ( .Y(n2438), .A(s_dvd[21]) );
  inv01 U1352 ( .Y(n2440), .A(s_dvd[22]) );
  inv01 U1353 ( .Y(n2442), .A(s_dvd[23]) );
  inv01 U1354 ( .Y(n2444), .A(s_dvd[24]) );
  inv01 U1355 ( .Y(n2447), .A(s_dvd[25]) );
  nand02 U1356 ( .Y(n2396), .A0(n____return556), .A1(n2387) );
  nand02 U1357 ( .Y(n2394), .A0(n2387), .A1(n2451) );
  inv01 U1358 ( .Y(n2395), .A(n____return927_0_) );
  inv01 U1359 ( .Y(n2399), .A(n____return927_1_) );
  inv01 U1360 ( .Y(n2401), .A(n____return927_2_) );
  inv01 U1361 ( .Y(n2403), .A(n____return927_3_) );
  inv01 U1362 ( .Y(n2405), .A(n____return927_4_) );
  inv01 U1363 ( .Y(n2407), .A(n____return927_5_) );
  inv01 U1364 ( .Y(n2409), .A(n____return927_6_) );
  inv01 U1365 ( .Y(n2411), .A(n____return927_7_) );
  inv01 U1366 ( .Y(n2413), .A(n____return927_8_) );
  inv01 U1367 ( .Y(n2415), .A(n____return927_9_) );
  inv01 U1368 ( .Y(n2417), .A(n____return927_10_) );
  inv01 U1369 ( .Y(n2419), .A(n____return927_11_) );
  inv01 U1370 ( .Y(n2421), .A(n____return927_12_) );
  inv01 U1371 ( .Y(n2423), .A(n____return927_13_) );
  inv01 U1372 ( .Y(n2425), .A(n____return927_14_) );
  inv01 U1373 ( .Y(n2427), .A(n____return927_15_) );
  inv01 U1374 ( .Y(n2429), .A(n____return927_16_) );
  inv01 U1375 ( .Y(n2431), .A(n____return927_17_) );
  inv01 U1376 ( .Y(n2433), .A(n____return927_18_) );
  inv01 U1377 ( .Y(n2435), .A(n____return927_19_) );
  inv01 U1378 ( .Y(n2437), .A(n____return927_20_) );
  inv01 U1379 ( .Y(n2439), .A(n____return927_21_) );
  inv01 U1380 ( .Y(n2441), .A(n____return927_22_) );
  inv01 U1381 ( .Y(n2443), .A(n____return927_23_) );
  inv01 U1382 ( .Y(n2445), .A(n____return927_24_) );
  inv01 U1383 ( .Y(n2453), .A(n2270) );
  inv01 U1384 ( .Y(n2448), .A(n____return927_25_) );
  inv01 U1385 ( .Y(n2455), .A(n2385) );
  inv01 U1386 ( .Y(n2451), .A(n____return556) );
  ao21 U1387 ( .Y(n2458), .A0(n2459), .A1(n2460), .B0(n2568) );
  ao21 U1388 ( .Y(n2462), .A0(n2364), .A1(n2459), .B0(n2557) );
  ao21 U1389 ( .Y(n2464), .A0(n2374), .A1(n2460), .B0(n2549) );
  ao21 U1390 ( .Y(n2466), .A0(n2374), .A1(n2364), .B0(n2548) );
  ao21 U1391 ( .Y(n2468), .A0(n2376), .A1(n2460), .B0(n2547) );
  ao21 U1392 ( .Y(n2470), .A0(n2376), .A1(n2364), .B0(n2546) );
  ao21 U1393 ( .Y(n2472), .A0(n2378), .A1(n2460), .B0(n2545) );
  ao21 U1394 ( .Y(n2476), .A0(n2378), .A1(n2364), .B0(n2544) );
  ao21 U1395 ( .Y(n2478), .A0(n2298), .A1(n2459), .B0(n2543) );
  ao21 U1396 ( .Y(n2479), .A0(n2302), .A1(n2459), .B0(n2542) );
  ao21 U1397 ( .Y(n2480), .A0(n2298), .A1(n2374), .B0(n2567) );
  ao21 U1398 ( .Y(n2481), .A0(n2302), .A1(n2374), .B0(n2566) );
  ao21 U1399 ( .Y(n2482), .A0(n2298), .A1(n2376), .B0(n2565) );
  ao21 U1400 ( .Y(n2483), .A0(n2302), .A1(n2376), .B0(n2564) );
  ao21 U1401 ( .Y(n2484), .A0(n2298), .A1(n2378), .B0(n2563) );
  ao21 U1402 ( .Y(n2485), .A0(n2302), .A1(n2378), .B0(n2562) );
  nand02 U1403 ( .Y(n2477), .A0(s_count[3]), .A1(n2486) );
  ao21 U1404 ( .Y(n2488), .A0(n2304), .A1(n2459), .B0(n2561) );
  ao21 U1405 ( .Y(n2489), .A0(n2300), .A1(n2459), .B0(n2560) );
  ao21 U1406 ( .Y(n2491), .A0(n2304), .A1(n2374), .B0(n2559) );
  nand02 U1407 ( .Y(n2463), .A0(n2246), .A1(n2492) );
  ao21 U1408 ( .Y(n2493), .A0(n2300), .A1(n2374), .B0(n2558) );
  nand02 U1409 ( .Y(n2465), .A0(n2248), .A1(n2492) );
  inv01 U1410 ( .Y(n2492), .A(n2494) );
  ao21 U1411 ( .Y(n2495), .A0(n2304), .A1(n2376), .B0(n2556) );
  nand02 U1412 ( .Y(n2467), .A0(n2237), .A1(n2245) );
  ao21 U1413 ( .Y(n2497), .A0(n2300), .A1(n2376), .B0(n2555) );
  inv01 U1414 ( .Y(n2498), .A(n2237) );
  nand02 U1415 ( .Y(n2469), .A0(n2238), .A1(n2248) );
  nor02 U1416 ( .Y(n2496), .A0(n2499), .A1(s_count[1]) );
  ao21 U1417 ( .Y(n2500), .A0(n2304), .A1(n2378), .B0(n2554) );
  nand02 U1418 ( .Y(n2471), .A0(n2230), .A1(n2244) );
  ao21 U1419 ( .Y(n2502), .A0(n2300), .A1(n2378), .B0(n2553) );
  inv01 U1420 ( .Y(n2503), .A(n2501) );
  nand02 U1421 ( .Y(n2487), .A0(s_count[4]), .A1(n2504) );
  nand02 U1422 ( .Y(n2475), .A0(n2501), .A1(n2248) );
  nor02 U1423 ( .Y(n2501), .A0(n2499), .A1(n2505) );
  ao21 U1424 ( .Y(n2507), .A0(n1911), .A1(n2508), .B0(n2552) );
  nand02 U1425 ( .Y(n2457), .A0(n2245), .A1(n2509) );
  ao21 U1426 ( .Y(n2510), .A0(n1911), .A1(n2390), .B0(n2551) );
  inv01 U1427 ( .Y(n2390), .A(n2370) );
  ao21 U1428 ( .Y(n2490), .A0(n2511), .A1(n2282), .B0(n2391) );
  nand02 U1429 ( .Y(n2461), .A0(n2248), .A1(n2509) );
  inv01 U1430 ( .Y(n2509), .A(n2511) );
  aoi21 U1431 ( .Y(n2513), .A0(n2512), .A1(n2282), .B0(n2391) );
  nand02 U1432 ( .Y(n2452), .A0(n2240), .A1(n2283) );
  nand02 U1433 ( .Y(n1685), .A0(n2514), .A1(n2289) );
  nand02 U1434 ( .Y(n1684), .A0(n2515), .A1(n2289) );
  ao22 U1435 ( .Y(n1683), .A0(s_count[2]), .A1(n2391), .B0(sum426_2_), .B1(
        n2516) );
  nand02 U1436 ( .Y(n2454), .A0(n2281), .A1(n2389) );
  nand02 U1437 ( .Y(n1682), .A0(n2517), .A1(n2289) );
  nor02 U1438 ( .Y(n2518), .A0(s_count[0]), .A1(n2293) );
  ao22 U1439 ( .Y(n1681), .A0(n2474), .A1(n2389), .B0(sum426_0_), .B1(n2519)
         );
  ao21 U1440 ( .Y(n2519), .A0(n2387), .A1(n2293), .B0(n2474) );
  nand02 U1441 ( .Y(n2511), .A0(n2499), .A1(n2505) );
  inv01 U1442 ( .Y(n2505), .A(s_count[1]) );
  nand02 U1443 ( .Y(n2456), .A0(n2486), .A1(n2504) );
  inv01 U1444 ( .Y(n2504), .A(s_count[3]) );
  inv01 U1445 ( .Y(n2486), .A(s_count[4]) );
  inv01 U1446 ( .Y(n2397), .A(n2393) );
  nand02 U1447 ( .Y(n2393), .A0(s_state), .A1(n2281) );
  nand02 U1448 ( .Y(n2508), .A0(s_count[0]), .A1(n2281) );
  nand04 U1449 ( .Y(n2523), .A0(n1385), .A1(n1390), .A2(n1807), .A3(n2263) );
  nand04 U1450 ( .Y(n2524), .A0(n2242), .A1(n2250), .A2(n2252), .A3(n2525) );
  nand04 U1451 ( .Y(n2529), .A0(n2580), .A1(n2530), .A2(n2531), .A3(n1909) );
  inv01 U1452 ( .Y(n2531), .A(s_dvdnd_i_29_) );
  inv01 U1453 ( .Y(n2530), .A(s_dvdnd_i_30_) );
  inv01 U1454 ( .Y(n2528), .A(n2229) );
  or03 U1455 ( .Y(n2532), .A0(s_dvdnd_i_37_), .A1(s_dvdnd_i_39_), .A2(
        s_dvdnd_i_38_) );
  nand04 U1456 ( .Y(n2527), .A0(n2533), .A1(n2534), .A2(n2589), .A3(n1907) );
  inv01 U1457 ( .Y(n2534), .A(s_dvdnd_i_41_) );
  inv01 U1458 ( .Y(n2533), .A(s_dvdnd_i_40_) );
  inv01 U1459 ( .Y(n2526), .A(n2227) );
  inv01 U1460 ( .Y(n2535), .A(n2225) );
  nand02 U1461 ( .Y(n2538), .A0(n2579), .A1(n2577) );
  nand03 U1462 ( .Y(n2537), .A0(n2585), .A1(n2583), .A2(n2578) );
  nand04 U1463 ( .Y(n2536), .A0(n2582), .A1(n2581), .A2(n2584), .A3(n2254) );
  nand03 U1464 ( .Y(n2539), .A0(n2575), .A1(n2574), .A2(n1397) );
  nand03 U1465 ( .Y(n2540), .A0(n1405), .A1(n1406), .A2(n1401) );
  nand04 U1466 ( .Y(n2522), .A0(n2569), .A1(n2570), .A2(n2571), .A3(n2261) );
  nand04 U1467 ( .Y(n2521), .A0(n1395), .A1(n1396), .A2(n1394), .A3(n2267) );
  nand04 U1468 ( .Y(n2520), .A0(n1388), .A1(n1389), .A2(n1387), .A3(n2265) );
  nor02 U1469 ( .Y(L546_26_), .A0(n2450), .A1(n2384) );
  inv01 U1470 ( .Y(n2450), .A(s_dvd[26]) );
  nand02 U1471 ( .Y(n2449), .A0(s_dvd[25]), .A1(n2512) );
  nand02 U1472 ( .Y(n2446), .A0(s_dvd[24]), .A1(n2512) );
  nand02 U1473 ( .Y(n2494), .A0(s_count[1]), .A1(n2499) );
  nand02 U1474 ( .Y(n2506), .A0(s_count[4]), .A1(s_count[3]) );
  serial_div_DW01_sub_27_0 sub_154_minus_minus ( .A({n2372, L546_25_, L546_24_, 
        L546_23_, L546_22_, L546_21_, L546_20_, L546_19_, L546_18_, L546_17_, 
        L546_16_, L546_15_, L546_14_, L546_13_, L546_12_, L546_11_, L546_10_, 
        L546_9_, L546_8_, L546_7_, L546_6_, L546_5_, L546_4_, L546_3_, L546_2_, 
        L546_1_, L546_0_}), .B({s_dvsor_i_26_, s_dvsor_i_25_, s_dvsor_i_24_, 
        s_dvsor_i_23_, s_dvsor_i_22_, s_dvsor_i_21_, s_dvsor_i_20_, 
        s_dvsor_i_19_, s_dvsor_i_18_, s_dvsor_i_17_, s_dvsor_i_16_, 
        s_dvsor_i_15_, s_dvsor_i_14_, s_dvsor_i_13_, s_dvsor_i_12_, 
        s_dvsor_i_11_, s_dvsor_i_10_, s_dvsor_i_9_, s_dvsor_i_8_, s_dvsor_i_7_, 
        s_dvsor_i_6_, s_dvsor_i_5_, s_dvsor_i_4_, s_dvsor_i_3_, s_dvsor_i_2_, 
        s_dvsor_i_1_, s_dvsor_i_0_}), .CI(1'b0), .DIFF({n____return927_26_, 
        n____return927_25_, n____return927_24_, n____return927_23_, 
        n____return927_22_, n____return927_21_, n____return927_20_, 
        n____return927_19_, n____return927_18_, n____return927_17_, 
        n____return927_16_, n____return927_15_, n____return927_14_, 
        n____return927_13_, n____return927_12_, n____return927_11_, 
        n____return927_10_, n____return927_9_, n____return927_8_, 
        n____return927_7_, n____return927_6_, n____return927_5_, 
        n____return927_4_, n____return927_3_, n____return927_2_, 
        n____return927_1_, n____return927_0_}) );
  serial_div_DW01_cmp2_27_0 lt_150_lt_lt ( .A({n2372, L546_25_, L546_24_, 
        L546_23_, L546_22_, L546_21_, L546_20_, L546_19_, L546_18_, L546_17_, 
        L546_16_, L546_15_, L546_14_, L546_13_, L546_12_, L546_11_, L546_10_, 
        L546_9_, L546_8_, L546_7_, L546_6_, L546_5_, L546_4_, L546_3_, L546_2_, 
        L546_1_, L546_0_}), .B({s_dvsor_i_26_, s_dvsor_i_25_, s_dvsor_i_24_, 
        s_dvsor_i_23_, s_dvsor_i_22_, s_dvsor_i_21_, s_dvsor_i_20_, 
        s_dvsor_i_19_, s_dvsor_i_18_, s_dvsor_i_17_, s_dvsor_i_16_, 
        s_dvsor_i_15_, s_dvsor_i_14_, s_dvsor_i_13_, s_dvsor_i_12_, 
        s_dvsor_i_11_, s_dvsor_i_10_, s_dvsor_i_9_, s_dvsor_i_8_, s_dvsor_i_7_, 
        s_dvsor_i_6_, s_dvsor_i_5_, s_dvsor_i_4_, s_dvsor_i_3_, s_dvsor_i_2_, 
        s_dvsor_i_1_, s_dvsor_i_0_}), .LEQ(1'b0), .TC(1'b0), .LT_LE(
        n____return556) );
  serial_div_DW01_dec_5_0 sub_127 ( .A({s_count[4:1], n2287}), .SUM({sum426_4_, 
        sum426_3_, sum426_2_, sum426_1_, sum426_0_}) );
endmodule


module sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_inc_52_0 ( A, SUM );
  input [51:0] A;
  output [51:0] SUM;
  wire   n2, carry_51_, carry_50_, carry_49_, carry_48_, carry_47_, carry_46_,
         carry_45_, carry_44_, carry_43_, carry_42_, carry_41_, carry_40_,
         carry_39_, carry_38_, carry_37_, carry_36_, carry_35_, carry_34_,
         carry_33_, carry_32_, carry_31_, carry_30_, carry_29_, carry_28_,
         carry_27_, carry_26_, carry_25_, carry_24_, carry_23_, carry_22_,
         carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, carry_6_, carry_5_, carry_4_, carry_3_,
         carry_2_;

  buf02 U5 ( .Y(SUM[0]), .A(n2) );
  inv01 U6 ( .Y(n2), .A(A[0]) );
  xor2 U7 ( .Y(SUM[51]), .A0(carry_51_), .A1(A[51]) );
  hadd1 U1_1_1 ( .S(SUM[1]), .CO(carry_2_), .A(A[1]), .B(A[0]) );
  hadd1 U1_1_2 ( .S(SUM[2]), .CO(carry_3_), .A(A[2]), .B(carry_2_) );
  hadd1 U1_1_3 ( .S(SUM[3]), .CO(carry_4_), .A(A[3]), .B(carry_3_) );
  hadd1 U1_1_4 ( .S(SUM[4]), .CO(carry_5_), .A(A[4]), .B(carry_4_) );
  hadd1 U1_1_5 ( .S(SUM[5]), .CO(carry_6_), .A(A[5]), .B(carry_5_) );
  hadd1 U1_1_6 ( .S(SUM[6]), .CO(carry_7_), .A(A[6]), .B(carry_6_) );
  hadd1 U1_1_7 ( .S(SUM[7]), .CO(carry_8_), .A(A[7]), .B(carry_7_) );
  hadd1 U1_1_8 ( .S(SUM[8]), .CO(carry_9_), .A(A[8]), .B(carry_8_) );
  hadd1 U1_1_9 ( .S(SUM[9]), .CO(carry_10_), .A(A[9]), .B(carry_9_) );
  hadd1 U1_1_10 ( .S(SUM[10]), .CO(carry_11_), .A(A[10]), .B(carry_10_) );
  hadd1 U1_1_11 ( .S(SUM[11]), .CO(carry_12_), .A(A[11]), .B(carry_11_) );
  hadd1 U1_1_12 ( .S(SUM[12]), .CO(carry_13_), .A(A[12]), .B(carry_12_) );
  hadd1 U1_1_13 ( .S(SUM[13]), .CO(carry_14_), .A(A[13]), .B(carry_13_) );
  hadd1 U1_1_14 ( .S(SUM[14]), .CO(carry_15_), .A(A[14]), .B(carry_14_) );
  hadd1 U1_1_15 ( .S(SUM[15]), .CO(carry_16_), .A(A[15]), .B(carry_15_) );
  hadd1 U1_1_16 ( .S(SUM[16]), .CO(carry_17_), .A(A[16]), .B(carry_16_) );
  hadd1 U1_1_17 ( .S(SUM[17]), .CO(carry_18_), .A(A[17]), .B(carry_17_) );
  hadd1 U1_1_18 ( .S(SUM[18]), .CO(carry_19_), .A(A[18]), .B(carry_18_) );
  hadd1 U1_1_19 ( .S(SUM[19]), .CO(carry_20_), .A(A[19]), .B(carry_19_) );
  hadd1 U1_1_20 ( .S(SUM[20]), .CO(carry_21_), .A(A[20]), .B(carry_20_) );
  hadd1 U1_1_21 ( .S(SUM[21]), .CO(carry_22_), .A(A[21]), .B(carry_21_) );
  hadd1 U1_1_22 ( .S(SUM[22]), .CO(carry_23_), .A(A[22]), .B(carry_22_) );
  hadd1 U1_1_23 ( .S(SUM[23]), .CO(carry_24_), .A(A[23]), .B(carry_23_) );
  hadd1 U1_1_24 ( .S(SUM[24]), .CO(carry_25_), .A(A[24]), .B(carry_24_) );
  hadd1 U1_1_25 ( .S(SUM[25]), .CO(carry_26_), .A(A[25]), .B(carry_25_) );
  hadd1 U1_1_26 ( .S(SUM[26]), .CO(carry_27_), .A(A[26]), .B(carry_26_) );
  hadd1 U1_1_27 ( .S(SUM[27]), .CO(carry_28_), .A(A[27]), .B(carry_27_) );
  hadd1 U1_1_28 ( .S(SUM[28]), .CO(carry_29_), .A(A[28]), .B(carry_28_) );
  hadd1 U1_1_29 ( .S(SUM[29]), .CO(carry_30_), .A(A[29]), .B(carry_29_) );
  hadd1 U1_1_30 ( .S(SUM[30]), .CO(carry_31_), .A(A[30]), .B(carry_30_) );
  hadd1 U1_1_31 ( .S(SUM[31]), .CO(carry_32_), .A(A[31]), .B(carry_31_) );
  hadd1 U1_1_32 ( .S(SUM[32]), .CO(carry_33_), .A(A[32]), .B(carry_32_) );
  hadd1 U1_1_33 ( .S(SUM[33]), .CO(carry_34_), .A(A[33]), .B(carry_33_) );
  hadd1 U1_1_34 ( .S(SUM[34]), .CO(carry_35_), .A(A[34]), .B(carry_34_) );
  hadd1 U1_1_35 ( .S(SUM[35]), .CO(carry_36_), .A(A[35]), .B(carry_35_) );
  hadd1 U1_1_36 ( .S(SUM[36]), .CO(carry_37_), .A(A[36]), .B(carry_36_) );
  hadd1 U1_1_37 ( .S(SUM[37]), .CO(carry_38_), .A(A[37]), .B(carry_37_) );
  hadd1 U1_1_38 ( .S(SUM[38]), .CO(carry_39_), .A(A[38]), .B(carry_38_) );
  hadd1 U1_1_39 ( .S(SUM[39]), .CO(carry_40_), .A(A[39]), .B(carry_39_) );
  hadd1 U1_1_40 ( .S(SUM[40]), .CO(carry_41_), .A(A[40]), .B(carry_40_) );
  hadd1 U1_1_41 ( .S(SUM[41]), .CO(carry_42_), .A(A[41]), .B(carry_41_) );
  hadd1 U1_1_42 ( .S(SUM[42]), .CO(carry_43_), .A(A[42]), .B(carry_42_) );
  hadd1 U1_1_43 ( .S(SUM[43]), .CO(carry_44_), .A(A[43]), .B(carry_43_) );
  hadd1 U1_1_44 ( .S(SUM[44]), .CO(carry_45_), .A(A[44]), .B(carry_44_) );
  hadd1 U1_1_45 ( .S(SUM[45]), .CO(carry_46_), .A(A[45]), .B(carry_45_) );
  hadd1 U1_1_46 ( .S(SUM[46]), .CO(carry_47_), .A(A[46]), .B(carry_46_) );
  hadd1 U1_1_47 ( .S(SUM[47]), .CO(carry_48_), .A(A[47]), .B(carry_47_) );
  hadd1 U1_1_48 ( .S(SUM[48]), .CO(carry_49_), .A(A[48]), .B(carry_48_) );
  hadd1 U1_1_49 ( .S(SUM[49]), .CO(carry_50_), .A(A[49]), .B(carry_49_) );
  hadd1 U1_1_50 ( .S(SUM[50]), .CO(carry_51_), .A(A[50]), .B(carry_50_) );
endmodule


module sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_sub_52_1 ( A, B, CI, DIFF, CO );
  input [51:0] A;
  input [51:0] B;
  output [51:0] DIFF;
  input CI;
  output CO;
  wire   carry_51_, carry_50_, carry_49_, carry_48_, carry_47_, carry_46_,
         carry_45_, carry_44_, carry_43_, carry_42_, carry_41_, carry_40_,
         carry_39_, carry_38_, carry_37_, carry_36_, carry_35_, carry_34_,
         carry_33_, carry_32_, carry_31_, carry_30_, carry_29_, carry_28_,
         carry_27_, carry_26_, carry_25_, carry_24_, carry_23_, carry_22_,
         carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, carry_6_, carry_5_, carry_4_, carry_3_,
         carry_2_, B_not_51_, B_not_50_, B_not_49_, B_not_48_, B_not_47_,
         B_not_46_, B_not_45_, B_not_44_, B_not_43_, B_not_42_, B_not_41_,
         B_not_40_, B_not_39_, B_not_38_, B_not_37_, B_not_36_, B_not_35_,
         B_not_34_, B_not_33_, B_not_32_, B_not_31_, B_not_30_, B_not_29_,
         B_not_28_, B_not_27_, B_not_26_, B_not_25_, B_not_24_, B_not_23_,
         B_not_22_, B_not_21_, B_not_20_, B_not_19_, B_not_18_, B_not_17_,
         B_not_16_, B_not_15_, B_not_14_, B_not_13_, B_not_12_, B_not_11_,
         B_not_10_, B_not_9_, B_not_8_, B_not_7_, B_not_6_, B_not_5_, B_not_4_,
         B_not_3_, B_not_2_, B_not_1_, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, A_0_, n15, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066;
  assign DIFF[0] = A_0_;
  assign A_0_ = A[0];

  buf02 U6 ( .Y(DIFF[19]), .A(n1069) );
  buf02 U7 ( .Y(DIFF[13]), .A(n1072) );
  buf02 U8 ( .Y(DIFF[15]), .A(n1070) );
  buf02 U9 ( .Y(DIFF[7]), .A(n1075) );
  buf02 U10 ( .Y(DIFF[4]), .A(n1076) );
  buf02 U11 ( .Y(DIFF[14]), .A(n1071) );
  buf02 U12 ( .Y(DIFF[9]), .A(n1073) );
  buf02 U13 ( .Y(DIFF[8]), .A(n1074) );
  buf02 U14 ( .Y(DIFF[20]), .A(n1068) );
  buf02 U15 ( .Y(DIFF[51]), .A(n1067) );
  xor2 U16 ( .Y(n15), .A0(B_not_1_), .A1(A[1]) );
  inv01 U17 ( .Y(DIFF[1]), .A(n15) );
  inv01 U18 ( .Y(DIFF[35]), .A(n17) );
  inv02 U19 ( .Y(carry_36_), .A(n18) );
  inv02 U20 ( .Y(n19), .A(B_not_35_) );
  inv02 U21 ( .Y(n20), .A(A[35]) );
  inv02 U22 ( .Y(n21), .A(carry_35_) );
  nor02 U23 ( .Y(n22), .A0(n19), .A1(n23) );
  nor02 U24 ( .Y(n24), .A0(n20), .A1(n25) );
  nor02 U25 ( .Y(n26), .A0(n21), .A1(n27) );
  nor02 U26 ( .Y(n28), .A0(n21), .A1(n29) );
  nor02 U27 ( .Y(n17), .A0(n30), .A1(n31) );
  nor02 U28 ( .Y(n32), .A0(n20), .A1(n21) );
  nor02 U29 ( .Y(n33), .A0(n19), .A1(n21) );
  nor02 U30 ( .Y(n34), .A0(n19), .A1(n20) );
  nor02 U31 ( .Y(n18), .A0(n34), .A1(n35) );
  nor02 U32 ( .Y(n36), .A0(A[35]), .A1(carry_35_) );
  inv01 U33 ( .Y(n23), .A(n36) );
  nor02 U34 ( .Y(n37), .A0(B_not_35_), .A1(carry_35_) );
  inv01 U35 ( .Y(n25), .A(n37) );
  nor02 U36 ( .Y(n38), .A0(B_not_35_), .A1(A[35]) );
  inv01 U37 ( .Y(n27), .A(n38) );
  nor02 U38 ( .Y(n39), .A0(n19), .A1(n20) );
  inv01 U39 ( .Y(n29), .A(n39) );
  nor02 U40 ( .Y(n40), .A0(n22), .A1(n24) );
  inv01 U41 ( .Y(n30), .A(n40) );
  nor02 U42 ( .Y(n41), .A0(n26), .A1(n28) );
  inv01 U43 ( .Y(n31), .A(n41) );
  nor02 U44 ( .Y(n42), .A0(n32), .A1(n33) );
  inv01 U45 ( .Y(n35), .A(n42) );
  inv01 U46 ( .Y(DIFF[29]), .A(n43) );
  inv02 U47 ( .Y(carry_30_), .A(n44) );
  inv02 U48 ( .Y(n45), .A(B_not_29_) );
  inv02 U49 ( .Y(n46), .A(A[29]) );
  inv02 U50 ( .Y(n47), .A(carry_29_) );
  nor02 U51 ( .Y(n48), .A0(n45), .A1(n49) );
  nor02 U52 ( .Y(n50), .A0(n46), .A1(n51) );
  nor02 U53 ( .Y(n52), .A0(n47), .A1(n53) );
  nor02 U54 ( .Y(n54), .A0(n47), .A1(n55) );
  nor02 U55 ( .Y(n43), .A0(n56), .A1(n57) );
  nor02 U56 ( .Y(n58), .A0(n46), .A1(n47) );
  nor02 U57 ( .Y(n59), .A0(n45), .A1(n47) );
  nor02 U58 ( .Y(n60), .A0(n45), .A1(n46) );
  nor02 U59 ( .Y(n44), .A0(n60), .A1(n61) );
  nor02 U60 ( .Y(n62), .A0(A[29]), .A1(carry_29_) );
  inv01 U61 ( .Y(n49), .A(n62) );
  nor02 U62 ( .Y(n63), .A0(B_not_29_), .A1(carry_29_) );
  inv01 U63 ( .Y(n51), .A(n63) );
  nor02 U64 ( .Y(n64), .A0(B_not_29_), .A1(A[29]) );
  inv01 U65 ( .Y(n53), .A(n64) );
  nor02 U66 ( .Y(n65), .A0(n45), .A1(n46) );
  inv01 U67 ( .Y(n55), .A(n65) );
  nor02 U68 ( .Y(n66), .A0(n48), .A1(n50) );
  inv01 U69 ( .Y(n56), .A(n66) );
  nor02 U70 ( .Y(n67), .A0(n52), .A1(n54) );
  inv01 U71 ( .Y(n57), .A(n67) );
  nor02 U72 ( .Y(n68), .A0(n58), .A1(n59) );
  inv01 U73 ( .Y(n61), .A(n68) );
  inv01 U74 ( .Y(DIFF[28]), .A(n69) );
  inv02 U75 ( .Y(carry_29_), .A(n70) );
  inv02 U76 ( .Y(n71), .A(B_not_28_) );
  inv02 U77 ( .Y(n72), .A(A[28]) );
  inv02 U78 ( .Y(n73), .A(carry_28_) );
  nor02 U79 ( .Y(n74), .A0(n71), .A1(n75) );
  nor02 U80 ( .Y(n76), .A0(n72), .A1(n77) );
  nor02 U81 ( .Y(n78), .A0(n73), .A1(n79) );
  nor02 U82 ( .Y(n80), .A0(n73), .A1(n81) );
  nor02 U83 ( .Y(n69), .A0(n82), .A1(n83) );
  nor02 U84 ( .Y(n84), .A0(n72), .A1(n73) );
  nor02 U85 ( .Y(n85), .A0(n71), .A1(n73) );
  nor02 U86 ( .Y(n86), .A0(n71), .A1(n72) );
  nor02 U87 ( .Y(n70), .A0(n86), .A1(n87) );
  nor02 U88 ( .Y(n88), .A0(A[28]), .A1(carry_28_) );
  inv01 U89 ( .Y(n75), .A(n88) );
  nor02 U90 ( .Y(n89), .A0(B_not_28_), .A1(carry_28_) );
  inv01 U91 ( .Y(n77), .A(n89) );
  nor02 U92 ( .Y(n90), .A0(B_not_28_), .A1(A[28]) );
  inv01 U93 ( .Y(n79), .A(n90) );
  nor02 U94 ( .Y(n91), .A0(n71), .A1(n72) );
  inv01 U95 ( .Y(n81), .A(n91) );
  nor02 U96 ( .Y(n92), .A0(n74), .A1(n76) );
  inv01 U97 ( .Y(n82), .A(n92) );
  nor02 U98 ( .Y(n93), .A0(n78), .A1(n80) );
  inv01 U99 ( .Y(n83), .A(n93) );
  nor02 U100 ( .Y(n94), .A0(n84), .A1(n85) );
  inv01 U101 ( .Y(n87), .A(n94) );
  inv02 U102 ( .Y(B_not_35_), .A(B[35]) );
  inv02 U103 ( .Y(B_not_29_), .A(B[29]) );
  inv02 U104 ( .Y(B_not_28_), .A(B[28]) );
  inv01 U105 ( .Y(DIFF[36]), .A(n95) );
  inv02 U106 ( .Y(carry_37_), .A(n96) );
  inv02 U107 ( .Y(n97), .A(B_not_36_) );
  inv02 U108 ( .Y(n98), .A(A[36]) );
  inv02 U109 ( .Y(n99), .A(carry_36_) );
  nor02 U110 ( .Y(n100), .A0(n97), .A1(n101) );
  nor02 U111 ( .Y(n102), .A0(n98), .A1(n103) );
  nor02 U112 ( .Y(n104), .A0(n99), .A1(n105) );
  nor02 U113 ( .Y(n106), .A0(n99), .A1(n107) );
  nor02 U114 ( .Y(n95), .A0(n108), .A1(n109) );
  nor02 U115 ( .Y(n110), .A0(n98), .A1(n99) );
  nor02 U116 ( .Y(n111), .A0(n97), .A1(n99) );
  nor02 U117 ( .Y(n112), .A0(n97), .A1(n98) );
  nor02 U118 ( .Y(n96), .A0(n112), .A1(n113) );
  nor02 U119 ( .Y(n114), .A0(A[36]), .A1(carry_36_) );
  inv01 U120 ( .Y(n101), .A(n114) );
  nor02 U121 ( .Y(n115), .A0(B_not_36_), .A1(carry_36_) );
  inv01 U122 ( .Y(n103), .A(n115) );
  nor02 U123 ( .Y(n116), .A0(B_not_36_), .A1(A[36]) );
  inv01 U124 ( .Y(n105), .A(n116) );
  nor02 U125 ( .Y(n117), .A0(n97), .A1(n98) );
  inv01 U126 ( .Y(n107), .A(n117) );
  nor02 U127 ( .Y(n118), .A0(n100), .A1(n102) );
  inv01 U128 ( .Y(n108), .A(n118) );
  nor02 U129 ( .Y(n119), .A0(n104), .A1(n106) );
  inv01 U130 ( .Y(n109), .A(n119) );
  nor02 U131 ( .Y(n120), .A0(n110), .A1(n111) );
  inv01 U132 ( .Y(n113), .A(n120) );
  inv01 U133 ( .Y(DIFF[30]), .A(n121) );
  inv02 U134 ( .Y(carry_31_), .A(n122) );
  inv02 U135 ( .Y(n123), .A(B_not_30_) );
  inv02 U136 ( .Y(n124), .A(A[30]) );
  inv02 U137 ( .Y(n125), .A(carry_30_) );
  nor02 U138 ( .Y(n126), .A0(n123), .A1(n127) );
  nor02 U139 ( .Y(n128), .A0(n124), .A1(n129) );
  nor02 U140 ( .Y(n130), .A0(n125), .A1(n131) );
  nor02 U141 ( .Y(n132), .A0(n125), .A1(n133) );
  nor02 U142 ( .Y(n121), .A0(n134), .A1(n135) );
  nor02 U143 ( .Y(n136), .A0(n124), .A1(n125) );
  nor02 U144 ( .Y(n137), .A0(n123), .A1(n125) );
  nor02 U145 ( .Y(n138), .A0(n123), .A1(n124) );
  nor02 U146 ( .Y(n122), .A0(n138), .A1(n139) );
  nor02 U147 ( .Y(n140), .A0(A[30]), .A1(carry_30_) );
  inv01 U148 ( .Y(n127), .A(n140) );
  nor02 U149 ( .Y(n141), .A0(B_not_30_), .A1(carry_30_) );
  inv01 U150 ( .Y(n129), .A(n141) );
  nor02 U151 ( .Y(n142), .A0(B_not_30_), .A1(A[30]) );
  inv01 U152 ( .Y(n131), .A(n142) );
  nor02 U153 ( .Y(n143), .A0(n123), .A1(n124) );
  inv01 U154 ( .Y(n133), .A(n143) );
  nor02 U155 ( .Y(n144), .A0(n126), .A1(n128) );
  inv01 U156 ( .Y(n134), .A(n144) );
  nor02 U157 ( .Y(n145), .A0(n130), .A1(n132) );
  inv01 U158 ( .Y(n135), .A(n145) );
  nor02 U159 ( .Y(n146), .A0(n136), .A1(n137) );
  inv01 U160 ( .Y(n139), .A(n146) );
  inv01 U161 ( .Y(DIFF[34]), .A(n147) );
  inv02 U162 ( .Y(carry_35_), .A(n148) );
  inv02 U163 ( .Y(n149), .A(B_not_34_) );
  inv02 U164 ( .Y(n150), .A(A[34]) );
  inv02 U165 ( .Y(n151), .A(carry_34_) );
  nor02 U166 ( .Y(n152), .A0(n149), .A1(n153) );
  nor02 U167 ( .Y(n154), .A0(n150), .A1(n155) );
  nor02 U168 ( .Y(n156), .A0(n151), .A1(n157) );
  nor02 U169 ( .Y(n158), .A0(n151), .A1(n159) );
  nor02 U170 ( .Y(n147), .A0(n160), .A1(n161) );
  nor02 U171 ( .Y(n162), .A0(n150), .A1(n151) );
  nor02 U172 ( .Y(n163), .A0(n149), .A1(n151) );
  nor02 U173 ( .Y(n164), .A0(n149), .A1(n150) );
  nor02 U174 ( .Y(n148), .A0(n164), .A1(n165) );
  nor02 U175 ( .Y(n166), .A0(A[34]), .A1(carry_34_) );
  inv01 U176 ( .Y(n153), .A(n166) );
  nor02 U177 ( .Y(n167), .A0(B_not_34_), .A1(carry_34_) );
  inv01 U178 ( .Y(n155), .A(n167) );
  nor02 U179 ( .Y(n168), .A0(B_not_34_), .A1(A[34]) );
  inv01 U180 ( .Y(n157), .A(n168) );
  nor02 U181 ( .Y(n169), .A0(n149), .A1(n150) );
  inv01 U182 ( .Y(n159), .A(n169) );
  nor02 U183 ( .Y(n170), .A0(n152), .A1(n154) );
  inv01 U184 ( .Y(n160), .A(n170) );
  nor02 U185 ( .Y(n171), .A0(n156), .A1(n158) );
  inv01 U186 ( .Y(n161), .A(n171) );
  nor02 U187 ( .Y(n172), .A0(n162), .A1(n163) );
  inv01 U188 ( .Y(n165), .A(n172) );
  inv02 U189 ( .Y(B_not_36_), .A(B[36]) );
  inv02 U190 ( .Y(B_not_30_), .A(B[30]) );
  inv02 U191 ( .Y(B_not_34_), .A(B[34]) );
  inv01 U192 ( .Y(DIFF[37]), .A(n173) );
  inv02 U193 ( .Y(carry_38_), .A(n174) );
  inv02 U194 ( .Y(n175), .A(B_not_37_) );
  inv02 U195 ( .Y(n176), .A(A[37]) );
  inv02 U196 ( .Y(n177), .A(carry_37_) );
  nor02 U197 ( .Y(n178), .A0(n175), .A1(n179) );
  nor02 U198 ( .Y(n180), .A0(n176), .A1(n181) );
  nor02 U199 ( .Y(n182), .A0(n177), .A1(n183) );
  nor02 U200 ( .Y(n184), .A0(n177), .A1(n185) );
  nor02 U201 ( .Y(n173), .A0(n186), .A1(n187) );
  nor02 U202 ( .Y(n188), .A0(n176), .A1(n177) );
  nor02 U203 ( .Y(n189), .A0(n175), .A1(n177) );
  nor02 U204 ( .Y(n190), .A0(n175), .A1(n176) );
  nor02 U205 ( .Y(n174), .A0(n190), .A1(n191) );
  nor02 U206 ( .Y(n192), .A0(A[37]), .A1(carry_37_) );
  inv01 U207 ( .Y(n179), .A(n192) );
  nor02 U208 ( .Y(n193), .A0(B_not_37_), .A1(carry_37_) );
  inv01 U209 ( .Y(n181), .A(n193) );
  nor02 U210 ( .Y(n194), .A0(B_not_37_), .A1(A[37]) );
  inv01 U211 ( .Y(n183), .A(n194) );
  nor02 U212 ( .Y(n195), .A0(n175), .A1(n176) );
  inv01 U213 ( .Y(n185), .A(n195) );
  nor02 U214 ( .Y(n196), .A0(n178), .A1(n180) );
  inv01 U215 ( .Y(n186), .A(n196) );
  nor02 U216 ( .Y(n197), .A0(n182), .A1(n184) );
  inv01 U217 ( .Y(n187), .A(n197) );
  nor02 U218 ( .Y(n198), .A0(n188), .A1(n189) );
  inv01 U219 ( .Y(n191), .A(n198) );
  inv01 U220 ( .Y(DIFF[31]), .A(n199) );
  inv02 U221 ( .Y(carry_32_), .A(n200) );
  inv02 U222 ( .Y(n201), .A(B_not_31_) );
  inv02 U223 ( .Y(n202), .A(A[31]) );
  inv02 U224 ( .Y(n203), .A(carry_31_) );
  nor02 U225 ( .Y(n204), .A0(n201), .A1(n205) );
  nor02 U226 ( .Y(n206), .A0(n202), .A1(n207) );
  nor02 U227 ( .Y(n208), .A0(n203), .A1(n209) );
  nor02 U228 ( .Y(n210), .A0(n203), .A1(n211) );
  nor02 U229 ( .Y(n199), .A0(n212), .A1(n213) );
  nor02 U230 ( .Y(n214), .A0(n202), .A1(n203) );
  nor02 U231 ( .Y(n215), .A0(n201), .A1(n203) );
  nor02 U232 ( .Y(n216), .A0(n201), .A1(n202) );
  nor02 U233 ( .Y(n200), .A0(n216), .A1(n217) );
  nor02 U234 ( .Y(n218), .A0(A[31]), .A1(carry_31_) );
  inv01 U235 ( .Y(n205), .A(n218) );
  nor02 U236 ( .Y(n219), .A0(B_not_31_), .A1(carry_31_) );
  inv01 U237 ( .Y(n207), .A(n219) );
  nor02 U238 ( .Y(n220), .A0(B_not_31_), .A1(A[31]) );
  inv01 U239 ( .Y(n209), .A(n220) );
  nor02 U240 ( .Y(n221), .A0(n201), .A1(n202) );
  inv01 U241 ( .Y(n211), .A(n221) );
  nor02 U242 ( .Y(n222), .A0(n204), .A1(n206) );
  inv01 U243 ( .Y(n212), .A(n222) );
  nor02 U244 ( .Y(n223), .A0(n208), .A1(n210) );
  inv01 U245 ( .Y(n213), .A(n223) );
  nor02 U246 ( .Y(n224), .A0(n214), .A1(n215) );
  inv01 U247 ( .Y(n217), .A(n224) );
  inv01 U248 ( .Y(DIFF[33]), .A(n225) );
  inv02 U249 ( .Y(carry_34_), .A(n226) );
  inv02 U250 ( .Y(n227), .A(B_not_33_) );
  inv02 U251 ( .Y(n228), .A(A[33]) );
  inv02 U252 ( .Y(n229), .A(carry_33_) );
  nor02 U253 ( .Y(n230), .A0(n227), .A1(n231) );
  nor02 U254 ( .Y(n232), .A0(n228), .A1(n233) );
  nor02 U255 ( .Y(n234), .A0(n229), .A1(n235) );
  nor02 U256 ( .Y(n236), .A0(n229), .A1(n237) );
  nor02 U257 ( .Y(n225), .A0(n238), .A1(n239) );
  nor02 U258 ( .Y(n240), .A0(n228), .A1(n229) );
  nor02 U259 ( .Y(n241), .A0(n227), .A1(n229) );
  nor02 U260 ( .Y(n242), .A0(n227), .A1(n228) );
  nor02 U261 ( .Y(n226), .A0(n242), .A1(n243) );
  nor02 U262 ( .Y(n244), .A0(A[33]), .A1(carry_33_) );
  inv01 U263 ( .Y(n231), .A(n244) );
  nor02 U264 ( .Y(n245), .A0(B_not_33_), .A1(carry_33_) );
  inv01 U265 ( .Y(n233), .A(n245) );
  nor02 U266 ( .Y(n246), .A0(B_not_33_), .A1(A[33]) );
  inv01 U267 ( .Y(n235), .A(n246) );
  nor02 U268 ( .Y(n247), .A0(n227), .A1(n228) );
  inv01 U269 ( .Y(n237), .A(n247) );
  nor02 U270 ( .Y(n248), .A0(n230), .A1(n232) );
  inv01 U271 ( .Y(n238), .A(n248) );
  nor02 U272 ( .Y(n249), .A0(n234), .A1(n236) );
  inv01 U273 ( .Y(n239), .A(n249) );
  nor02 U274 ( .Y(n250), .A0(n240), .A1(n241) );
  inv01 U275 ( .Y(n243), .A(n250) );
  inv02 U276 ( .Y(B_not_37_), .A(B[37]) );
  inv02 U277 ( .Y(B_not_31_), .A(B[31]) );
  inv02 U278 ( .Y(B_not_33_), .A(B[33]) );
  inv01 U279 ( .Y(DIFF[38]), .A(n251) );
  inv02 U280 ( .Y(carry_39_), .A(n252) );
  inv02 U281 ( .Y(n253), .A(B_not_38_) );
  inv02 U282 ( .Y(n254), .A(A[38]) );
  inv02 U283 ( .Y(n255), .A(carry_38_) );
  nor02 U284 ( .Y(n256), .A0(n253), .A1(n257) );
  nor02 U285 ( .Y(n258), .A0(n254), .A1(n259) );
  nor02 U286 ( .Y(n260), .A0(n255), .A1(n261) );
  nor02 U287 ( .Y(n262), .A0(n255), .A1(n263) );
  nor02 U288 ( .Y(n251), .A0(n264), .A1(n265) );
  nor02 U289 ( .Y(n266), .A0(n254), .A1(n255) );
  nor02 U290 ( .Y(n267), .A0(n253), .A1(n255) );
  nor02 U291 ( .Y(n268), .A0(n253), .A1(n254) );
  nor02 U292 ( .Y(n252), .A0(n268), .A1(n269) );
  nor02 U293 ( .Y(n270), .A0(A[38]), .A1(carry_38_) );
  inv01 U294 ( .Y(n257), .A(n270) );
  nor02 U295 ( .Y(n271), .A0(B_not_38_), .A1(carry_38_) );
  inv01 U296 ( .Y(n259), .A(n271) );
  nor02 U297 ( .Y(n272), .A0(B_not_38_), .A1(A[38]) );
  inv01 U298 ( .Y(n261), .A(n272) );
  nor02 U299 ( .Y(n273), .A0(n253), .A1(n254) );
  inv01 U300 ( .Y(n263), .A(n273) );
  nor02 U301 ( .Y(n274), .A0(n256), .A1(n258) );
  inv01 U302 ( .Y(n264), .A(n274) );
  nor02 U303 ( .Y(n275), .A0(n260), .A1(n262) );
  inv01 U304 ( .Y(n265), .A(n275) );
  nor02 U305 ( .Y(n276), .A0(n266), .A1(n267) );
  inv01 U306 ( .Y(n269), .A(n276) );
  inv01 U307 ( .Y(DIFF[27]), .A(n277) );
  inv02 U308 ( .Y(carry_28_), .A(n278) );
  inv02 U309 ( .Y(n279), .A(B_not_27_) );
  inv02 U310 ( .Y(n280), .A(A[27]) );
  inv02 U311 ( .Y(n281), .A(carry_27_) );
  nor02 U312 ( .Y(n282), .A0(n279), .A1(n283) );
  nor02 U313 ( .Y(n284), .A0(n280), .A1(n285) );
  nor02 U314 ( .Y(n286), .A0(n281), .A1(n287) );
  nor02 U315 ( .Y(n288), .A0(n281), .A1(n289) );
  nor02 U316 ( .Y(n277), .A0(n290), .A1(n291) );
  nor02 U317 ( .Y(n292), .A0(n280), .A1(n281) );
  nor02 U318 ( .Y(n293), .A0(n279), .A1(n281) );
  nor02 U319 ( .Y(n294), .A0(n279), .A1(n280) );
  nor02 U320 ( .Y(n278), .A0(n294), .A1(n295) );
  nor02 U321 ( .Y(n296), .A0(A[27]), .A1(carry_27_) );
  inv01 U322 ( .Y(n283), .A(n296) );
  nor02 U323 ( .Y(n297), .A0(B_not_27_), .A1(carry_27_) );
  inv01 U324 ( .Y(n285), .A(n297) );
  nor02 U325 ( .Y(n298), .A0(B_not_27_), .A1(A[27]) );
  inv01 U326 ( .Y(n287), .A(n298) );
  nor02 U327 ( .Y(n299), .A0(n279), .A1(n280) );
  inv01 U328 ( .Y(n289), .A(n299) );
  nor02 U329 ( .Y(n300), .A0(n282), .A1(n284) );
  inv01 U330 ( .Y(n290), .A(n300) );
  nor02 U331 ( .Y(n301), .A0(n286), .A1(n288) );
  inv01 U332 ( .Y(n291), .A(n301) );
  nor02 U333 ( .Y(n302), .A0(n292), .A1(n293) );
  inv01 U334 ( .Y(n295), .A(n302) );
  inv01 U335 ( .Y(DIFF[32]), .A(n303) );
  inv02 U336 ( .Y(carry_33_), .A(n304) );
  inv02 U337 ( .Y(n305), .A(B_not_32_) );
  inv02 U338 ( .Y(n306), .A(A[32]) );
  inv02 U339 ( .Y(n307), .A(carry_32_) );
  nor02 U340 ( .Y(n308), .A0(n305), .A1(n309) );
  nor02 U341 ( .Y(n310), .A0(n306), .A1(n311) );
  nor02 U342 ( .Y(n312), .A0(n307), .A1(n313) );
  nor02 U343 ( .Y(n314), .A0(n307), .A1(n315) );
  nor02 U344 ( .Y(n303), .A0(n316), .A1(n317) );
  nor02 U345 ( .Y(n318), .A0(n306), .A1(n307) );
  nor02 U346 ( .Y(n319), .A0(n305), .A1(n307) );
  nor02 U347 ( .Y(n320), .A0(n305), .A1(n306) );
  nor02 U348 ( .Y(n304), .A0(n320), .A1(n321) );
  nor02 U349 ( .Y(n322), .A0(A[32]), .A1(carry_32_) );
  inv01 U350 ( .Y(n309), .A(n322) );
  nor02 U351 ( .Y(n323), .A0(B_not_32_), .A1(carry_32_) );
  inv01 U352 ( .Y(n311), .A(n323) );
  nor02 U353 ( .Y(n324), .A0(B_not_32_), .A1(A[32]) );
  inv01 U354 ( .Y(n313), .A(n324) );
  nor02 U355 ( .Y(n325), .A0(n305), .A1(n306) );
  inv01 U356 ( .Y(n315), .A(n325) );
  nor02 U357 ( .Y(n326), .A0(n308), .A1(n310) );
  inv01 U358 ( .Y(n316), .A(n326) );
  nor02 U359 ( .Y(n327), .A0(n312), .A1(n314) );
  inv01 U360 ( .Y(n317), .A(n327) );
  nor02 U361 ( .Y(n328), .A0(n318), .A1(n319) );
  inv01 U362 ( .Y(n321), .A(n328) );
  inv02 U363 ( .Y(B_not_38_), .A(B[38]) );
  inv02 U364 ( .Y(B_not_27_), .A(B[27]) );
  inv02 U365 ( .Y(B_not_32_), .A(B[32]) );
  inv01 U366 ( .Y(DIFF[39]), .A(n329) );
  inv02 U367 ( .Y(carry_40_), .A(n330) );
  inv02 U368 ( .Y(n331), .A(B_not_39_) );
  inv02 U369 ( .Y(n332), .A(A[39]) );
  inv02 U370 ( .Y(n333), .A(carry_39_) );
  nor02 U371 ( .Y(n334), .A0(n331), .A1(n335) );
  nor02 U372 ( .Y(n336), .A0(n332), .A1(n337) );
  nor02 U373 ( .Y(n338), .A0(n333), .A1(n339) );
  nor02 U374 ( .Y(n340), .A0(n333), .A1(n341) );
  nor02 U375 ( .Y(n329), .A0(n342), .A1(n343) );
  nor02 U376 ( .Y(n344), .A0(n332), .A1(n333) );
  nor02 U377 ( .Y(n345), .A0(n331), .A1(n333) );
  nor02 U378 ( .Y(n346), .A0(n331), .A1(n332) );
  nor02 U379 ( .Y(n330), .A0(n346), .A1(n347) );
  nor02 U380 ( .Y(n348), .A0(A[39]), .A1(carry_39_) );
  inv01 U381 ( .Y(n335), .A(n348) );
  nor02 U382 ( .Y(n349), .A0(B_not_39_), .A1(carry_39_) );
  inv01 U383 ( .Y(n337), .A(n349) );
  nor02 U384 ( .Y(n350), .A0(B_not_39_), .A1(A[39]) );
  inv01 U385 ( .Y(n339), .A(n350) );
  nor02 U386 ( .Y(n351), .A0(n331), .A1(n332) );
  inv01 U387 ( .Y(n341), .A(n351) );
  nor02 U388 ( .Y(n352), .A0(n334), .A1(n336) );
  inv01 U389 ( .Y(n342), .A(n352) );
  nor02 U390 ( .Y(n353), .A0(n338), .A1(n340) );
  inv01 U391 ( .Y(n343), .A(n353) );
  nor02 U392 ( .Y(n354), .A0(n344), .A1(n345) );
  inv01 U393 ( .Y(n347), .A(n354) );
  inv01 U394 ( .Y(DIFF[26]), .A(n355) );
  inv02 U395 ( .Y(carry_27_), .A(n356) );
  inv02 U396 ( .Y(n357), .A(B_not_26_) );
  inv02 U397 ( .Y(n358), .A(A[26]) );
  inv02 U398 ( .Y(n359), .A(carry_26_) );
  nor02 U399 ( .Y(n360), .A0(n357), .A1(n361) );
  nor02 U400 ( .Y(n362), .A0(n358), .A1(n363) );
  nor02 U401 ( .Y(n364), .A0(n359), .A1(n365) );
  nor02 U402 ( .Y(n366), .A0(n359), .A1(n367) );
  nor02 U403 ( .Y(n355), .A0(n368), .A1(n369) );
  nor02 U404 ( .Y(n370), .A0(n358), .A1(n359) );
  nor02 U405 ( .Y(n371), .A0(n357), .A1(n359) );
  nor02 U406 ( .Y(n372), .A0(n357), .A1(n358) );
  nor02 U407 ( .Y(n356), .A0(n372), .A1(n373) );
  nor02 U408 ( .Y(n374), .A0(A[26]), .A1(carry_26_) );
  inv01 U409 ( .Y(n361), .A(n374) );
  nor02 U410 ( .Y(n375), .A0(B_not_26_), .A1(carry_26_) );
  inv01 U411 ( .Y(n363), .A(n375) );
  nor02 U412 ( .Y(n376), .A0(B_not_26_), .A1(A[26]) );
  inv01 U413 ( .Y(n365), .A(n376) );
  nor02 U414 ( .Y(n377), .A0(n357), .A1(n358) );
  inv01 U415 ( .Y(n367), .A(n377) );
  nor02 U416 ( .Y(n378), .A0(n360), .A1(n362) );
  inv01 U417 ( .Y(n368), .A(n378) );
  nor02 U418 ( .Y(n379), .A0(n364), .A1(n366) );
  inv01 U419 ( .Y(n369), .A(n379) );
  nor02 U420 ( .Y(n380), .A0(n370), .A1(n371) );
  inv01 U421 ( .Y(n373), .A(n380) );
  inv02 U422 ( .Y(B_not_39_), .A(B[39]) );
  inv02 U423 ( .Y(B_not_26_), .A(B[26]) );
  inv01 U424 ( .Y(DIFF[40]), .A(n381) );
  inv02 U425 ( .Y(carry_41_), .A(n382) );
  inv02 U426 ( .Y(n383), .A(B_not_40_) );
  inv02 U427 ( .Y(n384), .A(A[40]) );
  inv02 U428 ( .Y(n385), .A(carry_40_) );
  nor02 U429 ( .Y(n386), .A0(n383), .A1(n387) );
  nor02 U430 ( .Y(n388), .A0(n384), .A1(n389) );
  nor02 U431 ( .Y(n390), .A0(n385), .A1(n391) );
  nor02 U432 ( .Y(n392), .A0(n385), .A1(n393) );
  nor02 U433 ( .Y(n381), .A0(n394), .A1(n395) );
  nor02 U434 ( .Y(n396), .A0(n384), .A1(n385) );
  nor02 U435 ( .Y(n397), .A0(n383), .A1(n385) );
  nor02 U436 ( .Y(n398), .A0(n383), .A1(n384) );
  nor02 U437 ( .Y(n382), .A0(n398), .A1(n399) );
  nor02 U438 ( .Y(n400), .A0(A[40]), .A1(carry_40_) );
  inv01 U439 ( .Y(n387), .A(n400) );
  nor02 U440 ( .Y(n401), .A0(B_not_40_), .A1(carry_40_) );
  inv01 U441 ( .Y(n389), .A(n401) );
  nor02 U442 ( .Y(n402), .A0(B_not_40_), .A1(A[40]) );
  inv01 U443 ( .Y(n391), .A(n402) );
  nor02 U444 ( .Y(n403), .A0(n383), .A1(n384) );
  inv01 U445 ( .Y(n393), .A(n403) );
  nor02 U446 ( .Y(n404), .A0(n386), .A1(n388) );
  inv01 U447 ( .Y(n394), .A(n404) );
  nor02 U448 ( .Y(n405), .A0(n390), .A1(n392) );
  inv01 U449 ( .Y(n395), .A(n405) );
  nor02 U450 ( .Y(n406), .A0(n396), .A1(n397) );
  inv01 U451 ( .Y(n399), .A(n406) );
  inv01 U452 ( .Y(DIFF[25]), .A(n407) );
  inv02 U453 ( .Y(carry_26_), .A(n408) );
  inv02 U454 ( .Y(n409), .A(B_not_25_) );
  inv02 U455 ( .Y(n410), .A(A[25]) );
  inv02 U456 ( .Y(n411), .A(carry_25_) );
  nor02 U457 ( .Y(n412), .A0(n409), .A1(n413) );
  nor02 U458 ( .Y(n414), .A0(n410), .A1(n415) );
  nor02 U459 ( .Y(n416), .A0(n411), .A1(n417) );
  nor02 U460 ( .Y(n418), .A0(n411), .A1(n419) );
  nor02 U461 ( .Y(n407), .A0(n420), .A1(n421) );
  nor02 U462 ( .Y(n422), .A0(n410), .A1(n411) );
  nor02 U463 ( .Y(n423), .A0(n409), .A1(n411) );
  nor02 U464 ( .Y(n424), .A0(n409), .A1(n410) );
  nor02 U465 ( .Y(n408), .A0(n424), .A1(n425) );
  nor02 U466 ( .Y(n426), .A0(A[25]), .A1(carry_25_) );
  inv01 U467 ( .Y(n413), .A(n426) );
  nor02 U468 ( .Y(n427), .A0(B_not_25_), .A1(carry_25_) );
  inv01 U469 ( .Y(n415), .A(n427) );
  nor02 U470 ( .Y(n428), .A0(B_not_25_), .A1(A[25]) );
  inv01 U471 ( .Y(n417), .A(n428) );
  nor02 U472 ( .Y(n429), .A0(n409), .A1(n410) );
  inv01 U473 ( .Y(n419), .A(n429) );
  nor02 U474 ( .Y(n430), .A0(n412), .A1(n414) );
  inv01 U475 ( .Y(n420), .A(n430) );
  nor02 U476 ( .Y(n431), .A0(n416), .A1(n418) );
  inv01 U477 ( .Y(n421), .A(n431) );
  nor02 U478 ( .Y(n432), .A0(n422), .A1(n423) );
  inv01 U479 ( .Y(n425), .A(n432) );
  inv02 U480 ( .Y(B_not_40_), .A(B[40]) );
  inv02 U481 ( .Y(B_not_25_), .A(B[25]) );
  inv01 U482 ( .Y(DIFF[41]), .A(n433) );
  inv02 U483 ( .Y(carry_42_), .A(n434) );
  inv02 U484 ( .Y(n435), .A(B_not_41_) );
  inv02 U485 ( .Y(n436), .A(A[41]) );
  inv02 U486 ( .Y(n437), .A(carry_41_) );
  nor02 U487 ( .Y(n438), .A0(n435), .A1(n439) );
  nor02 U488 ( .Y(n440), .A0(n436), .A1(n441) );
  nor02 U489 ( .Y(n442), .A0(n437), .A1(n443) );
  nor02 U490 ( .Y(n444), .A0(n437), .A1(n445) );
  nor02 U491 ( .Y(n433), .A0(n446), .A1(n447) );
  nor02 U492 ( .Y(n448), .A0(n436), .A1(n437) );
  nor02 U493 ( .Y(n449), .A0(n435), .A1(n437) );
  nor02 U494 ( .Y(n450), .A0(n435), .A1(n436) );
  nor02 U495 ( .Y(n434), .A0(n450), .A1(n451) );
  nor02 U496 ( .Y(n452), .A0(A[41]), .A1(carry_41_) );
  inv01 U497 ( .Y(n439), .A(n452) );
  nor02 U498 ( .Y(n453), .A0(B_not_41_), .A1(carry_41_) );
  inv01 U499 ( .Y(n441), .A(n453) );
  nor02 U500 ( .Y(n454), .A0(B_not_41_), .A1(A[41]) );
  inv01 U501 ( .Y(n443), .A(n454) );
  nor02 U502 ( .Y(n455), .A0(n435), .A1(n436) );
  inv01 U503 ( .Y(n445), .A(n455) );
  nor02 U504 ( .Y(n456), .A0(n438), .A1(n440) );
  inv01 U505 ( .Y(n446), .A(n456) );
  nor02 U506 ( .Y(n457), .A0(n442), .A1(n444) );
  inv01 U507 ( .Y(n447), .A(n457) );
  nor02 U508 ( .Y(n458), .A0(n448), .A1(n449) );
  inv01 U509 ( .Y(n451), .A(n458) );
  inv01 U510 ( .Y(DIFF[24]), .A(n459) );
  inv02 U511 ( .Y(carry_25_), .A(n460) );
  inv02 U512 ( .Y(n461), .A(B_not_24_) );
  inv02 U513 ( .Y(n462), .A(A[24]) );
  inv02 U514 ( .Y(n463), .A(carry_24_) );
  nor02 U515 ( .Y(n464), .A0(n461), .A1(n465) );
  nor02 U516 ( .Y(n466), .A0(n462), .A1(n467) );
  nor02 U517 ( .Y(n468), .A0(n463), .A1(n469) );
  nor02 U518 ( .Y(n470), .A0(n463), .A1(n471) );
  nor02 U519 ( .Y(n459), .A0(n472), .A1(n473) );
  nor02 U520 ( .Y(n474), .A0(n462), .A1(n463) );
  nor02 U521 ( .Y(n475), .A0(n461), .A1(n463) );
  nor02 U522 ( .Y(n476), .A0(n461), .A1(n462) );
  nor02 U523 ( .Y(n460), .A0(n476), .A1(n477) );
  nor02 U524 ( .Y(n478), .A0(A[24]), .A1(carry_24_) );
  inv01 U525 ( .Y(n465), .A(n478) );
  nor02 U526 ( .Y(n479), .A0(B_not_24_), .A1(carry_24_) );
  inv01 U527 ( .Y(n467), .A(n479) );
  nor02 U528 ( .Y(n480), .A0(B_not_24_), .A1(A[24]) );
  inv01 U529 ( .Y(n469), .A(n480) );
  nor02 U530 ( .Y(n481), .A0(n461), .A1(n462) );
  inv01 U531 ( .Y(n471), .A(n481) );
  nor02 U532 ( .Y(n482), .A0(n464), .A1(n466) );
  inv01 U533 ( .Y(n472), .A(n482) );
  nor02 U534 ( .Y(n483), .A0(n468), .A1(n470) );
  inv01 U535 ( .Y(n473), .A(n483) );
  nor02 U536 ( .Y(n484), .A0(n474), .A1(n475) );
  inv01 U537 ( .Y(n477), .A(n484) );
  inv02 U538 ( .Y(B_not_41_), .A(B[41]) );
  inv02 U539 ( .Y(B_not_24_), .A(B[24]) );
  inv01 U540 ( .Y(DIFF[42]), .A(n485) );
  inv02 U541 ( .Y(carry_43_), .A(n486) );
  inv02 U542 ( .Y(n487), .A(B_not_42_) );
  inv02 U543 ( .Y(n488), .A(A[42]) );
  inv02 U544 ( .Y(n489), .A(carry_42_) );
  nor02 U545 ( .Y(n490), .A0(n487), .A1(n491) );
  nor02 U546 ( .Y(n492), .A0(n488), .A1(n493) );
  nor02 U547 ( .Y(n494), .A0(n489), .A1(n495) );
  nor02 U548 ( .Y(n496), .A0(n489), .A1(n497) );
  nor02 U549 ( .Y(n485), .A0(n498), .A1(n499) );
  nor02 U550 ( .Y(n500), .A0(n488), .A1(n489) );
  nor02 U551 ( .Y(n501), .A0(n487), .A1(n489) );
  nor02 U552 ( .Y(n502), .A0(n487), .A1(n488) );
  nor02 U553 ( .Y(n486), .A0(n502), .A1(n503) );
  nor02 U554 ( .Y(n504), .A0(A[42]), .A1(carry_42_) );
  inv01 U555 ( .Y(n491), .A(n504) );
  nor02 U556 ( .Y(n505), .A0(B_not_42_), .A1(carry_42_) );
  inv01 U557 ( .Y(n493), .A(n505) );
  nor02 U558 ( .Y(n506), .A0(B_not_42_), .A1(A[42]) );
  inv01 U559 ( .Y(n495), .A(n506) );
  nor02 U560 ( .Y(n507), .A0(n487), .A1(n488) );
  inv01 U561 ( .Y(n497), .A(n507) );
  nor02 U562 ( .Y(n508), .A0(n490), .A1(n492) );
  inv01 U563 ( .Y(n498), .A(n508) );
  nor02 U564 ( .Y(n509), .A0(n494), .A1(n496) );
  inv01 U565 ( .Y(n499), .A(n509) );
  nor02 U566 ( .Y(n510), .A0(n500), .A1(n501) );
  inv01 U567 ( .Y(n503), .A(n510) );
  inv01 U568 ( .Y(DIFF[50]), .A(n511) );
  inv02 U569 ( .Y(carry_51_), .A(n512) );
  inv02 U570 ( .Y(n513), .A(B_not_50_) );
  inv02 U571 ( .Y(n514), .A(A[50]) );
  inv02 U572 ( .Y(n515), .A(carry_50_) );
  nor02 U573 ( .Y(n516), .A0(n513), .A1(n517) );
  nor02 U574 ( .Y(n518), .A0(n514), .A1(n519) );
  nor02 U575 ( .Y(n520), .A0(n515), .A1(n521) );
  nor02 U576 ( .Y(n522), .A0(n515), .A1(n523) );
  nor02 U577 ( .Y(n511), .A0(n524), .A1(n525) );
  nor02 U578 ( .Y(n526), .A0(n514), .A1(n515) );
  nor02 U579 ( .Y(n527), .A0(n513), .A1(n515) );
  nor02 U580 ( .Y(n528), .A0(n513), .A1(n514) );
  nor02 U581 ( .Y(n512), .A0(n528), .A1(n529) );
  nor02 U582 ( .Y(n530), .A0(A[50]), .A1(carry_50_) );
  inv01 U583 ( .Y(n517), .A(n530) );
  nor02 U584 ( .Y(n531), .A0(B_not_50_), .A1(carry_50_) );
  inv01 U585 ( .Y(n519), .A(n531) );
  nor02 U586 ( .Y(n532), .A0(B_not_50_), .A1(A[50]) );
  inv01 U587 ( .Y(n521), .A(n532) );
  nor02 U588 ( .Y(n533), .A0(n513), .A1(n514) );
  inv01 U589 ( .Y(n523), .A(n533) );
  nor02 U590 ( .Y(n534), .A0(n516), .A1(n518) );
  inv01 U591 ( .Y(n524), .A(n534) );
  nor02 U592 ( .Y(n535), .A0(n520), .A1(n522) );
  inv01 U593 ( .Y(n525), .A(n535) );
  nor02 U594 ( .Y(n536), .A0(n526), .A1(n527) );
  inv01 U595 ( .Y(n529), .A(n536) );
  inv02 U596 ( .Y(B_not_42_), .A(B[42]) );
  inv02 U597 ( .Y(B_not_50_), .A(B[50]) );
  inv01 U598 ( .Y(DIFF[43]), .A(n537) );
  inv02 U599 ( .Y(carry_44_), .A(n538) );
  inv02 U600 ( .Y(n539), .A(B_not_43_) );
  inv02 U601 ( .Y(n540), .A(A[43]) );
  inv02 U602 ( .Y(n541), .A(carry_43_) );
  nor02 U603 ( .Y(n542), .A0(n539), .A1(n543) );
  nor02 U604 ( .Y(n544), .A0(n540), .A1(n545) );
  nor02 U605 ( .Y(n546), .A0(n541), .A1(n547) );
  nor02 U606 ( .Y(n548), .A0(n541), .A1(n549) );
  nor02 U607 ( .Y(n537), .A0(n550), .A1(n551) );
  nor02 U608 ( .Y(n552), .A0(n540), .A1(n541) );
  nor02 U609 ( .Y(n553), .A0(n539), .A1(n541) );
  nor02 U610 ( .Y(n554), .A0(n539), .A1(n540) );
  nor02 U611 ( .Y(n538), .A0(n554), .A1(n555) );
  nor02 U612 ( .Y(n556), .A0(A[43]), .A1(carry_43_) );
  inv01 U613 ( .Y(n543), .A(n556) );
  nor02 U614 ( .Y(n557), .A0(B_not_43_), .A1(carry_43_) );
  inv01 U615 ( .Y(n545), .A(n557) );
  nor02 U616 ( .Y(n558), .A0(B_not_43_), .A1(A[43]) );
  inv01 U617 ( .Y(n547), .A(n558) );
  nor02 U618 ( .Y(n559), .A0(n539), .A1(n540) );
  inv01 U619 ( .Y(n549), .A(n559) );
  nor02 U620 ( .Y(n560), .A0(n542), .A1(n544) );
  inv01 U621 ( .Y(n550), .A(n560) );
  nor02 U622 ( .Y(n561), .A0(n546), .A1(n548) );
  inv01 U623 ( .Y(n551), .A(n561) );
  nor02 U624 ( .Y(n562), .A0(n552), .A1(n553) );
  inv01 U625 ( .Y(n555), .A(n562) );
  inv01 U626 ( .Y(DIFF[49]), .A(n563) );
  inv02 U627 ( .Y(carry_50_), .A(n564) );
  inv02 U628 ( .Y(n565), .A(B_not_49_) );
  inv02 U629 ( .Y(n566), .A(A[49]) );
  inv02 U630 ( .Y(n567), .A(carry_49_) );
  nor02 U631 ( .Y(n568), .A0(n565), .A1(n569) );
  nor02 U632 ( .Y(n570), .A0(n566), .A1(n571) );
  nor02 U633 ( .Y(n572), .A0(n567), .A1(n573) );
  nor02 U634 ( .Y(n574), .A0(n567), .A1(n575) );
  nor02 U635 ( .Y(n563), .A0(n576), .A1(n577) );
  nor02 U636 ( .Y(n578), .A0(n566), .A1(n567) );
  nor02 U637 ( .Y(n579), .A0(n565), .A1(n567) );
  nor02 U638 ( .Y(n580), .A0(n565), .A1(n566) );
  nor02 U639 ( .Y(n564), .A0(n580), .A1(n581) );
  nor02 U640 ( .Y(n582), .A0(A[49]), .A1(carry_49_) );
  inv01 U641 ( .Y(n569), .A(n582) );
  nor02 U642 ( .Y(n583), .A0(B_not_49_), .A1(carry_49_) );
  inv01 U643 ( .Y(n571), .A(n583) );
  nor02 U644 ( .Y(n584), .A0(B_not_49_), .A1(A[49]) );
  inv01 U645 ( .Y(n573), .A(n584) );
  nor02 U646 ( .Y(n585), .A0(n565), .A1(n566) );
  inv01 U647 ( .Y(n575), .A(n585) );
  nor02 U648 ( .Y(n586), .A0(n568), .A1(n570) );
  inv01 U649 ( .Y(n576), .A(n586) );
  nor02 U650 ( .Y(n587), .A0(n572), .A1(n574) );
  inv01 U651 ( .Y(n577), .A(n587) );
  nor02 U652 ( .Y(n588), .A0(n578), .A1(n579) );
  inv01 U653 ( .Y(n581), .A(n588) );
  inv02 U654 ( .Y(B_not_43_), .A(B[43]) );
  inv02 U655 ( .Y(B_not_49_), .A(B[49]) );
  inv01 U656 ( .Y(DIFF[44]), .A(n589) );
  inv02 U657 ( .Y(carry_45_), .A(n590) );
  inv02 U658 ( .Y(n591), .A(B_not_44_) );
  inv02 U659 ( .Y(n592), .A(A[44]) );
  inv02 U660 ( .Y(n593), .A(carry_44_) );
  nor02 U661 ( .Y(n594), .A0(n591), .A1(n595) );
  nor02 U662 ( .Y(n596), .A0(n592), .A1(n597) );
  nor02 U663 ( .Y(n598), .A0(n593), .A1(n599) );
  nor02 U664 ( .Y(n600), .A0(n593), .A1(n601) );
  nor02 U665 ( .Y(n589), .A0(n602), .A1(n603) );
  nor02 U666 ( .Y(n604), .A0(n592), .A1(n593) );
  nor02 U667 ( .Y(n605), .A0(n591), .A1(n593) );
  nor02 U668 ( .Y(n606), .A0(n591), .A1(n592) );
  nor02 U669 ( .Y(n590), .A0(n606), .A1(n607) );
  nor02 U670 ( .Y(n608), .A0(A[44]), .A1(carry_44_) );
  inv01 U671 ( .Y(n595), .A(n608) );
  nor02 U672 ( .Y(n609), .A0(B_not_44_), .A1(carry_44_) );
  inv01 U673 ( .Y(n597), .A(n609) );
  nor02 U674 ( .Y(n610), .A0(B_not_44_), .A1(A[44]) );
  inv01 U675 ( .Y(n599), .A(n610) );
  nor02 U676 ( .Y(n611), .A0(n591), .A1(n592) );
  inv01 U677 ( .Y(n601), .A(n611) );
  nor02 U678 ( .Y(n612), .A0(n594), .A1(n596) );
  inv01 U679 ( .Y(n602), .A(n612) );
  nor02 U680 ( .Y(n613), .A0(n598), .A1(n600) );
  inv01 U681 ( .Y(n603), .A(n613) );
  nor02 U682 ( .Y(n614), .A0(n604), .A1(n605) );
  inv01 U683 ( .Y(n607), .A(n614) );
  inv01 U684 ( .Y(DIFF[48]), .A(n615) );
  inv02 U685 ( .Y(carry_49_), .A(n616) );
  inv02 U686 ( .Y(n617), .A(B_not_48_) );
  inv02 U687 ( .Y(n618), .A(A[48]) );
  inv02 U688 ( .Y(n619), .A(carry_48_) );
  nor02 U689 ( .Y(n620), .A0(n617), .A1(n621) );
  nor02 U690 ( .Y(n622), .A0(n618), .A1(n623) );
  nor02 U691 ( .Y(n624), .A0(n619), .A1(n625) );
  nor02 U692 ( .Y(n626), .A0(n619), .A1(n627) );
  nor02 U693 ( .Y(n615), .A0(n628), .A1(n629) );
  nor02 U694 ( .Y(n630), .A0(n618), .A1(n619) );
  nor02 U695 ( .Y(n631), .A0(n617), .A1(n619) );
  nor02 U696 ( .Y(n632), .A0(n617), .A1(n618) );
  nor02 U697 ( .Y(n616), .A0(n632), .A1(n633) );
  nor02 U698 ( .Y(n634), .A0(A[48]), .A1(carry_48_) );
  inv01 U699 ( .Y(n621), .A(n634) );
  nor02 U700 ( .Y(n635), .A0(B_not_48_), .A1(carry_48_) );
  inv01 U701 ( .Y(n623), .A(n635) );
  nor02 U702 ( .Y(n636), .A0(B_not_48_), .A1(A[48]) );
  inv01 U703 ( .Y(n625), .A(n636) );
  nor02 U704 ( .Y(n637), .A0(n617), .A1(n618) );
  inv01 U705 ( .Y(n627), .A(n637) );
  nor02 U706 ( .Y(n638), .A0(n620), .A1(n622) );
  inv01 U707 ( .Y(n628), .A(n638) );
  nor02 U708 ( .Y(n639), .A0(n624), .A1(n626) );
  inv01 U709 ( .Y(n629), .A(n639) );
  nor02 U710 ( .Y(n640), .A0(n630), .A1(n631) );
  inv01 U711 ( .Y(n633), .A(n640) );
  inv02 U712 ( .Y(B_not_44_), .A(B[44]) );
  inv02 U713 ( .Y(B_not_48_), .A(B[48]) );
  inv01 U714 ( .Y(DIFF[45]), .A(n641) );
  inv02 U715 ( .Y(carry_46_), .A(n642) );
  inv02 U716 ( .Y(n643), .A(B_not_45_) );
  inv02 U717 ( .Y(n644), .A(A[45]) );
  inv02 U718 ( .Y(n645), .A(carry_45_) );
  nor02 U719 ( .Y(n646), .A0(n643), .A1(n647) );
  nor02 U720 ( .Y(n648), .A0(n644), .A1(n649) );
  nor02 U721 ( .Y(n650), .A0(n645), .A1(n651) );
  nor02 U722 ( .Y(n652), .A0(n645), .A1(n653) );
  nor02 U723 ( .Y(n641), .A0(n654), .A1(n655) );
  nor02 U724 ( .Y(n656), .A0(n644), .A1(n645) );
  nor02 U725 ( .Y(n657), .A0(n643), .A1(n645) );
  nor02 U726 ( .Y(n658), .A0(n643), .A1(n644) );
  nor02 U727 ( .Y(n642), .A0(n658), .A1(n659) );
  nor02 U728 ( .Y(n660), .A0(A[45]), .A1(carry_45_) );
  inv01 U729 ( .Y(n647), .A(n660) );
  nor02 U730 ( .Y(n661), .A0(B_not_45_), .A1(carry_45_) );
  inv01 U731 ( .Y(n649), .A(n661) );
  nor02 U732 ( .Y(n662), .A0(B_not_45_), .A1(A[45]) );
  inv01 U733 ( .Y(n651), .A(n662) );
  nor02 U734 ( .Y(n663), .A0(n643), .A1(n644) );
  inv01 U735 ( .Y(n653), .A(n663) );
  nor02 U736 ( .Y(n664), .A0(n646), .A1(n648) );
  inv01 U737 ( .Y(n654), .A(n664) );
  nor02 U738 ( .Y(n665), .A0(n650), .A1(n652) );
  inv01 U739 ( .Y(n655), .A(n665) );
  nor02 U740 ( .Y(n666), .A0(n656), .A1(n657) );
  inv01 U741 ( .Y(n659), .A(n666) );
  inv01 U742 ( .Y(DIFF[47]), .A(n667) );
  inv02 U743 ( .Y(carry_48_), .A(n668) );
  inv02 U744 ( .Y(n669), .A(B_not_47_) );
  inv02 U745 ( .Y(n670), .A(A[47]) );
  inv02 U746 ( .Y(n671), .A(carry_47_) );
  nor02 U747 ( .Y(n672), .A0(n669), .A1(n673) );
  nor02 U748 ( .Y(n674), .A0(n670), .A1(n675) );
  nor02 U749 ( .Y(n676), .A0(n671), .A1(n677) );
  nor02 U750 ( .Y(n678), .A0(n671), .A1(n679) );
  nor02 U751 ( .Y(n667), .A0(n680), .A1(n681) );
  nor02 U752 ( .Y(n682), .A0(n670), .A1(n671) );
  nor02 U753 ( .Y(n683), .A0(n669), .A1(n671) );
  nor02 U754 ( .Y(n684), .A0(n669), .A1(n670) );
  nor02 U755 ( .Y(n668), .A0(n684), .A1(n685) );
  nor02 U756 ( .Y(n686), .A0(A[47]), .A1(carry_47_) );
  inv01 U757 ( .Y(n673), .A(n686) );
  nor02 U758 ( .Y(n687), .A0(B_not_47_), .A1(carry_47_) );
  inv01 U759 ( .Y(n675), .A(n687) );
  nor02 U760 ( .Y(n688), .A0(B_not_47_), .A1(A[47]) );
  inv01 U761 ( .Y(n677), .A(n688) );
  nor02 U762 ( .Y(n689), .A0(n669), .A1(n670) );
  inv01 U763 ( .Y(n679), .A(n689) );
  nor02 U764 ( .Y(n690), .A0(n672), .A1(n674) );
  inv01 U765 ( .Y(n680), .A(n690) );
  nor02 U766 ( .Y(n691), .A0(n676), .A1(n678) );
  inv01 U767 ( .Y(n681), .A(n691) );
  nor02 U768 ( .Y(n692), .A0(n682), .A1(n683) );
  inv01 U769 ( .Y(n685), .A(n692) );
  inv02 U770 ( .Y(B_not_45_), .A(B[45]) );
  inv02 U771 ( .Y(B_not_47_), .A(B[47]) );
  inv01 U772 ( .Y(DIFF[23]), .A(n693) );
  inv02 U773 ( .Y(carry_24_), .A(n694) );
  inv02 U774 ( .Y(n695), .A(B_not_23_) );
  inv02 U775 ( .Y(n696), .A(A[23]) );
  inv02 U776 ( .Y(n697), .A(carry_23_) );
  nor02 U777 ( .Y(n698), .A0(n695), .A1(n699) );
  nor02 U778 ( .Y(n700), .A0(n696), .A1(n701) );
  nor02 U779 ( .Y(n702), .A0(n697), .A1(n703) );
  nor02 U780 ( .Y(n704), .A0(n697), .A1(n705) );
  nor02 U781 ( .Y(n693), .A0(n706), .A1(n707) );
  nor02 U782 ( .Y(n708), .A0(n696), .A1(n697) );
  nor02 U783 ( .Y(n709), .A0(n695), .A1(n697) );
  nor02 U784 ( .Y(n710), .A0(n695), .A1(n696) );
  nor02 U785 ( .Y(n694), .A0(n710), .A1(n711) );
  nor02 U786 ( .Y(n712), .A0(A[23]), .A1(carry_23_) );
  inv01 U787 ( .Y(n699), .A(n712) );
  nor02 U788 ( .Y(n713), .A0(B_not_23_), .A1(carry_23_) );
  inv01 U789 ( .Y(n701), .A(n713) );
  nor02 U790 ( .Y(n714), .A0(B_not_23_), .A1(A[23]) );
  inv01 U791 ( .Y(n703), .A(n714) );
  nor02 U792 ( .Y(n715), .A0(n695), .A1(n696) );
  inv01 U793 ( .Y(n705), .A(n715) );
  nor02 U794 ( .Y(n716), .A0(n698), .A1(n700) );
  inv01 U795 ( .Y(n706), .A(n716) );
  nor02 U796 ( .Y(n717), .A0(n702), .A1(n704) );
  inv01 U797 ( .Y(n707), .A(n717) );
  nor02 U798 ( .Y(n718), .A0(n708), .A1(n709) );
  inv01 U799 ( .Y(n711), .A(n718) );
  inv01 U800 ( .Y(DIFF[46]), .A(n719) );
  inv02 U801 ( .Y(carry_47_), .A(n720) );
  inv02 U802 ( .Y(n721), .A(B_not_46_) );
  inv02 U803 ( .Y(n722), .A(A[46]) );
  inv02 U804 ( .Y(n723), .A(carry_46_) );
  nor02 U805 ( .Y(n724), .A0(n721), .A1(n725) );
  nor02 U806 ( .Y(n726), .A0(n722), .A1(n727) );
  nor02 U807 ( .Y(n728), .A0(n723), .A1(n729) );
  nor02 U808 ( .Y(n730), .A0(n723), .A1(n731) );
  nor02 U809 ( .Y(n719), .A0(n732), .A1(n733) );
  nor02 U810 ( .Y(n734), .A0(n722), .A1(n723) );
  nor02 U811 ( .Y(n735), .A0(n721), .A1(n723) );
  nor02 U812 ( .Y(n736), .A0(n721), .A1(n722) );
  nor02 U813 ( .Y(n720), .A0(n736), .A1(n737) );
  nor02 U814 ( .Y(n738), .A0(A[46]), .A1(carry_46_) );
  inv01 U815 ( .Y(n725), .A(n738) );
  nor02 U816 ( .Y(n739), .A0(B_not_46_), .A1(carry_46_) );
  inv01 U817 ( .Y(n727), .A(n739) );
  nor02 U818 ( .Y(n740), .A0(B_not_46_), .A1(A[46]) );
  inv01 U819 ( .Y(n729), .A(n740) );
  nor02 U820 ( .Y(n741), .A0(n721), .A1(n722) );
  inv01 U821 ( .Y(n731), .A(n741) );
  nor02 U822 ( .Y(n742), .A0(n724), .A1(n726) );
  inv01 U823 ( .Y(n732), .A(n742) );
  nor02 U824 ( .Y(n743), .A0(n728), .A1(n730) );
  inv01 U825 ( .Y(n733), .A(n743) );
  nor02 U826 ( .Y(n744), .A0(n734), .A1(n735) );
  inv01 U827 ( .Y(n737), .A(n744) );
  inv02 U828 ( .Y(B_not_23_), .A(B[23]) );
  inv02 U829 ( .Y(B_not_46_), .A(B[46]) );
  inv01 U830 ( .Y(DIFF[22]), .A(n745) );
  inv02 U831 ( .Y(carry_23_), .A(n746) );
  inv02 U832 ( .Y(n747), .A(B_not_22_) );
  inv02 U833 ( .Y(n748), .A(A[22]) );
  inv02 U834 ( .Y(n749), .A(carry_22_) );
  nor02 U835 ( .Y(n750), .A0(n747), .A1(n751) );
  nor02 U836 ( .Y(n752), .A0(n748), .A1(n753) );
  nor02 U837 ( .Y(n754), .A0(n749), .A1(n755) );
  nor02 U838 ( .Y(n756), .A0(n749), .A1(n757) );
  nor02 U839 ( .Y(n745), .A0(n758), .A1(n759) );
  nor02 U840 ( .Y(n760), .A0(n748), .A1(n749) );
  nor02 U841 ( .Y(n761), .A0(n747), .A1(n749) );
  nor02 U842 ( .Y(n762), .A0(n747), .A1(n748) );
  nor02 U843 ( .Y(n746), .A0(n762), .A1(n763) );
  nor02 U844 ( .Y(n764), .A0(A[22]), .A1(carry_22_) );
  inv01 U845 ( .Y(n751), .A(n764) );
  nor02 U846 ( .Y(n765), .A0(B_not_22_), .A1(carry_22_) );
  inv01 U847 ( .Y(n753), .A(n765) );
  nor02 U848 ( .Y(n766), .A0(B_not_22_), .A1(A[22]) );
  inv01 U849 ( .Y(n755), .A(n766) );
  nor02 U850 ( .Y(n767), .A0(n747), .A1(n748) );
  inv01 U851 ( .Y(n757), .A(n767) );
  nor02 U852 ( .Y(n768), .A0(n750), .A1(n752) );
  inv01 U853 ( .Y(n758), .A(n768) );
  nor02 U854 ( .Y(n769), .A0(n754), .A1(n756) );
  inv01 U855 ( .Y(n759), .A(n769) );
  nor02 U856 ( .Y(n770), .A0(n760), .A1(n761) );
  inv01 U857 ( .Y(n763), .A(n770) );
  inv02 U858 ( .Y(B_not_22_), .A(B[22]) );
  inv01 U859 ( .Y(DIFF[21]), .A(n771) );
  inv02 U860 ( .Y(carry_22_), .A(n772) );
  inv02 U861 ( .Y(n773), .A(B_not_21_) );
  inv02 U862 ( .Y(n774), .A(A[21]) );
  inv02 U863 ( .Y(n775), .A(n797) );
  nor02 U864 ( .Y(n776), .A0(n773), .A1(n777) );
  nor02 U865 ( .Y(n778), .A0(n774), .A1(n779) );
  nor02 U866 ( .Y(n780), .A0(n775), .A1(n781) );
  nor02 U867 ( .Y(n782), .A0(n775), .A1(n783) );
  nor02 U868 ( .Y(n771), .A0(n784), .A1(n785) );
  nor02 U869 ( .Y(n786), .A0(n774), .A1(n775) );
  nor02 U870 ( .Y(n787), .A0(n773), .A1(n775) );
  nor02 U871 ( .Y(n788), .A0(n773), .A1(n774) );
  nor02 U872 ( .Y(n772), .A0(n788), .A1(n789) );
  nor02 U873 ( .Y(n790), .A0(A[21]), .A1(n797) );
  inv01 U874 ( .Y(n777), .A(n790) );
  nor02 U875 ( .Y(n791), .A0(B_not_21_), .A1(n797) );
  inv01 U876 ( .Y(n779), .A(n791) );
  nor02 U877 ( .Y(n792), .A0(B_not_21_), .A1(A[21]) );
  inv01 U878 ( .Y(n781), .A(n792) );
  nor02 U879 ( .Y(n793), .A0(n773), .A1(n774) );
  inv01 U880 ( .Y(n783), .A(n793) );
  nor02 U881 ( .Y(n794), .A0(n776), .A1(n778) );
  inv01 U882 ( .Y(n784), .A(n794) );
  nor02 U883 ( .Y(n795), .A0(n780), .A1(n782) );
  inv01 U884 ( .Y(n785), .A(n795) );
  nor02 U885 ( .Y(n796), .A0(n786), .A1(n787) );
  inv01 U886 ( .Y(n789), .A(n796) );
  inv02 U887 ( .Y(B_not_21_), .A(B[21]) );
  buf02 U888 ( .Y(n797), .A(carry_21_) );
  buf02 U889 ( .Y(n798), .A(carry_20_) );
  inv01 U890 ( .Y(DIFF[18]), .A(n799) );
  inv02 U891 ( .Y(carry_19_), .A(n800) );
  inv02 U892 ( .Y(n801), .A(B_not_18_) );
  inv02 U893 ( .Y(n802), .A(A[18]) );
  inv02 U894 ( .Y(n803), .A(carry_18_) );
  nor02 U895 ( .Y(n804), .A0(n801), .A1(n805) );
  nor02 U896 ( .Y(n806), .A0(n802), .A1(n807) );
  nor02 U897 ( .Y(n808), .A0(n803), .A1(n809) );
  nor02 U898 ( .Y(n810), .A0(n803), .A1(n811) );
  nor02 U899 ( .Y(n799), .A0(n812), .A1(n813) );
  nor02 U900 ( .Y(n814), .A0(n802), .A1(n803) );
  nor02 U901 ( .Y(n815), .A0(n801), .A1(n803) );
  nor02 U902 ( .Y(n816), .A0(n801), .A1(n802) );
  nor02 U903 ( .Y(n800), .A0(n816), .A1(n817) );
  nor02 U904 ( .Y(n818), .A0(A[18]), .A1(carry_18_) );
  inv01 U905 ( .Y(n805), .A(n818) );
  nor02 U906 ( .Y(n819), .A0(B_not_18_), .A1(carry_18_) );
  inv01 U907 ( .Y(n807), .A(n819) );
  nor02 U908 ( .Y(n820), .A0(B_not_18_), .A1(A[18]) );
  inv01 U909 ( .Y(n809), .A(n820) );
  nor02 U910 ( .Y(n821), .A0(n801), .A1(n802) );
  inv01 U911 ( .Y(n811), .A(n821) );
  nor02 U912 ( .Y(n822), .A0(n804), .A1(n806) );
  inv01 U913 ( .Y(n812), .A(n822) );
  nor02 U914 ( .Y(n823), .A0(n808), .A1(n810) );
  inv01 U915 ( .Y(n813), .A(n823) );
  nor02 U916 ( .Y(n824), .A0(n814), .A1(n815) );
  inv01 U917 ( .Y(n817), .A(n824) );
  inv02 U918 ( .Y(B_not_18_), .A(B[18]) );
  inv01 U919 ( .Y(DIFF[17]), .A(n825) );
  inv02 U920 ( .Y(carry_18_), .A(n826) );
  inv02 U921 ( .Y(n827), .A(B_not_17_) );
  inv02 U922 ( .Y(n828), .A(A[17]) );
  inv02 U923 ( .Y(n829), .A(carry_17_) );
  nor02 U924 ( .Y(n830), .A0(n827), .A1(n831) );
  nor02 U925 ( .Y(n832), .A0(n828), .A1(n833) );
  nor02 U926 ( .Y(n834), .A0(n829), .A1(n835) );
  nor02 U927 ( .Y(n836), .A0(n829), .A1(n837) );
  nor02 U928 ( .Y(n825), .A0(n838), .A1(n839) );
  nor02 U929 ( .Y(n840), .A0(n828), .A1(n829) );
  nor02 U930 ( .Y(n841), .A0(n827), .A1(n829) );
  nor02 U931 ( .Y(n842), .A0(n827), .A1(n828) );
  nor02 U932 ( .Y(n826), .A0(n842), .A1(n843) );
  nor02 U933 ( .Y(n844), .A0(A[17]), .A1(carry_17_) );
  inv01 U934 ( .Y(n831), .A(n844) );
  nor02 U935 ( .Y(n845), .A0(B_not_17_), .A1(carry_17_) );
  inv01 U936 ( .Y(n833), .A(n845) );
  nor02 U937 ( .Y(n846), .A0(B_not_17_), .A1(A[17]) );
  inv01 U938 ( .Y(n835), .A(n846) );
  nor02 U939 ( .Y(n847), .A0(n827), .A1(n828) );
  inv01 U940 ( .Y(n837), .A(n847) );
  nor02 U941 ( .Y(n848), .A0(n830), .A1(n832) );
  inv01 U942 ( .Y(n838), .A(n848) );
  nor02 U943 ( .Y(n849), .A0(n834), .A1(n836) );
  inv01 U944 ( .Y(n839), .A(n849) );
  nor02 U945 ( .Y(n850), .A0(n840), .A1(n841) );
  inv01 U946 ( .Y(n843), .A(n850) );
  inv02 U947 ( .Y(B_not_17_), .A(B[17]) );
  inv01 U948 ( .Y(DIFF[16]), .A(n851) );
  inv02 U949 ( .Y(carry_17_), .A(n852) );
  inv02 U950 ( .Y(n853), .A(B_not_16_) );
  inv02 U951 ( .Y(n854), .A(A[16]) );
  inv02 U952 ( .Y(n855), .A(n877) );
  nor02 U953 ( .Y(n856), .A0(n853), .A1(n857) );
  nor02 U954 ( .Y(n858), .A0(n854), .A1(n859) );
  nor02 U955 ( .Y(n860), .A0(n855), .A1(n861) );
  nor02 U956 ( .Y(n862), .A0(n855), .A1(n863) );
  nor02 U957 ( .Y(n851), .A0(n864), .A1(n865) );
  nor02 U958 ( .Y(n866), .A0(n854), .A1(n855) );
  nor02 U959 ( .Y(n867), .A0(n853), .A1(n855) );
  nor02 U960 ( .Y(n868), .A0(n853), .A1(n854) );
  nor02 U961 ( .Y(n852), .A0(n868), .A1(n869) );
  nor02 U962 ( .Y(n870), .A0(A[16]), .A1(n877) );
  inv01 U963 ( .Y(n857), .A(n870) );
  nor02 U964 ( .Y(n871), .A0(B_not_16_), .A1(n877) );
  inv01 U965 ( .Y(n859), .A(n871) );
  nor02 U966 ( .Y(n872), .A0(B_not_16_), .A1(A[16]) );
  inv01 U967 ( .Y(n861), .A(n872) );
  nor02 U968 ( .Y(n873), .A0(n853), .A1(n854) );
  inv01 U969 ( .Y(n863), .A(n873) );
  nor02 U970 ( .Y(n874), .A0(n856), .A1(n858) );
  inv01 U971 ( .Y(n864), .A(n874) );
  nor02 U972 ( .Y(n875), .A0(n860), .A1(n862) );
  inv01 U973 ( .Y(n865), .A(n875) );
  nor02 U974 ( .Y(n876), .A0(n866), .A1(n867) );
  inv01 U975 ( .Y(n869), .A(n876) );
  inv02 U976 ( .Y(B_not_16_), .A(B[16]) );
  buf02 U977 ( .Y(n877), .A(carry_16_) );
  buf02 U978 ( .Y(n878), .A(carry_15_) );
  buf02 U979 ( .Y(n879), .A(carry_14_) );
  inv01 U980 ( .Y(DIFF[12]), .A(n880) );
  inv02 U981 ( .Y(carry_13_), .A(n881) );
  inv02 U982 ( .Y(n882), .A(B_not_12_) );
  inv02 U983 ( .Y(n883), .A(A[12]) );
  inv02 U984 ( .Y(n884), .A(carry_12_) );
  nor02 U985 ( .Y(n885), .A0(n882), .A1(n886) );
  nor02 U986 ( .Y(n887), .A0(n883), .A1(n888) );
  nor02 U987 ( .Y(n889), .A0(n884), .A1(n890) );
  nor02 U988 ( .Y(n891), .A0(n884), .A1(n892) );
  nor02 U989 ( .Y(n880), .A0(n893), .A1(n894) );
  nor02 U990 ( .Y(n895), .A0(n883), .A1(n884) );
  nor02 U991 ( .Y(n896), .A0(n882), .A1(n884) );
  nor02 U992 ( .Y(n897), .A0(n882), .A1(n883) );
  nor02 U993 ( .Y(n881), .A0(n897), .A1(n898) );
  nor02 U994 ( .Y(n899), .A0(A[12]), .A1(carry_12_) );
  inv01 U995 ( .Y(n886), .A(n899) );
  nor02 U996 ( .Y(n900), .A0(B_not_12_), .A1(carry_12_) );
  inv01 U997 ( .Y(n888), .A(n900) );
  nor02 U998 ( .Y(n901), .A0(B_not_12_), .A1(A[12]) );
  inv01 U999 ( .Y(n890), .A(n901) );
  nor02 U1000 ( .Y(n902), .A0(n882), .A1(n883) );
  inv01 U1001 ( .Y(n892), .A(n902) );
  nor02 U1002 ( .Y(n903), .A0(n885), .A1(n887) );
  inv01 U1003 ( .Y(n893), .A(n903) );
  nor02 U1004 ( .Y(n904), .A0(n889), .A1(n891) );
  inv01 U1005 ( .Y(n894), .A(n904) );
  nor02 U1006 ( .Y(n905), .A0(n895), .A1(n896) );
  inv01 U1007 ( .Y(n898), .A(n905) );
  inv02 U1008 ( .Y(B_not_12_), .A(B[12]) );
  inv01 U1009 ( .Y(DIFF[11]), .A(n906) );
  inv02 U1010 ( .Y(carry_12_), .A(n907) );
  inv02 U1011 ( .Y(n908), .A(B_not_11_) );
  inv02 U1012 ( .Y(n909), .A(A[11]) );
  inv02 U1013 ( .Y(n910), .A(carry_11_) );
  nor02 U1014 ( .Y(n911), .A0(n908), .A1(n912) );
  nor02 U1015 ( .Y(n913), .A0(n909), .A1(n914) );
  nor02 U1016 ( .Y(n915), .A0(n910), .A1(n916) );
  nor02 U1017 ( .Y(n917), .A0(n910), .A1(n918) );
  nor02 U1018 ( .Y(n906), .A0(n919), .A1(n920) );
  nor02 U1019 ( .Y(n921), .A0(n909), .A1(n910) );
  nor02 U1020 ( .Y(n922), .A0(n908), .A1(n910) );
  nor02 U1021 ( .Y(n923), .A0(n908), .A1(n909) );
  nor02 U1022 ( .Y(n907), .A0(n923), .A1(n924) );
  nor02 U1023 ( .Y(n925), .A0(A[11]), .A1(carry_11_) );
  inv01 U1024 ( .Y(n912), .A(n925) );
  nor02 U1025 ( .Y(n926), .A0(B_not_11_), .A1(carry_11_) );
  inv01 U1026 ( .Y(n914), .A(n926) );
  nor02 U1027 ( .Y(n927), .A0(B_not_11_), .A1(A[11]) );
  inv01 U1028 ( .Y(n916), .A(n927) );
  nor02 U1029 ( .Y(n928), .A0(n908), .A1(n909) );
  inv01 U1030 ( .Y(n918), .A(n928) );
  nor02 U1031 ( .Y(n929), .A0(n911), .A1(n913) );
  inv01 U1032 ( .Y(n919), .A(n929) );
  nor02 U1033 ( .Y(n930), .A0(n915), .A1(n917) );
  inv01 U1034 ( .Y(n920), .A(n930) );
  nor02 U1035 ( .Y(n931), .A0(n921), .A1(n922) );
  inv01 U1036 ( .Y(n924), .A(n931) );
  inv02 U1037 ( .Y(B_not_11_), .A(B[11]) );
  inv01 U1038 ( .Y(DIFF[10]), .A(n932) );
  inv02 U1039 ( .Y(carry_11_), .A(n933) );
  inv02 U1040 ( .Y(n934), .A(B_not_10_) );
  inv02 U1041 ( .Y(n935), .A(A[10]) );
  inv02 U1042 ( .Y(n936), .A(n958) );
  nor02 U1043 ( .Y(n937), .A0(n934), .A1(n938) );
  nor02 U1044 ( .Y(n939), .A0(n935), .A1(n940) );
  nor02 U1045 ( .Y(n941), .A0(n936), .A1(n942) );
  nor02 U1046 ( .Y(n943), .A0(n936), .A1(n944) );
  nor02 U1047 ( .Y(n932), .A0(n945), .A1(n946) );
  nor02 U1048 ( .Y(n947), .A0(n935), .A1(n936) );
  nor02 U1049 ( .Y(n948), .A0(n934), .A1(n936) );
  nor02 U1050 ( .Y(n949), .A0(n934), .A1(n935) );
  nor02 U1051 ( .Y(n933), .A0(n949), .A1(n950) );
  nor02 U1052 ( .Y(n951), .A0(A[10]), .A1(n958) );
  inv01 U1053 ( .Y(n938), .A(n951) );
  nor02 U1054 ( .Y(n952), .A0(B_not_10_), .A1(n958) );
  inv01 U1055 ( .Y(n940), .A(n952) );
  nor02 U1056 ( .Y(n953), .A0(B_not_10_), .A1(A[10]) );
  inv01 U1057 ( .Y(n942), .A(n953) );
  nor02 U1058 ( .Y(n954), .A0(n934), .A1(n935) );
  inv01 U1059 ( .Y(n944), .A(n954) );
  nor02 U1060 ( .Y(n955), .A0(n937), .A1(n939) );
  inv01 U1061 ( .Y(n945), .A(n955) );
  nor02 U1062 ( .Y(n956), .A0(n941), .A1(n943) );
  inv01 U1063 ( .Y(n946), .A(n956) );
  nor02 U1064 ( .Y(n957), .A0(n947), .A1(n948) );
  inv01 U1065 ( .Y(n950), .A(n957) );
  inv02 U1066 ( .Y(B_not_10_), .A(B[10]) );
  buf02 U1067 ( .Y(n958), .A(carry_10_) );
  buf02 U1068 ( .Y(n959), .A(carry_9_) );
  buf02 U1069 ( .Y(n960), .A(carry_8_) );
  inv01 U1070 ( .Y(DIFF[6]), .A(n961) );
  inv02 U1071 ( .Y(carry_7_), .A(n962) );
  inv02 U1072 ( .Y(n963), .A(B_not_6_) );
  inv02 U1073 ( .Y(n964), .A(A[6]) );
  inv02 U1074 ( .Y(n965), .A(carry_6_) );
  nor02 U1075 ( .Y(n966), .A0(n963), .A1(n967) );
  nor02 U1076 ( .Y(n968), .A0(n964), .A1(n969) );
  nor02 U1077 ( .Y(n970), .A0(n965), .A1(n971) );
  nor02 U1078 ( .Y(n972), .A0(n965), .A1(n973) );
  nor02 U1079 ( .Y(n961), .A0(n974), .A1(n975) );
  nor02 U1080 ( .Y(n976), .A0(n964), .A1(n965) );
  nor02 U1081 ( .Y(n977), .A0(n963), .A1(n965) );
  nor02 U1082 ( .Y(n978), .A0(n963), .A1(n964) );
  nor02 U1083 ( .Y(n962), .A0(n978), .A1(n979) );
  nor02 U1084 ( .Y(n980), .A0(A[6]), .A1(carry_6_) );
  inv01 U1085 ( .Y(n967), .A(n980) );
  nor02 U1086 ( .Y(n981), .A0(B_not_6_), .A1(carry_6_) );
  inv01 U1087 ( .Y(n969), .A(n981) );
  nor02 U1088 ( .Y(n982), .A0(B_not_6_), .A1(A[6]) );
  inv01 U1089 ( .Y(n971), .A(n982) );
  nor02 U1090 ( .Y(n983), .A0(n963), .A1(n964) );
  inv01 U1091 ( .Y(n973), .A(n983) );
  nor02 U1092 ( .Y(n984), .A0(n966), .A1(n968) );
  inv01 U1093 ( .Y(n974), .A(n984) );
  nor02 U1094 ( .Y(n985), .A0(n970), .A1(n972) );
  inv01 U1095 ( .Y(n975), .A(n985) );
  nor02 U1096 ( .Y(n986), .A0(n976), .A1(n977) );
  inv01 U1097 ( .Y(n979), .A(n986) );
  inv02 U1098 ( .Y(B_not_6_), .A(B[6]) );
  inv01 U1099 ( .Y(DIFF[5]), .A(n987) );
  inv02 U1100 ( .Y(carry_6_), .A(n988) );
  inv02 U1101 ( .Y(n989), .A(B_not_5_) );
  inv02 U1102 ( .Y(n990), .A(A[5]) );
  inv02 U1103 ( .Y(n991), .A(n1013) );
  nor02 U1104 ( .Y(n992), .A0(n989), .A1(n993) );
  nor02 U1105 ( .Y(n994), .A0(n990), .A1(n995) );
  nor02 U1106 ( .Y(n996), .A0(n991), .A1(n997) );
  nor02 U1107 ( .Y(n998), .A0(n991), .A1(n999) );
  nor02 U1108 ( .Y(n987), .A0(n1000), .A1(n1001) );
  nor02 U1109 ( .Y(n1002), .A0(n990), .A1(n991) );
  nor02 U1110 ( .Y(n1003), .A0(n989), .A1(n991) );
  nor02 U1111 ( .Y(n1004), .A0(n989), .A1(n990) );
  nor02 U1112 ( .Y(n988), .A0(n1004), .A1(n1005) );
  nor02 U1113 ( .Y(n1006), .A0(A[5]), .A1(n1013) );
  inv01 U1114 ( .Y(n993), .A(n1006) );
  nor02 U1115 ( .Y(n1007), .A0(B_not_5_), .A1(n1013) );
  inv01 U1116 ( .Y(n995), .A(n1007) );
  nor02 U1117 ( .Y(n1008), .A0(B_not_5_), .A1(A[5]) );
  inv01 U1118 ( .Y(n997), .A(n1008) );
  nor02 U1119 ( .Y(n1009), .A0(n989), .A1(n990) );
  inv01 U1120 ( .Y(n999), .A(n1009) );
  nor02 U1121 ( .Y(n1010), .A0(n992), .A1(n994) );
  inv01 U1122 ( .Y(n1000), .A(n1010) );
  nor02 U1123 ( .Y(n1011), .A0(n996), .A1(n998) );
  inv01 U1124 ( .Y(n1001), .A(n1011) );
  nor02 U1125 ( .Y(n1012), .A0(n1002), .A1(n1003) );
  inv01 U1126 ( .Y(n1005), .A(n1012) );
  inv02 U1127 ( .Y(B_not_5_), .A(B[5]) );
  buf02 U1128 ( .Y(n1013), .A(carry_5_) );
  inv01 U1129 ( .Y(DIFF[3]), .A(n1014) );
  inv02 U1130 ( .Y(carry_4_), .A(n1015) );
  inv02 U1131 ( .Y(n1016), .A(B_not_3_) );
  inv02 U1132 ( .Y(n1017), .A(A[3]) );
  inv02 U1133 ( .Y(n1018), .A(carry_3_) );
  nor02 U1134 ( .Y(n1019), .A0(n1016), .A1(n1020) );
  nor02 U1135 ( .Y(n1021), .A0(n1017), .A1(n1022) );
  nor02 U1136 ( .Y(n1023), .A0(n1018), .A1(n1024) );
  nor02 U1137 ( .Y(n1025), .A0(n1018), .A1(n1026) );
  nor02 U1138 ( .Y(n1014), .A0(n1027), .A1(n1028) );
  nor02 U1139 ( .Y(n1029), .A0(n1017), .A1(n1018) );
  nor02 U1140 ( .Y(n1030), .A0(n1016), .A1(n1018) );
  nor02 U1141 ( .Y(n1031), .A0(n1016), .A1(n1017) );
  nor02 U1142 ( .Y(n1015), .A0(n1031), .A1(n1032) );
  nor02 U1143 ( .Y(n1033), .A0(A[3]), .A1(carry_3_) );
  inv01 U1144 ( .Y(n1020), .A(n1033) );
  nor02 U1145 ( .Y(n1034), .A0(B_not_3_), .A1(carry_3_) );
  inv01 U1146 ( .Y(n1022), .A(n1034) );
  nor02 U1147 ( .Y(n1035), .A0(B_not_3_), .A1(A[3]) );
  inv01 U1148 ( .Y(n1024), .A(n1035) );
  nor02 U1149 ( .Y(n1036), .A0(n1016), .A1(n1017) );
  inv01 U1150 ( .Y(n1026), .A(n1036) );
  nor02 U1151 ( .Y(n1037), .A0(n1019), .A1(n1021) );
  inv01 U1152 ( .Y(n1027), .A(n1037) );
  nor02 U1153 ( .Y(n1038), .A0(n1023), .A1(n1025) );
  inv01 U1154 ( .Y(n1028), .A(n1038) );
  nor02 U1155 ( .Y(n1039), .A0(n1029), .A1(n1030) );
  inv01 U1156 ( .Y(n1032), .A(n1039) );
  inv02 U1157 ( .Y(B_not_3_), .A(B[3]) );
  inv01 U1158 ( .Y(n1040), .A(n1045) );
  inv01 U1159 ( .Y(DIFF[2]), .A(n1041) );
  inv02 U1160 ( .Y(carry_3_), .A(n1042) );
  inv02 U1161 ( .Y(n1043), .A(B_not_2_) );
  inv02 U1162 ( .Y(n1044), .A(A[2]) );
  inv02 U1163 ( .Y(n1045), .A(carry_2_) );
  nor02 U1164 ( .Y(n1046), .A0(n1043), .A1(n1047) );
  nor02 U1165 ( .Y(n1048), .A0(n1044), .A1(n1049) );
  nor02 U1166 ( .Y(n1050), .A0(n1045), .A1(n1051) );
  nor02 U1167 ( .Y(n1052), .A0(n1045), .A1(n1053) );
  nor02 U1168 ( .Y(n1041), .A0(n1054), .A1(n1055) );
  nor02 U1169 ( .Y(n1056), .A0(n1044), .A1(n1045) );
  nor02 U1170 ( .Y(n1057), .A0(n1043), .A1(n1045) );
  nor02 U1171 ( .Y(n1058), .A0(n1043), .A1(n1044) );
  nor02 U1172 ( .Y(n1042), .A0(n1058), .A1(n1059) );
  nor02 U1173 ( .Y(n1060), .A0(A[2]), .A1(carry_2_) );
  inv01 U1174 ( .Y(n1047), .A(n1060) );
  nor02 U1175 ( .Y(n1061), .A0(B_not_2_), .A1(n1040) );
  inv01 U1176 ( .Y(n1049), .A(n1061) );
  nor02 U1177 ( .Y(n1062), .A0(B_not_2_), .A1(A[2]) );
  inv01 U1178 ( .Y(n1051), .A(n1062) );
  nor02 U1179 ( .Y(n1063), .A0(n1043), .A1(n1044) );
  inv01 U1180 ( .Y(n1053), .A(n1063) );
  nor02 U1181 ( .Y(n1064), .A0(n1046), .A1(n1048) );
  inv01 U1182 ( .Y(n1054), .A(n1064) );
  nor02 U1183 ( .Y(n1065), .A0(n1050), .A1(n1052) );
  inv01 U1184 ( .Y(n1055), .A(n1065) );
  nor02 U1185 ( .Y(n1066), .A0(n1056), .A1(n1057) );
  inv01 U1186 ( .Y(n1059), .A(n1066) );
  inv02 U1187 ( .Y(B_not_2_), .A(B[2]) );
  or02 U1188 ( .Y(carry_2_), .A0(B_not_1_), .A1(A[1]) );
  inv04 U1189 ( .Y(B_not_9_), .A(B[9]) );
  inv04 U1190 ( .Y(B_not_8_), .A(B[8]) );
  inv04 U1191 ( .Y(B_not_7_), .A(B[7]) );
  inv04 U1192 ( .Y(B_not_51_), .A(B[51]) );
  inv04 U1193 ( .Y(B_not_4_), .A(B[4]) );
  inv04 U1194 ( .Y(B_not_20_), .A(B[20]) );
  inv04 U1195 ( .Y(B_not_1_), .A(B[1]) );
  inv04 U1196 ( .Y(B_not_19_), .A(B[19]) );
  inv04 U1197 ( .Y(B_not_15_), .A(B[15]) );
  inv04 U1198 ( .Y(B_not_14_), .A(B[14]) );
  inv04 U1199 ( .Y(B_not_13_), .A(B[13]) );
  fadd1 U2_4 ( .S(n1076), .CO(carry_5_), .A(A[4]), .B(B_not_4_), .CI(carry_4_)
         );
  fadd1 U2_7 ( .S(n1075), .CO(carry_8_), .A(A[7]), .B(B_not_7_), .CI(carry_7_)
         );
  fadd1 U2_8 ( .S(n1074), .CO(carry_9_), .A(A[8]), .B(B_not_8_), .CI(n960) );
  fadd1 U2_9 ( .S(n1073), .CO(carry_10_), .A(A[9]), .B(B_not_9_), .CI(n959) );
  fadd1 U2_13 ( .S(n1072), .CO(carry_14_), .A(A[13]), .B(B_not_13_), .CI(
        carry_13_) );
  fadd1 U2_14 ( .S(n1071), .CO(carry_15_), .A(A[14]), .B(B_not_14_), .CI(n879)
         );
  fadd1 U2_15 ( .S(n1070), .CO(carry_16_), .A(A[15]), .B(B_not_15_), .CI(n878)
         );
  fadd1 U2_19 ( .S(n1069), .CO(carry_20_), .A(A[19]), .B(B_not_19_), .CI(
        carry_19_) );
  fadd1 U2_20 ( .S(n1068), .CO(carry_21_), .A(A[20]), .B(B_not_20_), .CI(n798)
         );
  fadd1 U2_51 ( .S(n1067), .A(A[51]), .B(B_not_51_), .CI(carry_51_) );
endmodule


module sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_dec_26_0 ( A, SUM );
  input [25:0] A;
  output [25:0] SUM;
  wire   carry_25_, carry_23_, carry_22_, carry_20_, carry_19_, carry_17_,
         carry_16_, carry_15_, carry_14_, carry_13_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, carry_6_, carry_5_, carry_4_, carry_3_,
         carry_2_, n5, n7, n9, n11, n13, n15, n17, n19, n21, n23, n25, n27,
         n29, n31, n33, n35, n37, n39, n41, n43, n45, n47, n49, n51, n53, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  xor2 U6 ( .Y(n5), .A0(carry_25_), .A1(A[25]) );
  inv01 U7 ( .Y(SUM[25]), .A(n5) );
  xor2 U8 ( .Y(n7), .A0(A[1]), .A1(A[0]) );
  inv01 U9 ( .Y(SUM[1]), .A(n7) );
  xor2 U10 ( .Y(n9), .A0(A[22]), .A1(n65) );
  inv01 U11 ( .Y(SUM[22]), .A(n9) );
  xor2 U12 ( .Y(n11), .A0(A[4]), .A1(n71) );
  inv01 U13 ( .Y(SUM[4]), .A(n11) );
  xor2 U14 ( .Y(n13), .A0(A[24]), .A1(n64) );
  inv01 U15 ( .Y(SUM[24]), .A(n13) );
  xor2 U16 ( .Y(n15), .A0(A[10]), .A1(n77) );
  inv01 U17 ( .Y(SUM[10]), .A(n15) );
  xor2 U18 ( .Y(n17), .A0(A[15]), .A1(n75) );
  inv01 U19 ( .Y(SUM[15]), .A(n17) );
  xor2 U20 ( .Y(n19), .A0(A[16]), .A1(n73) );
  inv01 U21 ( .Y(SUM[16]), .A(n19) );
  xor2 U22 ( .Y(n21), .A0(A[9]), .A1(n74) );
  inv01 U23 ( .Y(SUM[9]), .A(n21) );
  xor2 U24 ( .Y(n23), .A0(A[5]), .A1(n76) );
  inv01 U25 ( .Y(SUM[5]), .A(n23) );
  xor2 U26 ( .Y(n25), .A0(A[2]), .A1(n55) );
  inv01 U27 ( .Y(SUM[2]), .A(n25) );
  xor2 U28 ( .Y(n27), .A0(A[21]), .A1(n59) );
  inv01 U29 ( .Y(SUM[21]), .A(n27) );
  xor2 U30 ( .Y(n29), .A0(A[17]), .A1(n78) );
  inv01 U31 ( .Y(SUM[17]), .A(n29) );
  xor2 U32 ( .Y(n31), .A0(A[20]), .A1(n80) );
  inv01 U33 ( .Y(SUM[20]), .A(n31) );
  xor2 U34 ( .Y(n33), .A0(A[11]), .A1(n79) );
  inv01 U35 ( .Y(SUM[11]), .A(n33) );
  xor2 U36 ( .Y(n35), .A0(A[23]), .A1(n81) );
  inv01 U37 ( .Y(SUM[23]), .A(n35) );
  xor2 U38 ( .Y(n37), .A0(A[13]), .A1(n69) );
  inv01 U39 ( .Y(SUM[13]), .A(n37) );
  xor2 U40 ( .Y(n39), .A0(A[7]), .A1(n67) );
  inv01 U41 ( .Y(SUM[7]), .A(n39) );
  xor2 U42 ( .Y(n41), .A0(A[6]), .A1(n60) );
  inv01 U43 ( .Y(SUM[6]), .A(n41) );
  xor2 U44 ( .Y(n43), .A0(A[8]), .A1(n70) );
  inv01 U45 ( .Y(SUM[8]), .A(n43) );
  xor2 U46 ( .Y(n45), .A0(A[14]), .A1(n72) );
  inv01 U47 ( .Y(SUM[14]), .A(n45) );
  xor2 U48 ( .Y(n47), .A0(A[3]), .A1(n68) );
  inv01 U49 ( .Y(SUM[3]), .A(n47) );
  xor2 U50 ( .Y(n49), .A0(A[12]), .A1(n62) );
  inv01 U51 ( .Y(SUM[12]), .A(n49) );
  xor2 U52 ( .Y(n51), .A0(A[18]), .A1(n57) );
  inv01 U53 ( .Y(SUM[18]), .A(n51) );
  xor2 U54 ( .Y(n53), .A0(A[19]), .A1(n66) );
  inv01 U55 ( .Y(SUM[19]), .A(n53) );
  buf02 U56 ( .Y(n55), .A(carry_2_) );
  nor02 U57 ( .Y(n56), .A0(A[17]), .A1(n78) );
  inv02 U58 ( .Y(n57), .A(n56) );
  nor02 U59 ( .Y(n58), .A0(A[20]), .A1(n80) );
  inv02 U60 ( .Y(n59), .A(n58) );
  buf02 U61 ( .Y(n60), .A(carry_6_) );
  nor02 U62 ( .Y(n61), .A0(A[11]), .A1(n79) );
  inv02 U63 ( .Y(n62), .A(n61) );
  nor02 U64 ( .Y(n63), .A0(A[23]), .A1(n81) );
  inv02 U65 ( .Y(n64), .A(n63) );
  buf02 U66 ( .Y(n65), .A(carry_22_) );
  buf02 U67 ( .Y(n66), .A(carry_19_) );
  buf02 U68 ( .Y(n67), .A(carry_7_) );
  buf02 U69 ( .Y(n68), .A(carry_3_) );
  buf02 U70 ( .Y(n69), .A(carry_13_) );
  buf02 U71 ( .Y(n70), .A(carry_8_) );
  buf02 U72 ( .Y(n71), .A(carry_4_) );
  buf02 U73 ( .Y(n72), .A(carry_14_) );
  buf02 U74 ( .Y(n73), .A(carry_16_) );
  buf02 U75 ( .Y(n74), .A(carry_9_) );
  buf02 U76 ( .Y(n75), .A(carry_15_) );
  buf02 U77 ( .Y(n76), .A(carry_5_) );
  buf02 U78 ( .Y(n77), .A(carry_10_) );
  buf02 U79 ( .Y(n78), .A(carry_17_) );
  buf02 U80 ( .Y(n79), .A(carry_11_) );
  buf02 U81 ( .Y(n80), .A(carry_20_) );
  buf02 U82 ( .Y(n81), .A(carry_23_) );
  inv01 U83 ( .Y(SUM[0]), .A(A[0]) );
  or02 U1_B_1 ( .Y(carry_2_), .A0(A[1]), .A1(A[0]) );
  or02 U1_B_2 ( .Y(carry_3_), .A0(A[2]), .A1(n55) );
  or02 U1_B_3 ( .Y(carry_4_), .A0(A[3]), .A1(n68) );
  or02 U1_B_4 ( .Y(carry_5_), .A0(A[4]), .A1(n71) );
  or02 U1_B_5 ( .Y(carry_6_), .A0(A[5]), .A1(n76) );
  or02 U1_B_6 ( .Y(carry_7_), .A0(A[6]), .A1(n60) );
  or02 U1_B_7 ( .Y(carry_8_), .A0(A[7]), .A1(n67) );
  or02 U1_B_8 ( .Y(carry_9_), .A0(A[8]), .A1(n70) );
  or02 U1_B_9 ( .Y(carry_10_), .A0(A[9]), .A1(n74) );
  or02 U1_B_10 ( .Y(carry_11_), .A0(A[10]), .A1(n77) );
  or02 U1_B_12 ( .Y(carry_13_), .A0(A[12]), .A1(n62) );
  or02 U1_B_13 ( .Y(carry_14_), .A0(A[13]), .A1(n69) );
  or02 U1_B_14 ( .Y(carry_15_), .A0(A[14]), .A1(n72) );
  or02 U1_B_15 ( .Y(carry_16_), .A0(A[15]), .A1(n75) );
  or02 U1_B_16 ( .Y(carry_17_), .A0(A[16]), .A1(n73) );
  or02 U1_B_18 ( .Y(carry_19_), .A0(A[18]), .A1(n57) );
  or02 U1_B_19 ( .Y(carry_20_), .A0(A[19]), .A1(n66) );
  or02 U1_B_21 ( .Y(carry_22_), .A0(A[21]), .A1(n59) );
  or02 U1_B_22 ( .Y(carry_23_), .A0(A[22]), .A1(n65) );
  or02 U1_B_24 ( .Y(carry_25_), .A0(A[24]), .A1(n64) );
endmodule


module sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_cmp2_52_1 ( A, B, LEQ, TC, LT_LE, GE_GT
 );
  input [51:0] A;
  input [51:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297;

  ao22 U6 ( .Y(n15), .A0(A[51]), .A1(n170), .B0(n171), .B1(n172) );
  inv01 U7 ( .Y(n16), .A(n15) );
  inv01 U8 ( .Y(n171), .A(n17) );
  nor02 U9 ( .Y(n18), .A0(B[50]), .A1(n173) );
  nor02 U10 ( .Y(n19), .A0(B[49]), .A1(n174) );
  inv01 U11 ( .Y(n20), .A(n175) );
  nor02 U12 ( .Y(n17), .A0(n20), .A1(n21) );
  nor02 U13 ( .Y(n22), .A0(n18), .A1(n19) );
  inv01 U14 ( .Y(n21), .A(n22) );
  nand02 U15 ( .Y(n293), .A0(n296), .A1(n23) );
  inv01 U16 ( .Y(n24), .A(n291) );
  inv01 U17 ( .Y(n25), .A(B[2]) );
  inv01 U18 ( .Y(n26), .A(n295) );
  inv01 U19 ( .Y(n27), .A(n294) );
  nand02 U20 ( .Y(n28), .A0(n24), .A1(n25) );
  nand02 U21 ( .Y(n29), .A0(n26), .A1(n27) );
  nand02 U22 ( .Y(n30), .A0(n28), .A1(n29) );
  inv01 U23 ( .Y(n23), .A(n30) );
  inv01 U24 ( .Y(n292), .A(n293) );
  inv01 U25 ( .Y(n295), .A(A[1]) );
  inv01 U26 ( .Y(n291), .A(A[2]) );
  inv01 U27 ( .Y(n228), .A(n31) );
  nor02 U28 ( .Y(n32), .A0(B[28]), .A1(n226) );
  nor02 U29 ( .Y(n33), .A0(B[27]), .A1(n229) );
  inv01 U30 ( .Y(n34), .A(n230) );
  nor02 U31 ( .Y(n31), .A0(n34), .A1(n35) );
  nor02 U32 ( .Y(n36), .A0(n32), .A1(n33) );
  inv01 U33 ( .Y(n35), .A(n36) );
  inv01 U34 ( .Y(n243), .A(n37) );
  nor02 U35 ( .Y(n38), .A0(B[22]), .A1(n241) );
  nor02 U36 ( .Y(n39), .A0(B[21]), .A1(n244) );
  inv01 U37 ( .Y(n40), .A(n245) );
  nor02 U38 ( .Y(n37), .A0(n40), .A1(n41) );
  nor02 U39 ( .Y(n42), .A0(n38), .A1(n39) );
  inv01 U40 ( .Y(n41), .A(n42) );
  inv01 U41 ( .Y(n227), .A(n228) );
  inv01 U42 ( .Y(n242), .A(n243) );
  inv01 U43 ( .Y(n258), .A(n43) );
  nor02 U44 ( .Y(n44), .A0(B[16]), .A1(n256) );
  nor02 U45 ( .Y(n45), .A0(B[15]), .A1(n259) );
  inv01 U46 ( .Y(n46), .A(n260) );
  nor02 U47 ( .Y(n43), .A0(n46), .A1(n47) );
  nor02 U48 ( .Y(n48), .A0(n44), .A1(n45) );
  inv01 U49 ( .Y(n47), .A(n48) );
  inv01 U50 ( .Y(n273), .A(n49) );
  nor02 U51 ( .Y(n50), .A0(B[9]), .A1(n274) );
  nor02 U52 ( .Y(n51), .A0(B[10]), .A1(n271) );
  inv01 U53 ( .Y(n52), .A(n275) );
  nor02 U54 ( .Y(n49), .A0(n52), .A1(n53) );
  nor02 U55 ( .Y(n54), .A0(n50), .A1(n51) );
  inv01 U56 ( .Y(n53), .A(n54) );
  inv01 U57 ( .Y(n257), .A(n258) );
  inv01 U58 ( .Y(n272), .A(n273) );
  inv01 U59 ( .Y(n218), .A(n55) );
  nor02 U60 ( .Y(n56), .A0(B[32]), .A1(n216) );
  nor02 U61 ( .Y(n57), .A0(B[31]), .A1(n219) );
  inv01 U62 ( .Y(n58), .A(n220) );
  nor02 U63 ( .Y(n55), .A0(n58), .A1(n59) );
  nor02 U64 ( .Y(n60), .A0(n56), .A1(n57) );
  inv01 U65 ( .Y(n59), .A(n60) );
  inv01 U66 ( .Y(n188), .A(n61) );
  nor02 U67 ( .Y(n62), .A0(B[44]), .A1(n186) );
  nor02 U68 ( .Y(n63), .A0(B[43]), .A1(n189) );
  inv01 U69 ( .Y(n64), .A(n190) );
  nor02 U70 ( .Y(n61), .A0(n64), .A1(n65) );
  nor02 U71 ( .Y(n66), .A0(n62), .A1(n63) );
  inv01 U72 ( .Y(n65), .A(n66) );
  inv01 U73 ( .Y(n217), .A(n218) );
  inv01 U74 ( .Y(n187), .A(n188) );
  inv02 U75 ( .Y(n186), .A(A[44]) );
  inv01 U76 ( .Y(n283), .A(n67) );
  nor02 U77 ( .Y(n68), .A0(B[6]), .A1(n281) );
  nor02 U78 ( .Y(n69), .A0(B[5]), .A1(n284) );
  inv01 U79 ( .Y(n70), .A(n285) );
  nor02 U80 ( .Y(n67), .A0(n70), .A1(n71) );
  nor02 U81 ( .Y(n72), .A0(n68), .A1(n69) );
  inv01 U82 ( .Y(n71), .A(n72) );
  inv01 U83 ( .Y(n198), .A(n73) );
  nor02 U84 ( .Y(n74), .A0(B[40]), .A1(n196) );
  nor02 U85 ( .Y(n75), .A0(B[39]), .A1(n199) );
  inv01 U86 ( .Y(n76), .A(n200) );
  nor02 U87 ( .Y(n73), .A0(n76), .A1(n77) );
  nor02 U88 ( .Y(n78), .A0(n74), .A1(n75) );
  inv01 U89 ( .Y(n77), .A(n78) );
  inv01 U90 ( .Y(n282), .A(n283) );
  inv01 U91 ( .Y(n197), .A(n198) );
  inv01 U92 ( .Y(n183), .A(n79) );
  nor02 U93 ( .Y(n80), .A0(B[46]), .A1(n181) );
  nor02 U94 ( .Y(n81), .A0(B[45]), .A1(n184) );
  inv01 U95 ( .Y(n82), .A(n185) );
  nor02 U96 ( .Y(n79), .A0(n82), .A1(n83) );
  nor02 U97 ( .Y(n84), .A0(n80), .A1(n81) );
  inv01 U98 ( .Y(n83), .A(n84) );
  inv01 U99 ( .Y(n213), .A(n85) );
  nor02 U100 ( .Y(n86), .A0(B[34]), .A1(n211) );
  nor02 U101 ( .Y(n87), .A0(B[33]), .A1(n214) );
  inv01 U102 ( .Y(n88), .A(n215) );
  nor02 U103 ( .Y(n85), .A0(n88), .A1(n89) );
  nor02 U104 ( .Y(n90), .A0(n86), .A1(n87) );
  inv01 U105 ( .Y(n89), .A(n90) );
  inv01 U106 ( .Y(n182), .A(n183) );
  inv01 U107 ( .Y(n212), .A(n213) );
  inv01 U108 ( .Y(n248), .A(n91) );
  nor02 U109 ( .Y(n92), .A0(B[20]), .A1(n246) );
  nor02 U110 ( .Y(n93), .A0(B[19]), .A1(n249) );
  inv01 U111 ( .Y(n94), .A(n250) );
  nor02 U112 ( .Y(n91), .A0(n94), .A1(n95) );
  nor02 U113 ( .Y(n96), .A0(n92), .A1(n93) );
  inv01 U114 ( .Y(n95), .A(n96) );
  inv01 U115 ( .Y(n247), .A(n248) );
  inv01 U116 ( .Y(n268), .A(n97) );
  nor02 U117 ( .Y(n98), .A0(B[12]), .A1(n266) );
  nor02 U118 ( .Y(n99), .A0(B[11]), .A1(n269) );
  inv01 U119 ( .Y(n100), .A(n270) );
  nor02 U120 ( .Y(n97), .A0(n100), .A1(n101) );
  nor02 U121 ( .Y(n102), .A0(n98), .A1(n99) );
  inv01 U122 ( .Y(n101), .A(n102) );
  inv01 U123 ( .Y(n203), .A(n103) );
  nor02 U124 ( .Y(n104), .A0(B[38]), .A1(n201) );
  nor02 U125 ( .Y(n105), .A0(B[37]), .A1(n204) );
  inv01 U126 ( .Y(n106), .A(n205) );
  nor02 U127 ( .Y(n103), .A0(n106), .A1(n107) );
  nor02 U128 ( .Y(n108), .A0(n104), .A1(n105) );
  inv01 U129 ( .Y(n107), .A(n108) );
  inv01 U130 ( .Y(n267), .A(n268) );
  inv01 U131 ( .Y(n202), .A(n203) );
  inv01 U132 ( .Y(n223), .A(n109) );
  nor02 U133 ( .Y(n110), .A0(B[30]), .A1(n221) );
  nor02 U134 ( .Y(n111), .A0(B[29]), .A1(n224) );
  inv01 U135 ( .Y(n112), .A(n225) );
  nor02 U136 ( .Y(n109), .A0(n112), .A1(n113) );
  nor02 U137 ( .Y(n114), .A0(n110), .A1(n111) );
  inv01 U138 ( .Y(n113), .A(n114) );
  inv01 U139 ( .Y(n278), .A(n115) );
  nor02 U140 ( .Y(n116), .A0(B[8]), .A1(n276) );
  nor02 U141 ( .Y(n117), .A0(B[7]), .A1(n279) );
  inv01 U142 ( .Y(n118), .A(n280) );
  nor02 U143 ( .Y(n115), .A0(n118), .A1(n119) );
  nor02 U144 ( .Y(n120), .A0(n116), .A1(n117) );
  inv01 U145 ( .Y(n119), .A(n120) );
  inv01 U146 ( .Y(n222), .A(n223) );
  inv01 U147 ( .Y(n277), .A(n278) );
  inv01 U148 ( .Y(n238), .A(n121) );
  nor02 U149 ( .Y(n122), .A0(B[24]), .A1(n236) );
  nor02 U150 ( .Y(n123), .A0(B[23]), .A1(n239) );
  inv01 U151 ( .Y(n124), .A(n240) );
  nor02 U152 ( .Y(n121), .A0(n124), .A1(n125) );
  nor02 U153 ( .Y(n126), .A0(n122), .A1(n123) );
  inv01 U154 ( .Y(n125), .A(n126) );
  inv01 U155 ( .Y(n193), .A(n127) );
  nor02 U156 ( .Y(n128), .A0(B[42]), .A1(n191) );
  nor02 U157 ( .Y(n129), .A0(B[41]), .A1(n194) );
  inv01 U158 ( .Y(n130), .A(n195) );
  nor02 U159 ( .Y(n127), .A0(n130), .A1(n131) );
  nor02 U160 ( .Y(n132), .A0(n128), .A1(n129) );
  inv01 U161 ( .Y(n131), .A(n132) );
  inv01 U162 ( .Y(n237), .A(n238) );
  inv01 U163 ( .Y(n192), .A(n193) );
  inv01 U164 ( .Y(n288), .A(n133) );
  nor02 U165 ( .Y(n134), .A0(B[4]), .A1(n286) );
  nor02 U166 ( .Y(n135), .A0(B[3]), .A1(n289) );
  inv01 U167 ( .Y(n136), .A(n290) );
  nor02 U168 ( .Y(n133), .A0(n136), .A1(n137) );
  nor02 U169 ( .Y(n138), .A0(n134), .A1(n135) );
  inv01 U170 ( .Y(n137), .A(n138) );
  inv01 U171 ( .Y(n263), .A(n139) );
  nor02 U172 ( .Y(n140), .A0(B[14]), .A1(n261) );
  nor02 U173 ( .Y(n141), .A0(B[13]), .A1(n264) );
  inv01 U174 ( .Y(n142), .A(n265) );
  nor02 U175 ( .Y(n139), .A0(n142), .A1(n143) );
  nor02 U176 ( .Y(n144), .A0(n140), .A1(n141) );
  inv01 U177 ( .Y(n143), .A(n144) );
  inv01 U178 ( .Y(n287), .A(n288) );
  inv01 U179 ( .Y(n262), .A(n263) );
  inv01 U180 ( .Y(n253), .A(n145) );
  nor02 U181 ( .Y(n146), .A0(B[18]), .A1(n251) );
  nor02 U182 ( .Y(n147), .A0(B[17]), .A1(n254) );
  inv01 U183 ( .Y(n148), .A(n255) );
  nor02 U184 ( .Y(n145), .A0(n148), .A1(n149) );
  nor02 U185 ( .Y(n150), .A0(n146), .A1(n147) );
  inv01 U186 ( .Y(n149), .A(n150) );
  inv01 U187 ( .Y(n208), .A(n151) );
  nor02 U188 ( .Y(n152), .A0(B[36]), .A1(n206) );
  nor02 U189 ( .Y(n153), .A0(B[35]), .A1(n209) );
  inv01 U190 ( .Y(n154), .A(n210) );
  nor02 U191 ( .Y(n151), .A0(n154), .A1(n155) );
  nor02 U192 ( .Y(n156), .A0(n152), .A1(n153) );
  inv01 U193 ( .Y(n155), .A(n156) );
  inv01 U194 ( .Y(n252), .A(n253) );
  inv01 U195 ( .Y(n207), .A(n208) );
  inv01 U196 ( .Y(n178), .A(n157) );
  nor02 U197 ( .Y(n158), .A0(B[48]), .A1(n176) );
  nor02 U198 ( .Y(n159), .A0(B[47]), .A1(n179) );
  inv01 U199 ( .Y(n160), .A(n180) );
  nor02 U200 ( .Y(n157), .A0(n160), .A1(n161) );
  nor02 U201 ( .Y(n162), .A0(n158), .A1(n159) );
  inv01 U202 ( .Y(n161), .A(n162) );
  inv01 U203 ( .Y(n233), .A(n163) );
  nor02 U204 ( .Y(n164), .A0(B[26]), .A1(n231) );
  nor02 U205 ( .Y(n165), .A0(B[25]), .A1(n234) );
  inv01 U206 ( .Y(n166), .A(n235) );
  nor02 U207 ( .Y(n163), .A0(n166), .A1(n167) );
  nor02 U208 ( .Y(n168), .A0(n164), .A1(n165) );
  inv01 U209 ( .Y(n167), .A(n168) );
  inv01 U210 ( .Y(n177), .A(n178) );
  inv01 U211 ( .Y(n232), .A(n233) );
  inv01 U212 ( .Y(n224), .A(A[29]) );
  inv02 U213 ( .Y(n206), .A(A[36]) );
  inv02 U214 ( .Y(n241), .A(A[22]) );
  inv02 U215 ( .Y(n181), .A(A[46]) );
  inv02 U216 ( .Y(n276), .A(A[8]) );
  inv02 U217 ( .Y(n266), .A(A[12]) );
  inv02 U218 ( .Y(n236), .A(A[24]) );
  inv01 U219 ( .Y(n194), .A(A[41]) );
  inv01 U220 ( .Y(n239), .A(A[23]) );
  inv02 U221 ( .Y(n211), .A(A[34]) );
  inv02 U222 ( .Y(n256), .A(A[16]) );
  inv01 U223 ( .Y(n209), .A(A[35]) );
  inv01 U224 ( .Y(n184), .A(A[45]) );
  inv01 U225 ( .Y(n269), .A(A[11]) );
  inv02 U226 ( .Y(n251), .A(A[18]) );
  inv01 U227 ( .Y(n279), .A(A[7]) );
  inv01 U228 ( .Y(n214), .A(A[33]) );
  inv02 U229 ( .Y(n176), .A(A[48]) );
  inv01 U230 ( .Y(n244), .A(A[21]) );
  inv01 U231 ( .Y(n289), .A(A[3]) );
  inv01 U232 ( .Y(n271), .A(A[10]) );
  inv02 U233 ( .Y(n226), .A(A[28]) );
  inv02 U234 ( .Y(n196), .A(A[40]) );
  inv01 U235 ( .Y(n204), .A(A[37]) );
  inv01 U236 ( .Y(n179), .A(A[47]) );
  inv01 U237 ( .Y(n254), .A(A[17]) );
  inv02 U238 ( .Y(n281), .A(A[6]) );
  inv02 U239 ( .Y(n274), .A(A[9]) );
  inv01 U240 ( .Y(n229), .A(A[27]) );
  inv02 U241 ( .Y(n201), .A(A[38]) );
  inv02 U242 ( .Y(n173), .A(A[50]) );
  inv01 U243 ( .Y(n259), .A(A[15]) );
  inv01 U244 ( .Y(n249), .A(A[19]) );
  inv01 U245 ( .Y(n284), .A(A[5]) );
  inv02 U246 ( .Y(n246), .A(A[20]) );
  inv01 U247 ( .Y(n189), .A(A[43]) );
  inv02 U248 ( .Y(n216), .A(A[32]) );
  inv01 U249 ( .Y(n234), .A(A[25]) );
  inv01 U250 ( .Y(n264), .A(A[13]) );
  inv01 U251 ( .Y(n219), .A(A[31]) );
  inv02 U252 ( .Y(n221), .A(A[30]) );
  inv01 U253 ( .Y(n174), .A(A[49]) );
  inv02 U254 ( .Y(n286), .A(A[4]) );
  inv02 U255 ( .Y(n261), .A(A[14]) );
  inv02 U256 ( .Y(n231), .A(A[26]) );
  inv02 U257 ( .Y(n191), .A(A[42]) );
  inv01 U258 ( .Y(n199), .A(A[39]) );
  inv01 U259 ( .Y(n169), .A(A[51]) );
  inv01 U260 ( .Y(n297), .A(B[0]) );
  inv01 U261 ( .Y(n170), .A(B[51]) );
  ao21 U262 ( .Y(LT_LE), .A0(B[51]), .A1(n169), .B0(n16) );
  nand02 U263 ( .Y(n172), .A0(B[50]), .A1(n173) );
  ao221 U264 ( .Y(n175), .A0(n176), .A1(B[48]), .B0(n174), .B1(B[49]), .C0(
        n177) );
  ao221 U265 ( .Y(n180), .A0(n181), .A1(B[46]), .B0(n179), .B1(B[47]), .C0(
        n182) );
  ao221 U266 ( .Y(n185), .A0(n186), .A1(B[44]), .B0(n184), .B1(B[45]), .C0(
        n187) );
  ao221 U267 ( .Y(n190), .A0(n191), .A1(B[42]), .B0(n189), .B1(B[43]), .C0(
        n192) );
  ao221 U268 ( .Y(n195), .A0(n196), .A1(B[40]), .B0(n194), .B1(B[41]), .C0(
        n197) );
  ao221 U269 ( .Y(n200), .A0(n201), .A1(B[38]), .B0(n199), .B1(B[39]), .C0(
        n202) );
  ao221 U270 ( .Y(n205), .A0(n206), .A1(B[36]), .B0(n204), .B1(B[37]), .C0(
        n207) );
  ao221 U271 ( .Y(n210), .A0(n211), .A1(B[34]), .B0(n209), .B1(B[35]), .C0(
        n212) );
  ao221 U272 ( .Y(n215), .A0(n216), .A1(B[32]), .B0(n214), .B1(B[33]), .C0(
        n217) );
  ao221 U273 ( .Y(n220), .A0(n221), .A1(B[30]), .B0(n219), .B1(B[31]), .C0(
        n222) );
  ao221 U274 ( .Y(n225), .A0(n226), .A1(B[28]), .B0(n224), .B1(B[29]), .C0(
        n227) );
  ao221 U275 ( .Y(n230), .A0(n231), .A1(B[26]), .B0(n229), .B1(B[27]), .C0(
        n232) );
  ao221 U276 ( .Y(n235), .A0(n236), .A1(B[24]), .B0(n234), .B1(B[25]), .C0(
        n237) );
  ao221 U277 ( .Y(n240), .A0(n241), .A1(B[22]), .B0(n239), .B1(B[23]), .C0(
        n242) );
  ao221 U278 ( .Y(n245), .A0(n246), .A1(B[20]), .B0(n244), .B1(B[21]), .C0(
        n247) );
  ao221 U279 ( .Y(n250), .A0(n251), .A1(B[18]), .B0(n249), .B1(B[19]), .C0(
        n252) );
  ao221 U280 ( .Y(n255), .A0(n256), .A1(B[16]), .B0(n254), .B1(B[17]), .C0(
        n257) );
  ao221 U281 ( .Y(n260), .A0(n261), .A1(B[14]), .B0(n259), .B1(B[15]), .C0(
        n262) );
  ao221 U282 ( .Y(n265), .A0(n266), .A1(B[12]), .B0(n264), .B1(B[13]), .C0(
        n267) );
  ao221 U283 ( .Y(n270), .A0(n271), .A1(B[10]), .B0(n269), .B1(B[11]), .C0(
        n272) );
  ao221 U284 ( .Y(n275), .A0(n276), .A1(B[8]), .B0(n274), .B1(B[9]), .C0(n277)
         );
  ao221 U285 ( .Y(n280), .A0(n281), .A1(B[6]), .B0(n279), .B1(B[7]), .C0(n282)
         );
  ao221 U286 ( .Y(n285), .A0(n286), .A1(B[4]), .B0(n284), .B1(B[5]), .C0(n287)
         );
  ao221 U287 ( .Y(n290), .A0(n291), .A1(B[2]), .B0(n289), .B1(B[3]), .C0(n292)
         );
  ao21 U288 ( .Y(n296), .A0(n294), .A1(n295), .B0(B[1]) );
  nor02 U289 ( .Y(n294), .A0(n297), .A1(A[0]) );
endmodule


module sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_cmp2_52_0 ( A, B, LEQ, TC, LT_LE, GE_GT
 );
  input [51:0] A;
  input [51:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301;

  buf02 U6 ( .Y(n15), .A(n173) );
  inv01 U7 ( .Y(n175), .A(n16) );
  nor02 U8 ( .Y(n17), .A0(B[50]), .A1(n177) );
  nor02 U9 ( .Y(n18), .A0(B[49]), .A1(n178) );
  inv01 U10 ( .Y(n19), .A(n179) );
  nor02 U11 ( .Y(n16), .A0(n19), .A1(n20) );
  nor02 U12 ( .Y(n21), .A0(n17), .A1(n18) );
  inv01 U13 ( .Y(n20), .A(n21) );
  nand02 U14 ( .Y(n297), .A0(n300), .A1(n22) );
  inv01 U15 ( .Y(n23), .A(n295) );
  inv01 U16 ( .Y(n24), .A(B[2]) );
  inv01 U17 ( .Y(n25), .A(n299) );
  inv01 U18 ( .Y(n26), .A(n298) );
  nand02 U19 ( .Y(n27), .A0(n23), .A1(n24) );
  nand02 U20 ( .Y(n28), .A0(n25), .A1(n26) );
  nand02 U21 ( .Y(n29), .A0(n27), .A1(n28) );
  inv01 U22 ( .Y(n22), .A(n29) );
  inv01 U23 ( .Y(n296), .A(n297) );
  inv01 U24 ( .Y(n277), .A(n30) );
  nor02 U25 ( .Y(n31), .A0(B[9]), .A1(n278) );
  nor02 U26 ( .Y(n32), .A0(B[10]), .A1(n275) );
  inv01 U27 ( .Y(n33), .A(n279) );
  nor02 U28 ( .Y(n30), .A0(n33), .A1(n34) );
  nor02 U29 ( .Y(n35), .A0(n31), .A1(n32) );
  inv01 U30 ( .Y(n34), .A(n35) );
  inv01 U31 ( .Y(n252), .A(n36) );
  nor02 U32 ( .Y(n37), .A0(B[20]), .A1(n250) );
  nor02 U33 ( .Y(n38), .A0(B[19]), .A1(n253) );
  inv01 U34 ( .Y(n39), .A(n254) );
  nor02 U35 ( .Y(n36), .A0(n39), .A1(n40) );
  nor02 U36 ( .Y(n41), .A0(n37), .A1(n38) );
  inv01 U37 ( .Y(n40), .A(n41) );
  inv01 U38 ( .Y(n276), .A(n277) );
  inv01 U39 ( .Y(n251), .A(n252) );
  inv01 U40 ( .Y(n212), .A(n42) );
  nor02 U41 ( .Y(n43), .A0(B[36]), .A1(n210) );
  nor02 U42 ( .Y(n44), .A0(B[35]), .A1(n213) );
  inv01 U43 ( .Y(n45), .A(n214) );
  nor02 U44 ( .Y(n42), .A0(n45), .A1(n46) );
  nor02 U45 ( .Y(n47), .A0(n43), .A1(n44) );
  inv01 U46 ( .Y(n46), .A(n47) );
  inv01 U47 ( .Y(n287), .A(n48) );
  nor02 U48 ( .Y(n49), .A0(B[6]), .A1(n285) );
  nor02 U49 ( .Y(n50), .A0(B[5]), .A1(n288) );
  inv01 U50 ( .Y(n51), .A(n289) );
  nor02 U51 ( .Y(n48), .A0(n51), .A1(n52) );
  nor02 U52 ( .Y(n53), .A0(n49), .A1(n50) );
  inv01 U53 ( .Y(n52), .A(n53) );
  inv01 U54 ( .Y(n211), .A(n212) );
  inv01 U55 ( .Y(n210), .A(A[36]) );
  inv01 U56 ( .Y(n286), .A(n287) );
  inv01 U57 ( .Y(n285), .A(A[6]) );
  inv01 U58 ( .Y(n202), .A(n54) );
  nor02 U59 ( .Y(n55), .A0(B[40]), .A1(n200) );
  nor02 U60 ( .Y(n56), .A0(B[39]), .A1(n203) );
  inv01 U61 ( .Y(n57), .A(n204) );
  nor02 U62 ( .Y(n54), .A0(n57), .A1(n58) );
  nor02 U63 ( .Y(n59), .A0(n55), .A1(n56) );
  inv01 U64 ( .Y(n58), .A(n59) );
  inv01 U65 ( .Y(n192), .A(n60) );
  nor02 U66 ( .Y(n61), .A0(B[44]), .A1(n190) );
  nor02 U67 ( .Y(n62), .A0(B[43]), .A1(n193) );
  inv01 U68 ( .Y(n63), .A(n194) );
  nor02 U69 ( .Y(n60), .A0(n63), .A1(n64) );
  nor02 U70 ( .Y(n65), .A0(n61), .A1(n62) );
  inv01 U71 ( .Y(n64), .A(n65) );
  inv01 U72 ( .Y(n201), .A(n202) );
  inv01 U73 ( .Y(n200), .A(A[40]) );
  inv01 U74 ( .Y(n191), .A(n192) );
  inv02 U75 ( .Y(n190), .A(A[44]) );
  inv01 U76 ( .Y(n222), .A(n66) );
  nor02 U77 ( .Y(n67), .A0(B[32]), .A1(n220) );
  nor02 U78 ( .Y(n68), .A0(B[31]), .A1(n223) );
  inv01 U79 ( .Y(n69), .A(n224) );
  nor02 U80 ( .Y(n66), .A0(n69), .A1(n70) );
  nor02 U81 ( .Y(n71), .A0(n67), .A1(n68) );
  inv01 U82 ( .Y(n70), .A(n71) );
  inv01 U83 ( .Y(n262), .A(n72) );
  nor02 U84 ( .Y(n73), .A0(B[16]), .A1(n260) );
  nor02 U85 ( .Y(n74), .A0(B[15]), .A1(n263) );
  inv01 U86 ( .Y(n75), .A(n264) );
  nor02 U87 ( .Y(n72), .A0(n75), .A1(n76) );
  nor02 U88 ( .Y(n77), .A0(n73), .A1(n74) );
  inv01 U89 ( .Y(n76), .A(n77) );
  inv01 U90 ( .Y(n221), .A(n222) );
  inv01 U91 ( .Y(n261), .A(n262) );
  inv01 U92 ( .Y(n260), .A(A[16]) );
  inv01 U93 ( .Y(n247), .A(n78) );
  nor02 U94 ( .Y(n79), .A0(B[22]), .A1(n245) );
  nor02 U95 ( .Y(n80), .A0(B[21]), .A1(n248) );
  inv01 U96 ( .Y(n81), .A(n249) );
  nor02 U97 ( .Y(n78), .A0(n81), .A1(n82) );
  nor02 U98 ( .Y(n83), .A0(n79), .A1(n80) );
  inv01 U99 ( .Y(n82), .A(n83) );
  inv01 U100 ( .Y(n272), .A(n84) );
  nor02 U101 ( .Y(n85), .A0(B[12]), .A1(n270) );
  nor02 U102 ( .Y(n86), .A0(B[11]), .A1(n273) );
  inv01 U103 ( .Y(n87), .A(n274) );
  nor02 U104 ( .Y(n84), .A0(n87), .A1(n88) );
  nor02 U105 ( .Y(n89), .A0(n85), .A1(n86) );
  inv01 U106 ( .Y(n88), .A(n89) );
  inv01 U107 ( .Y(n246), .A(n247) );
  inv01 U108 ( .Y(n245), .A(A[22]) );
  inv01 U109 ( .Y(n271), .A(n272) );
  inv01 U110 ( .Y(n242), .A(n90) );
  nor02 U111 ( .Y(n91), .A0(B[24]), .A1(n240) );
  nor02 U112 ( .Y(n92), .A0(B[23]), .A1(n243) );
  inv01 U113 ( .Y(n93), .A(n244) );
  nor02 U114 ( .Y(n90), .A0(n93), .A1(n94) );
  nor02 U115 ( .Y(n95), .A0(n91), .A1(n92) );
  inv01 U116 ( .Y(n94), .A(n95) );
  inv01 U117 ( .Y(n217), .A(n96) );
  nor02 U118 ( .Y(n97), .A0(B[34]), .A1(n215) );
  nor02 U119 ( .Y(n98), .A0(B[33]), .A1(n218) );
  inv01 U120 ( .Y(n99), .A(n219) );
  nor02 U121 ( .Y(n96), .A0(n99), .A1(n100) );
  nor02 U122 ( .Y(n101), .A0(n97), .A1(n98) );
  inv01 U123 ( .Y(n100), .A(n101) );
  inv01 U124 ( .Y(n241), .A(n242) );
  inv01 U125 ( .Y(n216), .A(n217) );
  inv01 U126 ( .Y(n215), .A(A[34]) );
  inv01 U127 ( .Y(n187), .A(n102) );
  nor02 U128 ( .Y(n103), .A0(B[46]), .A1(n185) );
  nor02 U129 ( .Y(n104), .A0(B[45]), .A1(n188) );
  inv01 U130 ( .Y(n105), .A(n189) );
  nor02 U131 ( .Y(n102), .A0(n105), .A1(n106) );
  nor02 U132 ( .Y(n107), .A0(n103), .A1(n104) );
  inv01 U133 ( .Y(n106), .A(n107) );
  inv01 U134 ( .Y(n292), .A(n108) );
  nor02 U135 ( .Y(n109), .A0(B[4]), .A1(n290) );
  nor02 U136 ( .Y(n110), .A0(B[3]), .A1(n293) );
  inv01 U137 ( .Y(n111), .A(n294) );
  nor02 U138 ( .Y(n108), .A0(n111), .A1(n112) );
  nor02 U139 ( .Y(n113), .A0(n109), .A1(n110) );
  inv01 U140 ( .Y(n112), .A(n113) );
  inv01 U141 ( .Y(n186), .A(n187) );
  inv01 U142 ( .Y(n185), .A(A[46]) );
  inv01 U143 ( .Y(n291), .A(n292) );
  inv01 U144 ( .Y(n257), .A(n114) );
  nor02 U145 ( .Y(n115), .A0(B[18]), .A1(n255) );
  nor02 U146 ( .Y(n116), .A0(B[17]), .A1(n258) );
  inv01 U147 ( .Y(n117), .A(n259) );
  nor02 U148 ( .Y(n114), .A0(n117), .A1(n118) );
  nor02 U149 ( .Y(n119), .A0(n115), .A1(n116) );
  inv01 U150 ( .Y(n118), .A(n119) );
  inv01 U151 ( .Y(n282), .A(n120) );
  nor02 U152 ( .Y(n121), .A0(B[8]), .A1(n280) );
  nor02 U153 ( .Y(n122), .A0(B[7]), .A1(n283) );
  inv01 U154 ( .Y(n123), .A(n284) );
  nor02 U155 ( .Y(n120), .A0(n123), .A1(n124) );
  nor02 U156 ( .Y(n125), .A0(n121), .A1(n122) );
  inv01 U157 ( .Y(n124), .A(n125) );
  inv01 U158 ( .Y(n256), .A(n257) );
  inv01 U159 ( .Y(n255), .A(A[18]) );
  inv01 U160 ( .Y(n281), .A(n282) );
  inv01 U161 ( .Y(n232), .A(n126) );
  nor02 U162 ( .Y(n127), .A0(B[28]), .A1(n230) );
  nor02 U163 ( .Y(n128), .A0(B[27]), .A1(n233) );
  inv01 U164 ( .Y(n129), .A(n234) );
  nor02 U165 ( .Y(n126), .A0(n129), .A1(n130) );
  nor02 U166 ( .Y(n131), .A0(n127), .A1(n128) );
  inv01 U167 ( .Y(n130), .A(n131) );
  inv01 U168 ( .Y(n237), .A(n132) );
  nor02 U169 ( .Y(n133), .A0(B[26]), .A1(n235) );
  nor02 U170 ( .Y(n134), .A0(B[25]), .A1(n238) );
  inv01 U171 ( .Y(n135), .A(n239) );
  nor02 U172 ( .Y(n132), .A0(n135), .A1(n136) );
  nor02 U173 ( .Y(n137), .A0(n133), .A1(n134) );
  inv01 U174 ( .Y(n136), .A(n137) );
  inv01 U175 ( .Y(n231), .A(n232) );
  inv01 U176 ( .Y(n230), .A(A[28]) );
  inv01 U177 ( .Y(n236), .A(n237) );
  inv01 U178 ( .Y(n207), .A(n138) );
  nor02 U179 ( .Y(n139), .A0(B[38]), .A1(n205) );
  nor02 U180 ( .Y(n140), .A0(B[37]), .A1(n208) );
  inv01 U181 ( .Y(n141), .A(n209) );
  nor02 U182 ( .Y(n138), .A0(n141), .A1(n142) );
  nor02 U183 ( .Y(n143), .A0(n139), .A1(n140) );
  inv01 U184 ( .Y(n142), .A(n143) );
  inv01 U185 ( .Y(n197), .A(n144) );
  nor02 U186 ( .Y(n145), .A0(B[42]), .A1(n195) );
  nor02 U187 ( .Y(n146), .A0(B[41]), .A1(n198) );
  inv01 U188 ( .Y(n147), .A(n199) );
  nor02 U189 ( .Y(n144), .A0(n147), .A1(n148) );
  nor02 U190 ( .Y(n149), .A0(n145), .A1(n146) );
  inv01 U191 ( .Y(n148), .A(n149) );
  inv01 U192 ( .Y(n206), .A(n207) );
  inv01 U193 ( .Y(n196), .A(n197) );
  inv01 U194 ( .Y(n227), .A(n150) );
  nor02 U195 ( .Y(n151), .A0(B[30]), .A1(n225) );
  nor02 U196 ( .Y(n152), .A0(B[29]), .A1(n228) );
  inv01 U197 ( .Y(n153), .A(n229) );
  nor02 U198 ( .Y(n150), .A0(n153), .A1(n154) );
  nor02 U199 ( .Y(n155), .A0(n151), .A1(n152) );
  inv01 U200 ( .Y(n154), .A(n155) );
  inv01 U201 ( .Y(n267), .A(n156) );
  nor02 U202 ( .Y(n157), .A0(B[14]), .A1(n265) );
  nor02 U203 ( .Y(n158), .A0(B[13]), .A1(n268) );
  inv01 U204 ( .Y(n159), .A(n269) );
  nor02 U205 ( .Y(n156), .A0(n159), .A1(n160) );
  nor02 U206 ( .Y(n161), .A0(n157), .A1(n158) );
  inv01 U207 ( .Y(n160), .A(n161) );
  inv01 U208 ( .Y(n226), .A(n227) );
  inv01 U209 ( .Y(n225), .A(A[30]) );
  inv01 U210 ( .Y(n266), .A(n267) );
  inv01 U211 ( .Y(n182), .A(n162) );
  nor02 U212 ( .Y(n163), .A0(B[48]), .A1(n180) );
  nor02 U213 ( .Y(n164), .A0(B[47]), .A1(n183) );
  inv01 U214 ( .Y(n165), .A(n184) );
  nor02 U215 ( .Y(n162), .A0(n165), .A1(n166) );
  nor02 U216 ( .Y(n167), .A0(n163), .A1(n164) );
  inv01 U217 ( .Y(n166), .A(n167) );
  inv01 U218 ( .Y(n181), .A(n182) );
  inv01 U219 ( .Y(n180), .A(A[48]) );
  inv01 U220 ( .Y(n228), .A(A[29]) );
  inv02 U221 ( .Y(n280), .A(A[8]) );
  inv02 U222 ( .Y(n270), .A(A[12]) );
  inv02 U223 ( .Y(n240), .A(A[24]) );
  inv01 U224 ( .Y(n198), .A(A[41]) );
  inv01 U225 ( .Y(n243), .A(A[23]) );
  inv01 U226 ( .Y(n213), .A(A[35]) );
  inv01 U227 ( .Y(n188), .A(A[45]) );
  inv01 U228 ( .Y(n273), .A(A[11]) );
  inv02 U229 ( .Y(n295), .A(A[2]) );
  inv01 U230 ( .Y(n283), .A(A[7]) );
  inv01 U231 ( .Y(n218), .A(A[33]) );
  inv01 U232 ( .Y(n248), .A(A[21]) );
  inv01 U233 ( .Y(n293), .A(A[3]) );
  inv01 U234 ( .Y(n275), .A(A[10]) );
  inv01 U235 ( .Y(n208), .A(A[37]) );
  inv01 U236 ( .Y(n183), .A(A[47]) );
  inv01 U237 ( .Y(n258), .A(A[17]) );
  inv02 U238 ( .Y(n278), .A(A[9]) );
  inv01 U239 ( .Y(n233), .A(A[27]) );
  inv02 U240 ( .Y(n205), .A(A[38]) );
  inv02 U241 ( .Y(n177), .A(A[50]) );
  inv01 U242 ( .Y(n263), .A(A[15]) );
  inv01 U243 ( .Y(n253), .A(A[19]) );
  inv01 U244 ( .Y(n288), .A(A[5]) );
  inv02 U245 ( .Y(n299), .A(A[1]) );
  inv02 U246 ( .Y(n250), .A(A[20]) );
  inv01 U247 ( .Y(n193), .A(A[43]) );
  inv02 U248 ( .Y(n220), .A(A[32]) );
  inv01 U249 ( .Y(n238), .A(A[25]) );
  inv01 U250 ( .Y(n268), .A(A[13]) );
  inv01 U251 ( .Y(n223), .A(A[31]) );
  inv01 U252 ( .Y(n178), .A(A[49]) );
  inv02 U253 ( .Y(n290), .A(A[4]) );
  inv02 U254 ( .Y(n265), .A(A[14]) );
  inv02 U255 ( .Y(n235), .A(A[26]) );
  inv02 U256 ( .Y(n195), .A(A[42]) );
  inv01 U257 ( .Y(n203), .A(A[39]) );
  inv02 U258 ( .Y(LT_LE), .A(n168) );
  inv01 U259 ( .Y(n169), .A(n172) );
  inv01 U260 ( .Y(n170), .A(B[51]) );
  nor02 U261 ( .Y(n171), .A0(n169), .A1(n170) );
  nor02 U262 ( .Y(n168), .A0(n171), .A1(n15) );
  inv01 U263 ( .Y(n172), .A(A[51]) );
  inv04 U264 ( .Y(n301), .A(B[0]) );
  inv04 U265 ( .Y(n174), .A(B[51]) );
  aoi22 U266 ( .Y(n173), .A0(A[51]), .A1(n174), .B0(n175), .B1(n176) );
  nand02 U267 ( .Y(n176), .A0(B[50]), .A1(n177) );
  ao221 U268 ( .Y(n179), .A0(n180), .A1(B[48]), .B0(n178), .B1(B[49]), .C0(
        n181) );
  ao221 U269 ( .Y(n184), .A0(n185), .A1(B[46]), .B0(n183), .B1(B[47]), .C0(
        n186) );
  ao221 U270 ( .Y(n189), .A0(n190), .A1(B[44]), .B0(n188), .B1(B[45]), .C0(
        n191) );
  ao221 U271 ( .Y(n194), .A0(n195), .A1(B[42]), .B0(n193), .B1(B[43]), .C0(
        n196) );
  ao221 U272 ( .Y(n199), .A0(n200), .A1(B[40]), .B0(n198), .B1(B[41]), .C0(
        n201) );
  ao221 U273 ( .Y(n204), .A0(n205), .A1(B[38]), .B0(n203), .B1(B[39]), .C0(
        n206) );
  ao221 U274 ( .Y(n209), .A0(n210), .A1(B[36]), .B0(n208), .B1(B[37]), .C0(
        n211) );
  ao221 U275 ( .Y(n214), .A0(n215), .A1(B[34]), .B0(n213), .B1(B[35]), .C0(
        n216) );
  ao221 U276 ( .Y(n219), .A0(n220), .A1(B[32]), .B0(n218), .B1(B[33]), .C0(
        n221) );
  ao221 U277 ( .Y(n224), .A0(n225), .A1(B[30]), .B0(n223), .B1(B[31]), .C0(
        n226) );
  ao221 U278 ( .Y(n229), .A0(n230), .A1(B[28]), .B0(n228), .B1(B[29]), .C0(
        n231) );
  ao221 U279 ( .Y(n234), .A0(n235), .A1(B[26]), .B0(n233), .B1(B[27]), .C0(
        n236) );
  ao221 U280 ( .Y(n239), .A0(n240), .A1(B[24]), .B0(n238), .B1(B[25]), .C0(
        n241) );
  ao221 U281 ( .Y(n244), .A0(n245), .A1(B[22]), .B0(n243), .B1(B[23]), .C0(
        n246) );
  ao221 U282 ( .Y(n249), .A0(n250), .A1(B[20]), .B0(n248), .B1(B[21]), .C0(
        n251) );
  ao221 U283 ( .Y(n254), .A0(n255), .A1(B[18]), .B0(n253), .B1(B[19]), .C0(
        n256) );
  ao221 U284 ( .Y(n259), .A0(n260), .A1(B[16]), .B0(n258), .B1(B[17]), .C0(
        n261) );
  ao221 U285 ( .Y(n264), .A0(n265), .A1(B[14]), .B0(n263), .B1(B[15]), .C0(
        n266) );
  ao221 U286 ( .Y(n269), .A0(n270), .A1(B[12]), .B0(n268), .B1(B[13]), .C0(
        n271) );
  ao221 U287 ( .Y(n274), .A0(n275), .A1(B[10]), .B0(n273), .B1(B[11]), .C0(
        n276) );
  ao221 U288 ( .Y(n279), .A0(n280), .A1(B[8]), .B0(n278), .B1(B[9]), .C0(n281)
         );
  ao221 U289 ( .Y(n284), .A0(n285), .A1(B[6]), .B0(n283), .B1(B[7]), .C0(n286)
         );
  ao221 U290 ( .Y(n289), .A0(n290), .A1(B[4]), .B0(n288), .B1(B[5]), .C0(n291)
         );
  ao221 U291 ( .Y(n294), .A0(n295), .A1(B[2]), .B0(n293), .B1(B[3]), .C0(n296)
         );
  ao21 U292 ( .Y(n300), .A0(n298), .A1(n299), .B0(B[1]) );
  nor02 U293 ( .Y(n298), .A0(n301), .A1(A[0]) );
endmodule


module sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_add_52_1 ( A, B, CI, SUM, CO );
  input [51:0] A;
  input [51:0] B;
  output [51:0] SUM;
  input CI;
  output CO;
  wire   carry_51_, carry_50_, carry_49_, carry_48_, carry_47_, carry_46_,
         carry_45_, carry_44_, carry_43_, carry_42_, carry_41_, carry_40_,
         carry_39_, carry_38_, carry_37_, carry_36_, carry_35_, carry_34_,
         carry_33_, carry_32_, carry_31_, carry_30_, carry_29_, carry_28_,
         carry_27_, carry_26_, carry_25_, carry_24_, carry_23_, carry_22_,
         carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, carry_6_, carry_5_, carry_4_, carry_3_,
         carry_2_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303;

  nand02 U4 ( .Y(n1), .A0(A[0]), .A1(B[0]) );
  inv02 U5 ( .Y(n2), .A(n1) );
  inv01 U6 ( .Y(SUM[50]), .A(n3) );
  inv02 U7 ( .Y(carry_51_), .A(n4) );
  inv02 U8 ( .Y(n5), .A(B[50]) );
  inv02 U9 ( .Y(n6), .A(A[50]) );
  inv02 U10 ( .Y(n7), .A(carry_50_) );
  nor02 U11 ( .Y(n8), .A0(n5), .A1(n9) );
  nor02 U12 ( .Y(n10), .A0(n6), .A1(n11) );
  nor02 U13 ( .Y(n12), .A0(n7), .A1(n13) );
  nor02 U14 ( .Y(n14), .A0(n7), .A1(n15) );
  nor02 U15 ( .Y(n3), .A0(n16), .A1(n17) );
  nor02 U16 ( .Y(n18), .A0(n6), .A1(n7) );
  nor02 U17 ( .Y(n19), .A0(n5), .A1(n7) );
  nor02 U18 ( .Y(n20), .A0(n5), .A1(n6) );
  nor02 U19 ( .Y(n4), .A0(n20), .A1(n21) );
  nor02 U20 ( .Y(n22), .A0(A[50]), .A1(carry_50_) );
  inv01 U21 ( .Y(n9), .A(n22) );
  nor02 U22 ( .Y(n23), .A0(B[50]), .A1(carry_50_) );
  inv01 U23 ( .Y(n11), .A(n23) );
  nor02 U24 ( .Y(n24), .A0(B[50]), .A1(A[50]) );
  inv01 U25 ( .Y(n13), .A(n24) );
  nor02 U26 ( .Y(n25), .A0(n5), .A1(n6) );
  inv01 U27 ( .Y(n15), .A(n25) );
  nor02 U28 ( .Y(n26), .A0(n8), .A1(n10) );
  inv01 U29 ( .Y(n16), .A(n26) );
  nor02 U30 ( .Y(n27), .A0(n12), .A1(n14) );
  inv01 U31 ( .Y(n17), .A(n27) );
  nor02 U32 ( .Y(n28), .A0(n18), .A1(n19) );
  inv01 U33 ( .Y(n21), .A(n28) );
  inv01 U34 ( .Y(SUM[49]), .A(n29) );
  inv02 U35 ( .Y(carry_50_), .A(n30) );
  inv02 U36 ( .Y(n31), .A(B[49]) );
  inv02 U37 ( .Y(n32), .A(A[49]) );
  inv02 U38 ( .Y(n33), .A(carry_49_) );
  nor02 U39 ( .Y(n34), .A0(n31), .A1(n35) );
  nor02 U40 ( .Y(n36), .A0(n32), .A1(n37) );
  nor02 U41 ( .Y(n38), .A0(n33), .A1(n39) );
  nor02 U42 ( .Y(n40), .A0(n33), .A1(n41) );
  nor02 U43 ( .Y(n29), .A0(n42), .A1(n43) );
  nor02 U44 ( .Y(n44), .A0(n32), .A1(n33) );
  nor02 U45 ( .Y(n45), .A0(n31), .A1(n33) );
  nor02 U46 ( .Y(n46), .A0(n31), .A1(n32) );
  nor02 U47 ( .Y(n30), .A0(n46), .A1(n47) );
  nor02 U48 ( .Y(n48), .A0(A[49]), .A1(carry_49_) );
  inv01 U49 ( .Y(n35), .A(n48) );
  nor02 U50 ( .Y(n49), .A0(B[49]), .A1(carry_49_) );
  inv01 U51 ( .Y(n37), .A(n49) );
  nor02 U52 ( .Y(n50), .A0(B[49]), .A1(A[49]) );
  inv01 U53 ( .Y(n39), .A(n50) );
  nor02 U54 ( .Y(n51), .A0(n31), .A1(n32) );
  inv01 U55 ( .Y(n41), .A(n51) );
  nor02 U56 ( .Y(n52), .A0(n34), .A1(n36) );
  inv01 U57 ( .Y(n42), .A(n52) );
  nor02 U58 ( .Y(n53), .A0(n38), .A1(n40) );
  inv01 U59 ( .Y(n43), .A(n53) );
  nor02 U60 ( .Y(n54), .A0(n44), .A1(n45) );
  inv01 U61 ( .Y(n47), .A(n54) );
  inv01 U62 ( .Y(SUM[48]), .A(n55) );
  inv02 U63 ( .Y(carry_49_), .A(n56) );
  inv02 U64 ( .Y(n57), .A(B[48]) );
  inv02 U65 ( .Y(n58), .A(A[48]) );
  inv02 U66 ( .Y(n59), .A(carry_48_) );
  nor02 U67 ( .Y(n60), .A0(n57), .A1(n61) );
  nor02 U68 ( .Y(n62), .A0(n58), .A1(n63) );
  nor02 U69 ( .Y(n64), .A0(n59), .A1(n65) );
  nor02 U70 ( .Y(n66), .A0(n59), .A1(n67) );
  nor02 U71 ( .Y(n55), .A0(n68), .A1(n69) );
  nor02 U72 ( .Y(n70), .A0(n58), .A1(n59) );
  nor02 U73 ( .Y(n71), .A0(n57), .A1(n59) );
  nor02 U74 ( .Y(n72), .A0(n57), .A1(n58) );
  nor02 U75 ( .Y(n56), .A0(n72), .A1(n73) );
  nor02 U76 ( .Y(n74), .A0(A[48]), .A1(carry_48_) );
  inv01 U77 ( .Y(n61), .A(n74) );
  nor02 U78 ( .Y(n75), .A0(B[48]), .A1(carry_48_) );
  inv01 U79 ( .Y(n63), .A(n75) );
  nor02 U80 ( .Y(n76), .A0(B[48]), .A1(A[48]) );
  inv01 U81 ( .Y(n65), .A(n76) );
  nor02 U82 ( .Y(n77), .A0(n57), .A1(n58) );
  inv01 U83 ( .Y(n67), .A(n77) );
  nor02 U84 ( .Y(n78), .A0(n60), .A1(n62) );
  inv01 U85 ( .Y(n68), .A(n78) );
  nor02 U86 ( .Y(n79), .A0(n64), .A1(n66) );
  inv01 U87 ( .Y(n69), .A(n79) );
  nor02 U88 ( .Y(n80), .A0(n70), .A1(n71) );
  inv01 U89 ( .Y(n73), .A(n80) );
  inv01 U90 ( .Y(SUM[47]), .A(n81) );
  inv02 U91 ( .Y(carry_48_), .A(n82) );
  inv02 U92 ( .Y(n83), .A(B[47]) );
  inv02 U93 ( .Y(n84), .A(A[47]) );
  inv02 U94 ( .Y(n85), .A(carry_47_) );
  nor02 U95 ( .Y(n86), .A0(n83), .A1(n87) );
  nor02 U96 ( .Y(n88), .A0(n84), .A1(n89) );
  nor02 U97 ( .Y(n90), .A0(n85), .A1(n91) );
  nor02 U98 ( .Y(n92), .A0(n85), .A1(n93) );
  nor02 U99 ( .Y(n81), .A0(n94), .A1(n95) );
  nor02 U100 ( .Y(n96), .A0(n84), .A1(n85) );
  nor02 U101 ( .Y(n97), .A0(n83), .A1(n85) );
  nor02 U102 ( .Y(n98), .A0(n83), .A1(n84) );
  nor02 U103 ( .Y(n82), .A0(n98), .A1(n99) );
  nor02 U104 ( .Y(n100), .A0(A[47]), .A1(carry_47_) );
  inv01 U105 ( .Y(n87), .A(n100) );
  nor02 U106 ( .Y(n101), .A0(B[47]), .A1(carry_47_) );
  inv01 U107 ( .Y(n89), .A(n101) );
  nor02 U108 ( .Y(n102), .A0(B[47]), .A1(A[47]) );
  inv01 U109 ( .Y(n91), .A(n102) );
  nor02 U110 ( .Y(n103), .A0(n83), .A1(n84) );
  inv01 U111 ( .Y(n93), .A(n103) );
  nor02 U112 ( .Y(n104), .A0(n86), .A1(n88) );
  inv01 U113 ( .Y(n94), .A(n104) );
  nor02 U114 ( .Y(n105), .A0(n90), .A1(n92) );
  inv01 U115 ( .Y(n95), .A(n105) );
  nor02 U116 ( .Y(n106), .A0(n96), .A1(n97) );
  inv01 U117 ( .Y(n99), .A(n106) );
  inv01 U118 ( .Y(SUM[46]), .A(n107) );
  inv02 U119 ( .Y(carry_47_), .A(n108) );
  inv02 U120 ( .Y(n109), .A(B[46]) );
  inv02 U121 ( .Y(n110), .A(A[46]) );
  inv02 U122 ( .Y(n111), .A(carry_46_) );
  nor02 U123 ( .Y(n112), .A0(n109), .A1(n113) );
  nor02 U124 ( .Y(n114), .A0(n110), .A1(n115) );
  nor02 U125 ( .Y(n116), .A0(n111), .A1(n117) );
  nor02 U126 ( .Y(n118), .A0(n111), .A1(n119) );
  nor02 U127 ( .Y(n107), .A0(n120), .A1(n121) );
  nor02 U128 ( .Y(n122), .A0(n110), .A1(n111) );
  nor02 U129 ( .Y(n123), .A0(n109), .A1(n111) );
  nor02 U130 ( .Y(n124), .A0(n109), .A1(n110) );
  nor02 U131 ( .Y(n108), .A0(n124), .A1(n125) );
  nor02 U132 ( .Y(n126), .A0(A[46]), .A1(carry_46_) );
  inv01 U133 ( .Y(n113), .A(n126) );
  nor02 U134 ( .Y(n127), .A0(B[46]), .A1(carry_46_) );
  inv01 U135 ( .Y(n115), .A(n127) );
  nor02 U136 ( .Y(n128), .A0(B[46]), .A1(A[46]) );
  inv01 U137 ( .Y(n117), .A(n128) );
  nor02 U138 ( .Y(n129), .A0(n109), .A1(n110) );
  inv01 U139 ( .Y(n119), .A(n129) );
  nor02 U140 ( .Y(n130), .A0(n112), .A1(n114) );
  inv01 U141 ( .Y(n120), .A(n130) );
  nor02 U142 ( .Y(n131), .A0(n116), .A1(n118) );
  inv01 U143 ( .Y(n121), .A(n131) );
  nor02 U144 ( .Y(n132), .A0(n122), .A1(n123) );
  inv01 U145 ( .Y(n125), .A(n132) );
  inv01 U146 ( .Y(SUM[45]), .A(n133) );
  inv02 U147 ( .Y(carry_46_), .A(n134) );
  inv02 U148 ( .Y(n135), .A(B[45]) );
  inv02 U149 ( .Y(n136), .A(A[45]) );
  inv02 U150 ( .Y(n137), .A(carry_45_) );
  nor02 U151 ( .Y(n138), .A0(n135), .A1(n139) );
  nor02 U152 ( .Y(n140), .A0(n136), .A1(n141) );
  nor02 U153 ( .Y(n142), .A0(n137), .A1(n143) );
  nor02 U154 ( .Y(n144), .A0(n137), .A1(n145) );
  nor02 U155 ( .Y(n133), .A0(n146), .A1(n147) );
  nor02 U156 ( .Y(n148), .A0(n136), .A1(n137) );
  nor02 U157 ( .Y(n149), .A0(n135), .A1(n137) );
  nor02 U158 ( .Y(n150), .A0(n135), .A1(n136) );
  nor02 U159 ( .Y(n134), .A0(n150), .A1(n151) );
  nor02 U160 ( .Y(n152), .A0(A[45]), .A1(carry_45_) );
  inv01 U161 ( .Y(n139), .A(n152) );
  nor02 U162 ( .Y(n153), .A0(B[45]), .A1(carry_45_) );
  inv01 U163 ( .Y(n141), .A(n153) );
  nor02 U164 ( .Y(n154), .A0(B[45]), .A1(A[45]) );
  inv01 U165 ( .Y(n143), .A(n154) );
  nor02 U166 ( .Y(n155), .A0(n135), .A1(n136) );
  inv01 U167 ( .Y(n145), .A(n155) );
  nor02 U168 ( .Y(n156), .A0(n138), .A1(n140) );
  inv01 U169 ( .Y(n146), .A(n156) );
  nor02 U170 ( .Y(n157), .A0(n142), .A1(n144) );
  inv01 U171 ( .Y(n147), .A(n157) );
  nor02 U172 ( .Y(n158), .A0(n148), .A1(n149) );
  inv01 U173 ( .Y(n151), .A(n158) );
  inv01 U174 ( .Y(SUM[44]), .A(n159) );
  inv02 U175 ( .Y(carry_45_), .A(n160) );
  inv02 U176 ( .Y(n161), .A(B[44]) );
  inv02 U177 ( .Y(n162), .A(A[44]) );
  inv02 U178 ( .Y(n163), .A(carry_44_) );
  nor02 U179 ( .Y(n164), .A0(n161), .A1(n165) );
  nor02 U180 ( .Y(n166), .A0(n162), .A1(n167) );
  nor02 U181 ( .Y(n168), .A0(n163), .A1(n169) );
  nor02 U182 ( .Y(n170), .A0(n163), .A1(n171) );
  nor02 U183 ( .Y(n159), .A0(n172), .A1(n173) );
  nor02 U184 ( .Y(n174), .A0(n162), .A1(n163) );
  nor02 U185 ( .Y(n175), .A0(n161), .A1(n163) );
  nor02 U186 ( .Y(n176), .A0(n161), .A1(n162) );
  nor02 U187 ( .Y(n160), .A0(n176), .A1(n177) );
  nor02 U188 ( .Y(n178), .A0(A[44]), .A1(carry_44_) );
  inv01 U189 ( .Y(n165), .A(n178) );
  nor02 U190 ( .Y(n179), .A0(B[44]), .A1(carry_44_) );
  inv01 U191 ( .Y(n167), .A(n179) );
  nor02 U192 ( .Y(n180), .A0(B[44]), .A1(A[44]) );
  inv01 U193 ( .Y(n169), .A(n180) );
  nor02 U194 ( .Y(n181), .A0(n161), .A1(n162) );
  inv01 U195 ( .Y(n171), .A(n181) );
  nor02 U196 ( .Y(n182), .A0(n164), .A1(n166) );
  inv01 U197 ( .Y(n172), .A(n182) );
  nor02 U198 ( .Y(n183), .A0(n168), .A1(n170) );
  inv01 U199 ( .Y(n173), .A(n183) );
  nor02 U200 ( .Y(n184), .A0(n174), .A1(n175) );
  inv01 U201 ( .Y(n177), .A(n184) );
  inv01 U202 ( .Y(SUM[43]), .A(n185) );
  inv02 U203 ( .Y(carry_44_), .A(n186) );
  inv02 U204 ( .Y(n187), .A(B[43]) );
  inv02 U205 ( .Y(n188), .A(A[43]) );
  inv02 U206 ( .Y(n189), .A(carry_43_) );
  nor02 U207 ( .Y(n190), .A0(n187), .A1(n191) );
  nor02 U208 ( .Y(n192), .A0(n188), .A1(n193) );
  nor02 U209 ( .Y(n194), .A0(n189), .A1(n195) );
  nor02 U210 ( .Y(n196), .A0(n189), .A1(n197) );
  nor02 U211 ( .Y(n185), .A0(n198), .A1(n199) );
  nor02 U212 ( .Y(n200), .A0(n188), .A1(n189) );
  nor02 U213 ( .Y(n201), .A0(n187), .A1(n189) );
  nor02 U214 ( .Y(n202), .A0(n187), .A1(n188) );
  nor02 U215 ( .Y(n186), .A0(n202), .A1(n203) );
  nor02 U216 ( .Y(n204), .A0(A[43]), .A1(carry_43_) );
  inv01 U217 ( .Y(n191), .A(n204) );
  nor02 U218 ( .Y(n205), .A0(B[43]), .A1(carry_43_) );
  inv01 U219 ( .Y(n193), .A(n205) );
  nor02 U220 ( .Y(n206), .A0(B[43]), .A1(A[43]) );
  inv01 U221 ( .Y(n195), .A(n206) );
  nor02 U222 ( .Y(n207), .A0(n187), .A1(n188) );
  inv01 U223 ( .Y(n197), .A(n207) );
  nor02 U224 ( .Y(n208), .A0(n190), .A1(n192) );
  inv01 U225 ( .Y(n198), .A(n208) );
  nor02 U226 ( .Y(n209), .A0(n194), .A1(n196) );
  inv01 U227 ( .Y(n199), .A(n209) );
  nor02 U228 ( .Y(n210), .A0(n200), .A1(n201) );
  inv01 U229 ( .Y(n203), .A(n210) );
  inv01 U230 ( .Y(SUM[42]), .A(n211) );
  inv02 U231 ( .Y(carry_43_), .A(n212) );
  inv02 U232 ( .Y(n213), .A(B[42]) );
  inv02 U233 ( .Y(n214), .A(A[42]) );
  inv02 U234 ( .Y(n215), .A(carry_42_) );
  nor02 U235 ( .Y(n216), .A0(n213), .A1(n217) );
  nor02 U236 ( .Y(n218), .A0(n214), .A1(n219) );
  nor02 U237 ( .Y(n220), .A0(n215), .A1(n221) );
  nor02 U238 ( .Y(n222), .A0(n215), .A1(n223) );
  nor02 U239 ( .Y(n211), .A0(n224), .A1(n225) );
  nor02 U240 ( .Y(n226), .A0(n214), .A1(n215) );
  nor02 U241 ( .Y(n227), .A0(n213), .A1(n215) );
  nor02 U242 ( .Y(n228), .A0(n213), .A1(n214) );
  nor02 U243 ( .Y(n212), .A0(n228), .A1(n229) );
  nor02 U244 ( .Y(n230), .A0(A[42]), .A1(carry_42_) );
  inv01 U245 ( .Y(n217), .A(n230) );
  nor02 U246 ( .Y(n231), .A0(B[42]), .A1(carry_42_) );
  inv01 U247 ( .Y(n219), .A(n231) );
  nor02 U248 ( .Y(n232), .A0(B[42]), .A1(A[42]) );
  inv01 U249 ( .Y(n221), .A(n232) );
  nor02 U250 ( .Y(n233), .A0(n213), .A1(n214) );
  inv01 U251 ( .Y(n223), .A(n233) );
  nor02 U252 ( .Y(n234), .A0(n216), .A1(n218) );
  inv01 U253 ( .Y(n224), .A(n234) );
  nor02 U254 ( .Y(n235), .A0(n220), .A1(n222) );
  inv01 U255 ( .Y(n225), .A(n235) );
  nor02 U256 ( .Y(n236), .A0(n226), .A1(n227) );
  inv01 U257 ( .Y(n229), .A(n236) );
  inv01 U258 ( .Y(SUM[41]), .A(n237) );
  inv02 U259 ( .Y(carry_42_), .A(n238) );
  inv02 U260 ( .Y(n239), .A(B[41]) );
  inv02 U261 ( .Y(n240), .A(A[41]) );
  inv02 U262 ( .Y(n241), .A(carry_41_) );
  nor02 U263 ( .Y(n242), .A0(n239), .A1(n243) );
  nor02 U264 ( .Y(n244), .A0(n240), .A1(n245) );
  nor02 U265 ( .Y(n246), .A0(n241), .A1(n247) );
  nor02 U266 ( .Y(n248), .A0(n241), .A1(n249) );
  nor02 U267 ( .Y(n237), .A0(n250), .A1(n251) );
  nor02 U268 ( .Y(n252), .A0(n240), .A1(n241) );
  nor02 U269 ( .Y(n253), .A0(n239), .A1(n241) );
  nor02 U270 ( .Y(n254), .A0(n239), .A1(n240) );
  nor02 U271 ( .Y(n238), .A0(n254), .A1(n255) );
  nor02 U272 ( .Y(n256), .A0(A[41]), .A1(carry_41_) );
  inv01 U273 ( .Y(n243), .A(n256) );
  nor02 U274 ( .Y(n257), .A0(B[41]), .A1(carry_41_) );
  inv01 U275 ( .Y(n245), .A(n257) );
  nor02 U276 ( .Y(n258), .A0(B[41]), .A1(A[41]) );
  inv01 U277 ( .Y(n247), .A(n258) );
  nor02 U278 ( .Y(n259), .A0(n239), .A1(n240) );
  inv01 U279 ( .Y(n249), .A(n259) );
  nor02 U280 ( .Y(n260), .A0(n242), .A1(n244) );
  inv01 U281 ( .Y(n250), .A(n260) );
  nor02 U282 ( .Y(n261), .A0(n246), .A1(n248) );
  inv01 U283 ( .Y(n251), .A(n261) );
  nor02 U284 ( .Y(n262), .A0(n252), .A1(n253) );
  inv01 U285 ( .Y(n255), .A(n262) );
  inv01 U286 ( .Y(SUM[40]), .A(n263) );
  inv02 U287 ( .Y(carry_41_), .A(n264) );
  inv02 U288 ( .Y(n265), .A(B[40]) );
  inv02 U289 ( .Y(n266), .A(A[40]) );
  inv02 U290 ( .Y(n267), .A(carry_40_) );
  nor02 U291 ( .Y(n268), .A0(n265), .A1(n269) );
  nor02 U292 ( .Y(n270), .A0(n266), .A1(n271) );
  nor02 U293 ( .Y(n272), .A0(n267), .A1(n273) );
  nor02 U294 ( .Y(n274), .A0(n267), .A1(n275) );
  nor02 U295 ( .Y(n263), .A0(n276), .A1(n277) );
  nor02 U296 ( .Y(n278), .A0(n266), .A1(n267) );
  nor02 U297 ( .Y(n279), .A0(n265), .A1(n267) );
  nor02 U298 ( .Y(n280), .A0(n265), .A1(n266) );
  nor02 U299 ( .Y(n264), .A0(n280), .A1(n281) );
  nor02 U300 ( .Y(n282), .A0(A[40]), .A1(carry_40_) );
  inv01 U301 ( .Y(n269), .A(n282) );
  nor02 U302 ( .Y(n283), .A0(B[40]), .A1(carry_40_) );
  inv01 U303 ( .Y(n271), .A(n283) );
  nor02 U304 ( .Y(n284), .A0(B[40]), .A1(A[40]) );
  inv01 U305 ( .Y(n273), .A(n284) );
  nor02 U306 ( .Y(n285), .A0(n265), .A1(n266) );
  inv01 U307 ( .Y(n275), .A(n285) );
  nor02 U308 ( .Y(n286), .A0(n268), .A1(n270) );
  inv01 U309 ( .Y(n276), .A(n286) );
  nor02 U310 ( .Y(n287), .A0(n272), .A1(n274) );
  inv01 U311 ( .Y(n277), .A(n287) );
  nor02 U312 ( .Y(n288), .A0(n278), .A1(n279) );
  inv01 U313 ( .Y(n281), .A(n288) );
  inv01 U314 ( .Y(SUM[39]), .A(n289) );
  inv02 U315 ( .Y(carry_40_), .A(n290) );
  inv02 U316 ( .Y(n291), .A(B[39]) );
  inv02 U317 ( .Y(n292), .A(A[39]) );
  inv02 U318 ( .Y(n293), .A(carry_39_) );
  nor02 U319 ( .Y(n294), .A0(n291), .A1(n295) );
  nor02 U320 ( .Y(n296), .A0(n292), .A1(n297) );
  nor02 U321 ( .Y(n298), .A0(n293), .A1(n299) );
  nor02 U322 ( .Y(n300), .A0(n293), .A1(n301) );
  nor02 U323 ( .Y(n289), .A0(n302), .A1(n303) );
  nor02 U324 ( .Y(n304), .A0(n292), .A1(n293) );
  nor02 U325 ( .Y(n305), .A0(n291), .A1(n293) );
  nor02 U326 ( .Y(n306), .A0(n291), .A1(n292) );
  nor02 U327 ( .Y(n290), .A0(n306), .A1(n307) );
  nor02 U328 ( .Y(n308), .A0(A[39]), .A1(carry_39_) );
  inv01 U329 ( .Y(n295), .A(n308) );
  nor02 U330 ( .Y(n309), .A0(B[39]), .A1(carry_39_) );
  inv01 U331 ( .Y(n297), .A(n309) );
  nor02 U332 ( .Y(n310), .A0(B[39]), .A1(A[39]) );
  inv01 U333 ( .Y(n299), .A(n310) );
  nor02 U334 ( .Y(n311), .A0(n291), .A1(n292) );
  inv01 U335 ( .Y(n301), .A(n311) );
  nor02 U336 ( .Y(n312), .A0(n294), .A1(n296) );
  inv01 U337 ( .Y(n302), .A(n312) );
  nor02 U338 ( .Y(n313), .A0(n298), .A1(n300) );
  inv01 U339 ( .Y(n303), .A(n313) );
  nor02 U340 ( .Y(n314), .A0(n304), .A1(n305) );
  inv01 U341 ( .Y(n307), .A(n314) );
  inv01 U342 ( .Y(SUM[38]), .A(n315) );
  inv02 U343 ( .Y(carry_39_), .A(n316) );
  inv02 U344 ( .Y(n317), .A(B[38]) );
  inv02 U345 ( .Y(n318), .A(A[38]) );
  inv02 U346 ( .Y(n319), .A(carry_38_) );
  nor02 U347 ( .Y(n320), .A0(n317), .A1(n321) );
  nor02 U348 ( .Y(n322), .A0(n318), .A1(n323) );
  nor02 U349 ( .Y(n324), .A0(n319), .A1(n325) );
  nor02 U350 ( .Y(n326), .A0(n319), .A1(n327) );
  nor02 U351 ( .Y(n315), .A0(n328), .A1(n329) );
  nor02 U352 ( .Y(n330), .A0(n318), .A1(n319) );
  nor02 U353 ( .Y(n331), .A0(n317), .A1(n319) );
  nor02 U354 ( .Y(n332), .A0(n317), .A1(n318) );
  nor02 U355 ( .Y(n316), .A0(n332), .A1(n333) );
  nor02 U356 ( .Y(n334), .A0(A[38]), .A1(carry_38_) );
  inv01 U357 ( .Y(n321), .A(n334) );
  nor02 U358 ( .Y(n335), .A0(B[38]), .A1(carry_38_) );
  inv01 U359 ( .Y(n323), .A(n335) );
  nor02 U360 ( .Y(n336), .A0(B[38]), .A1(A[38]) );
  inv01 U361 ( .Y(n325), .A(n336) );
  nor02 U362 ( .Y(n337), .A0(n317), .A1(n318) );
  inv01 U363 ( .Y(n327), .A(n337) );
  nor02 U364 ( .Y(n338), .A0(n320), .A1(n322) );
  inv01 U365 ( .Y(n328), .A(n338) );
  nor02 U366 ( .Y(n339), .A0(n324), .A1(n326) );
  inv01 U367 ( .Y(n329), .A(n339) );
  nor02 U368 ( .Y(n340), .A0(n330), .A1(n331) );
  inv01 U369 ( .Y(n333), .A(n340) );
  inv01 U370 ( .Y(SUM[37]), .A(n341) );
  inv02 U371 ( .Y(carry_38_), .A(n342) );
  inv02 U372 ( .Y(n343), .A(B[37]) );
  inv02 U373 ( .Y(n344), .A(A[37]) );
  inv02 U374 ( .Y(n345), .A(carry_37_) );
  nor02 U375 ( .Y(n346), .A0(n343), .A1(n347) );
  nor02 U376 ( .Y(n348), .A0(n344), .A1(n349) );
  nor02 U377 ( .Y(n350), .A0(n345), .A1(n351) );
  nor02 U378 ( .Y(n352), .A0(n345), .A1(n353) );
  nor02 U379 ( .Y(n341), .A0(n354), .A1(n355) );
  nor02 U380 ( .Y(n356), .A0(n344), .A1(n345) );
  nor02 U381 ( .Y(n357), .A0(n343), .A1(n345) );
  nor02 U382 ( .Y(n358), .A0(n343), .A1(n344) );
  nor02 U383 ( .Y(n342), .A0(n358), .A1(n359) );
  nor02 U384 ( .Y(n360), .A0(A[37]), .A1(carry_37_) );
  inv01 U385 ( .Y(n347), .A(n360) );
  nor02 U386 ( .Y(n361), .A0(B[37]), .A1(carry_37_) );
  inv01 U387 ( .Y(n349), .A(n361) );
  nor02 U388 ( .Y(n362), .A0(B[37]), .A1(A[37]) );
  inv01 U389 ( .Y(n351), .A(n362) );
  nor02 U390 ( .Y(n363), .A0(n343), .A1(n344) );
  inv01 U391 ( .Y(n353), .A(n363) );
  nor02 U392 ( .Y(n364), .A0(n346), .A1(n348) );
  inv01 U393 ( .Y(n354), .A(n364) );
  nor02 U394 ( .Y(n365), .A0(n350), .A1(n352) );
  inv01 U395 ( .Y(n355), .A(n365) );
  nor02 U396 ( .Y(n366), .A0(n356), .A1(n357) );
  inv01 U397 ( .Y(n359), .A(n366) );
  inv01 U398 ( .Y(SUM[36]), .A(n367) );
  inv02 U399 ( .Y(carry_37_), .A(n368) );
  inv02 U400 ( .Y(n369), .A(B[36]) );
  inv02 U401 ( .Y(n370), .A(A[36]) );
  inv02 U402 ( .Y(n371), .A(carry_36_) );
  nor02 U403 ( .Y(n372), .A0(n369), .A1(n373) );
  nor02 U404 ( .Y(n374), .A0(n370), .A1(n375) );
  nor02 U405 ( .Y(n376), .A0(n371), .A1(n377) );
  nor02 U406 ( .Y(n378), .A0(n371), .A1(n379) );
  nor02 U407 ( .Y(n367), .A0(n380), .A1(n381) );
  nor02 U408 ( .Y(n382), .A0(n370), .A1(n371) );
  nor02 U409 ( .Y(n383), .A0(n369), .A1(n371) );
  nor02 U410 ( .Y(n384), .A0(n369), .A1(n370) );
  nor02 U411 ( .Y(n368), .A0(n384), .A1(n385) );
  nor02 U412 ( .Y(n386), .A0(A[36]), .A1(carry_36_) );
  inv01 U413 ( .Y(n373), .A(n386) );
  nor02 U414 ( .Y(n387), .A0(B[36]), .A1(carry_36_) );
  inv01 U415 ( .Y(n375), .A(n387) );
  nor02 U416 ( .Y(n388), .A0(B[36]), .A1(A[36]) );
  inv01 U417 ( .Y(n377), .A(n388) );
  nor02 U418 ( .Y(n389), .A0(n369), .A1(n370) );
  inv01 U419 ( .Y(n379), .A(n389) );
  nor02 U420 ( .Y(n390), .A0(n372), .A1(n374) );
  inv01 U421 ( .Y(n380), .A(n390) );
  nor02 U422 ( .Y(n391), .A0(n376), .A1(n378) );
  inv01 U423 ( .Y(n381), .A(n391) );
  nor02 U424 ( .Y(n392), .A0(n382), .A1(n383) );
  inv01 U425 ( .Y(n385), .A(n392) );
  inv01 U426 ( .Y(SUM[35]), .A(n393) );
  inv02 U427 ( .Y(carry_36_), .A(n394) );
  inv02 U428 ( .Y(n395), .A(B[35]) );
  inv02 U429 ( .Y(n396), .A(A[35]) );
  inv02 U430 ( .Y(n397), .A(carry_35_) );
  nor02 U431 ( .Y(n398), .A0(n395), .A1(n399) );
  nor02 U432 ( .Y(n400), .A0(n396), .A1(n401) );
  nor02 U433 ( .Y(n402), .A0(n397), .A1(n403) );
  nor02 U434 ( .Y(n404), .A0(n397), .A1(n405) );
  nor02 U435 ( .Y(n393), .A0(n406), .A1(n407) );
  nor02 U436 ( .Y(n408), .A0(n396), .A1(n397) );
  nor02 U437 ( .Y(n409), .A0(n395), .A1(n397) );
  nor02 U438 ( .Y(n410), .A0(n395), .A1(n396) );
  nor02 U439 ( .Y(n394), .A0(n410), .A1(n411) );
  nor02 U440 ( .Y(n412), .A0(A[35]), .A1(carry_35_) );
  inv01 U441 ( .Y(n399), .A(n412) );
  nor02 U442 ( .Y(n413), .A0(B[35]), .A1(carry_35_) );
  inv01 U443 ( .Y(n401), .A(n413) );
  nor02 U444 ( .Y(n414), .A0(B[35]), .A1(A[35]) );
  inv01 U445 ( .Y(n403), .A(n414) );
  nor02 U446 ( .Y(n415), .A0(n395), .A1(n396) );
  inv01 U447 ( .Y(n405), .A(n415) );
  nor02 U448 ( .Y(n416), .A0(n398), .A1(n400) );
  inv01 U449 ( .Y(n406), .A(n416) );
  nor02 U450 ( .Y(n417), .A0(n402), .A1(n404) );
  inv01 U451 ( .Y(n407), .A(n417) );
  nor02 U452 ( .Y(n418), .A0(n408), .A1(n409) );
  inv01 U453 ( .Y(n411), .A(n418) );
  inv01 U454 ( .Y(SUM[34]), .A(n419) );
  inv02 U455 ( .Y(carry_35_), .A(n420) );
  inv02 U456 ( .Y(n421), .A(B[34]) );
  inv02 U457 ( .Y(n422), .A(A[34]) );
  inv02 U458 ( .Y(n423), .A(carry_34_) );
  nor02 U459 ( .Y(n424), .A0(n421), .A1(n425) );
  nor02 U460 ( .Y(n426), .A0(n422), .A1(n427) );
  nor02 U461 ( .Y(n428), .A0(n423), .A1(n429) );
  nor02 U462 ( .Y(n430), .A0(n423), .A1(n431) );
  nor02 U463 ( .Y(n419), .A0(n432), .A1(n433) );
  nor02 U464 ( .Y(n434), .A0(n422), .A1(n423) );
  nor02 U465 ( .Y(n435), .A0(n421), .A1(n423) );
  nor02 U466 ( .Y(n436), .A0(n421), .A1(n422) );
  nor02 U467 ( .Y(n420), .A0(n436), .A1(n437) );
  nor02 U468 ( .Y(n438), .A0(A[34]), .A1(carry_34_) );
  inv01 U469 ( .Y(n425), .A(n438) );
  nor02 U470 ( .Y(n439), .A0(B[34]), .A1(carry_34_) );
  inv01 U471 ( .Y(n427), .A(n439) );
  nor02 U472 ( .Y(n440), .A0(B[34]), .A1(A[34]) );
  inv01 U473 ( .Y(n429), .A(n440) );
  nor02 U474 ( .Y(n441), .A0(n421), .A1(n422) );
  inv01 U475 ( .Y(n431), .A(n441) );
  nor02 U476 ( .Y(n442), .A0(n424), .A1(n426) );
  inv01 U477 ( .Y(n432), .A(n442) );
  nor02 U478 ( .Y(n443), .A0(n428), .A1(n430) );
  inv01 U479 ( .Y(n433), .A(n443) );
  nor02 U480 ( .Y(n444), .A0(n434), .A1(n435) );
  inv01 U481 ( .Y(n437), .A(n444) );
  inv01 U482 ( .Y(SUM[33]), .A(n445) );
  inv02 U483 ( .Y(carry_34_), .A(n446) );
  inv02 U484 ( .Y(n447), .A(B[33]) );
  inv02 U485 ( .Y(n448), .A(A[33]) );
  inv02 U486 ( .Y(n449), .A(carry_33_) );
  nor02 U487 ( .Y(n450), .A0(n447), .A1(n451) );
  nor02 U488 ( .Y(n452), .A0(n448), .A1(n453) );
  nor02 U489 ( .Y(n454), .A0(n449), .A1(n455) );
  nor02 U490 ( .Y(n456), .A0(n449), .A1(n457) );
  nor02 U491 ( .Y(n445), .A0(n458), .A1(n459) );
  nor02 U492 ( .Y(n460), .A0(n448), .A1(n449) );
  nor02 U493 ( .Y(n461), .A0(n447), .A1(n449) );
  nor02 U494 ( .Y(n462), .A0(n447), .A1(n448) );
  nor02 U495 ( .Y(n446), .A0(n462), .A1(n463) );
  nor02 U496 ( .Y(n464), .A0(A[33]), .A1(carry_33_) );
  inv01 U497 ( .Y(n451), .A(n464) );
  nor02 U498 ( .Y(n465), .A0(B[33]), .A1(carry_33_) );
  inv01 U499 ( .Y(n453), .A(n465) );
  nor02 U500 ( .Y(n466), .A0(B[33]), .A1(A[33]) );
  inv01 U501 ( .Y(n455), .A(n466) );
  nor02 U502 ( .Y(n467), .A0(n447), .A1(n448) );
  inv01 U503 ( .Y(n457), .A(n467) );
  nor02 U504 ( .Y(n468), .A0(n450), .A1(n452) );
  inv01 U505 ( .Y(n458), .A(n468) );
  nor02 U506 ( .Y(n469), .A0(n454), .A1(n456) );
  inv01 U507 ( .Y(n459), .A(n469) );
  nor02 U508 ( .Y(n470), .A0(n460), .A1(n461) );
  inv01 U509 ( .Y(n463), .A(n470) );
  inv01 U510 ( .Y(SUM[32]), .A(n471) );
  inv02 U511 ( .Y(carry_33_), .A(n472) );
  inv02 U512 ( .Y(n473), .A(B[32]) );
  inv02 U513 ( .Y(n474), .A(A[32]) );
  inv02 U514 ( .Y(n475), .A(carry_32_) );
  nor02 U515 ( .Y(n476), .A0(n473), .A1(n477) );
  nor02 U516 ( .Y(n478), .A0(n474), .A1(n479) );
  nor02 U517 ( .Y(n480), .A0(n475), .A1(n481) );
  nor02 U518 ( .Y(n482), .A0(n475), .A1(n483) );
  nor02 U519 ( .Y(n471), .A0(n484), .A1(n485) );
  nor02 U520 ( .Y(n486), .A0(n474), .A1(n475) );
  nor02 U521 ( .Y(n487), .A0(n473), .A1(n475) );
  nor02 U522 ( .Y(n488), .A0(n473), .A1(n474) );
  nor02 U523 ( .Y(n472), .A0(n488), .A1(n489) );
  nor02 U524 ( .Y(n490), .A0(A[32]), .A1(carry_32_) );
  inv01 U525 ( .Y(n477), .A(n490) );
  nor02 U526 ( .Y(n491), .A0(B[32]), .A1(carry_32_) );
  inv01 U527 ( .Y(n479), .A(n491) );
  nor02 U528 ( .Y(n492), .A0(B[32]), .A1(A[32]) );
  inv01 U529 ( .Y(n481), .A(n492) );
  nor02 U530 ( .Y(n493), .A0(n473), .A1(n474) );
  inv01 U531 ( .Y(n483), .A(n493) );
  nor02 U532 ( .Y(n494), .A0(n476), .A1(n478) );
  inv01 U533 ( .Y(n484), .A(n494) );
  nor02 U534 ( .Y(n495), .A0(n480), .A1(n482) );
  inv01 U535 ( .Y(n485), .A(n495) );
  nor02 U536 ( .Y(n496), .A0(n486), .A1(n487) );
  inv01 U537 ( .Y(n489), .A(n496) );
  inv01 U538 ( .Y(SUM[31]), .A(n497) );
  inv02 U539 ( .Y(carry_32_), .A(n498) );
  inv02 U540 ( .Y(n499), .A(B[31]) );
  inv02 U541 ( .Y(n500), .A(A[31]) );
  inv02 U542 ( .Y(n501), .A(carry_31_) );
  nor02 U543 ( .Y(n502), .A0(n499), .A1(n503) );
  nor02 U544 ( .Y(n504), .A0(n500), .A1(n505) );
  nor02 U545 ( .Y(n506), .A0(n501), .A1(n507) );
  nor02 U546 ( .Y(n508), .A0(n501), .A1(n509) );
  nor02 U547 ( .Y(n497), .A0(n510), .A1(n511) );
  nor02 U548 ( .Y(n512), .A0(n500), .A1(n501) );
  nor02 U549 ( .Y(n513), .A0(n499), .A1(n501) );
  nor02 U550 ( .Y(n514), .A0(n499), .A1(n500) );
  nor02 U551 ( .Y(n498), .A0(n514), .A1(n515) );
  nor02 U552 ( .Y(n516), .A0(A[31]), .A1(carry_31_) );
  inv01 U553 ( .Y(n503), .A(n516) );
  nor02 U554 ( .Y(n517), .A0(B[31]), .A1(carry_31_) );
  inv01 U555 ( .Y(n505), .A(n517) );
  nor02 U556 ( .Y(n518), .A0(B[31]), .A1(A[31]) );
  inv01 U557 ( .Y(n507), .A(n518) );
  nor02 U558 ( .Y(n519), .A0(n499), .A1(n500) );
  inv01 U559 ( .Y(n509), .A(n519) );
  nor02 U560 ( .Y(n520), .A0(n502), .A1(n504) );
  inv01 U561 ( .Y(n510), .A(n520) );
  nor02 U562 ( .Y(n521), .A0(n506), .A1(n508) );
  inv01 U563 ( .Y(n511), .A(n521) );
  nor02 U564 ( .Y(n522), .A0(n512), .A1(n513) );
  inv01 U565 ( .Y(n515), .A(n522) );
  inv01 U566 ( .Y(SUM[30]), .A(n523) );
  inv02 U567 ( .Y(carry_31_), .A(n524) );
  inv02 U568 ( .Y(n525), .A(B[30]) );
  inv02 U569 ( .Y(n526), .A(A[30]) );
  inv02 U570 ( .Y(n527), .A(carry_30_) );
  nor02 U571 ( .Y(n528), .A0(n525), .A1(n529) );
  nor02 U572 ( .Y(n530), .A0(n526), .A1(n531) );
  nor02 U573 ( .Y(n532), .A0(n527), .A1(n533) );
  nor02 U574 ( .Y(n534), .A0(n527), .A1(n535) );
  nor02 U575 ( .Y(n523), .A0(n536), .A1(n537) );
  nor02 U576 ( .Y(n538), .A0(n526), .A1(n527) );
  nor02 U577 ( .Y(n539), .A0(n525), .A1(n527) );
  nor02 U578 ( .Y(n540), .A0(n525), .A1(n526) );
  nor02 U579 ( .Y(n524), .A0(n540), .A1(n541) );
  nor02 U580 ( .Y(n542), .A0(A[30]), .A1(carry_30_) );
  inv01 U581 ( .Y(n529), .A(n542) );
  nor02 U582 ( .Y(n543), .A0(B[30]), .A1(carry_30_) );
  inv01 U583 ( .Y(n531), .A(n543) );
  nor02 U584 ( .Y(n544), .A0(B[30]), .A1(A[30]) );
  inv01 U585 ( .Y(n533), .A(n544) );
  nor02 U586 ( .Y(n545), .A0(n525), .A1(n526) );
  inv01 U587 ( .Y(n535), .A(n545) );
  nor02 U588 ( .Y(n546), .A0(n528), .A1(n530) );
  inv01 U589 ( .Y(n536), .A(n546) );
  nor02 U590 ( .Y(n547), .A0(n532), .A1(n534) );
  inv01 U591 ( .Y(n537), .A(n547) );
  nor02 U592 ( .Y(n548), .A0(n538), .A1(n539) );
  inv01 U593 ( .Y(n541), .A(n548) );
  inv01 U594 ( .Y(SUM[29]), .A(n549) );
  inv02 U595 ( .Y(carry_30_), .A(n550) );
  inv02 U596 ( .Y(n551), .A(B[29]) );
  inv02 U597 ( .Y(n552), .A(A[29]) );
  inv02 U598 ( .Y(n553), .A(carry_29_) );
  nor02 U599 ( .Y(n554), .A0(n551), .A1(n555) );
  nor02 U600 ( .Y(n556), .A0(n552), .A1(n557) );
  nor02 U601 ( .Y(n558), .A0(n553), .A1(n559) );
  nor02 U602 ( .Y(n560), .A0(n553), .A1(n561) );
  nor02 U603 ( .Y(n549), .A0(n562), .A1(n563) );
  nor02 U604 ( .Y(n564), .A0(n552), .A1(n553) );
  nor02 U605 ( .Y(n565), .A0(n551), .A1(n553) );
  nor02 U606 ( .Y(n566), .A0(n551), .A1(n552) );
  nor02 U607 ( .Y(n550), .A0(n566), .A1(n567) );
  nor02 U608 ( .Y(n568), .A0(A[29]), .A1(carry_29_) );
  inv01 U609 ( .Y(n555), .A(n568) );
  nor02 U610 ( .Y(n569), .A0(B[29]), .A1(carry_29_) );
  inv01 U611 ( .Y(n557), .A(n569) );
  nor02 U612 ( .Y(n570), .A0(B[29]), .A1(A[29]) );
  inv01 U613 ( .Y(n559), .A(n570) );
  nor02 U614 ( .Y(n571), .A0(n551), .A1(n552) );
  inv01 U615 ( .Y(n561), .A(n571) );
  nor02 U616 ( .Y(n572), .A0(n554), .A1(n556) );
  inv01 U617 ( .Y(n562), .A(n572) );
  nor02 U618 ( .Y(n573), .A0(n558), .A1(n560) );
  inv01 U619 ( .Y(n563), .A(n573) );
  nor02 U620 ( .Y(n574), .A0(n564), .A1(n565) );
  inv01 U621 ( .Y(n567), .A(n574) );
  inv01 U622 ( .Y(SUM[28]), .A(n575) );
  inv02 U623 ( .Y(carry_29_), .A(n576) );
  inv02 U624 ( .Y(n577), .A(B[28]) );
  inv02 U625 ( .Y(n578), .A(A[28]) );
  inv02 U626 ( .Y(n579), .A(carry_28_) );
  nor02 U627 ( .Y(n580), .A0(n577), .A1(n581) );
  nor02 U628 ( .Y(n582), .A0(n578), .A1(n583) );
  nor02 U629 ( .Y(n584), .A0(n579), .A1(n585) );
  nor02 U630 ( .Y(n586), .A0(n579), .A1(n587) );
  nor02 U631 ( .Y(n575), .A0(n588), .A1(n589) );
  nor02 U632 ( .Y(n590), .A0(n578), .A1(n579) );
  nor02 U633 ( .Y(n591), .A0(n577), .A1(n579) );
  nor02 U634 ( .Y(n592), .A0(n577), .A1(n578) );
  nor02 U635 ( .Y(n576), .A0(n592), .A1(n593) );
  nor02 U636 ( .Y(n594), .A0(A[28]), .A1(carry_28_) );
  inv01 U637 ( .Y(n581), .A(n594) );
  nor02 U638 ( .Y(n595), .A0(B[28]), .A1(carry_28_) );
  inv01 U639 ( .Y(n583), .A(n595) );
  nor02 U640 ( .Y(n596), .A0(B[28]), .A1(A[28]) );
  inv01 U641 ( .Y(n585), .A(n596) );
  nor02 U642 ( .Y(n597), .A0(n577), .A1(n578) );
  inv01 U643 ( .Y(n587), .A(n597) );
  nor02 U644 ( .Y(n598), .A0(n580), .A1(n582) );
  inv01 U645 ( .Y(n588), .A(n598) );
  nor02 U646 ( .Y(n599), .A0(n584), .A1(n586) );
  inv01 U647 ( .Y(n589), .A(n599) );
  nor02 U648 ( .Y(n600), .A0(n590), .A1(n591) );
  inv01 U649 ( .Y(n593), .A(n600) );
  inv01 U650 ( .Y(SUM[27]), .A(n601) );
  inv02 U651 ( .Y(carry_28_), .A(n602) );
  inv02 U652 ( .Y(n603), .A(B[27]) );
  inv02 U653 ( .Y(n604), .A(A[27]) );
  inv02 U654 ( .Y(n605), .A(carry_27_) );
  nor02 U655 ( .Y(n606), .A0(n603), .A1(n607) );
  nor02 U656 ( .Y(n608), .A0(n604), .A1(n609) );
  nor02 U657 ( .Y(n610), .A0(n605), .A1(n611) );
  nor02 U658 ( .Y(n612), .A0(n605), .A1(n613) );
  nor02 U659 ( .Y(n601), .A0(n614), .A1(n615) );
  nor02 U660 ( .Y(n616), .A0(n604), .A1(n605) );
  nor02 U661 ( .Y(n617), .A0(n603), .A1(n605) );
  nor02 U662 ( .Y(n618), .A0(n603), .A1(n604) );
  nor02 U663 ( .Y(n602), .A0(n618), .A1(n619) );
  nor02 U664 ( .Y(n620), .A0(A[27]), .A1(carry_27_) );
  inv01 U665 ( .Y(n607), .A(n620) );
  nor02 U666 ( .Y(n621), .A0(B[27]), .A1(carry_27_) );
  inv01 U667 ( .Y(n609), .A(n621) );
  nor02 U668 ( .Y(n622), .A0(B[27]), .A1(A[27]) );
  inv01 U669 ( .Y(n611), .A(n622) );
  nor02 U670 ( .Y(n623), .A0(n603), .A1(n604) );
  inv01 U671 ( .Y(n613), .A(n623) );
  nor02 U672 ( .Y(n624), .A0(n606), .A1(n608) );
  inv01 U673 ( .Y(n614), .A(n624) );
  nor02 U674 ( .Y(n625), .A0(n610), .A1(n612) );
  inv01 U675 ( .Y(n615), .A(n625) );
  nor02 U676 ( .Y(n626), .A0(n616), .A1(n617) );
  inv01 U677 ( .Y(n619), .A(n626) );
  inv01 U678 ( .Y(SUM[26]), .A(n627) );
  inv02 U679 ( .Y(carry_27_), .A(n628) );
  inv02 U680 ( .Y(n629), .A(B[26]) );
  inv02 U681 ( .Y(n630), .A(A[26]) );
  inv02 U682 ( .Y(n631), .A(carry_26_) );
  nor02 U683 ( .Y(n632), .A0(n629), .A1(n633) );
  nor02 U684 ( .Y(n634), .A0(n630), .A1(n635) );
  nor02 U685 ( .Y(n636), .A0(n631), .A1(n637) );
  nor02 U686 ( .Y(n638), .A0(n631), .A1(n639) );
  nor02 U687 ( .Y(n627), .A0(n640), .A1(n641) );
  nor02 U688 ( .Y(n642), .A0(n630), .A1(n631) );
  nor02 U689 ( .Y(n643), .A0(n629), .A1(n631) );
  nor02 U690 ( .Y(n644), .A0(n629), .A1(n630) );
  nor02 U691 ( .Y(n628), .A0(n644), .A1(n645) );
  nor02 U692 ( .Y(n646), .A0(A[26]), .A1(carry_26_) );
  inv01 U693 ( .Y(n633), .A(n646) );
  nor02 U694 ( .Y(n647), .A0(B[26]), .A1(carry_26_) );
  inv01 U695 ( .Y(n635), .A(n647) );
  nor02 U696 ( .Y(n648), .A0(B[26]), .A1(A[26]) );
  inv01 U697 ( .Y(n637), .A(n648) );
  nor02 U698 ( .Y(n649), .A0(n629), .A1(n630) );
  inv01 U699 ( .Y(n639), .A(n649) );
  nor02 U700 ( .Y(n650), .A0(n632), .A1(n634) );
  inv01 U701 ( .Y(n640), .A(n650) );
  nor02 U702 ( .Y(n651), .A0(n636), .A1(n638) );
  inv01 U703 ( .Y(n641), .A(n651) );
  nor02 U704 ( .Y(n652), .A0(n642), .A1(n643) );
  inv01 U705 ( .Y(n645), .A(n652) );
  inv01 U706 ( .Y(SUM[25]), .A(n653) );
  inv02 U707 ( .Y(carry_26_), .A(n654) );
  inv02 U708 ( .Y(n655), .A(B[25]) );
  inv02 U709 ( .Y(n656), .A(A[25]) );
  inv02 U710 ( .Y(n657), .A(carry_25_) );
  nor02 U711 ( .Y(n658), .A0(n655), .A1(n659) );
  nor02 U712 ( .Y(n660), .A0(n656), .A1(n661) );
  nor02 U713 ( .Y(n662), .A0(n657), .A1(n663) );
  nor02 U714 ( .Y(n664), .A0(n657), .A1(n665) );
  nor02 U715 ( .Y(n653), .A0(n666), .A1(n667) );
  nor02 U716 ( .Y(n668), .A0(n656), .A1(n657) );
  nor02 U717 ( .Y(n669), .A0(n655), .A1(n657) );
  nor02 U718 ( .Y(n670), .A0(n655), .A1(n656) );
  nor02 U719 ( .Y(n654), .A0(n670), .A1(n671) );
  nor02 U720 ( .Y(n672), .A0(A[25]), .A1(carry_25_) );
  inv01 U721 ( .Y(n659), .A(n672) );
  nor02 U722 ( .Y(n673), .A0(B[25]), .A1(carry_25_) );
  inv01 U723 ( .Y(n661), .A(n673) );
  nor02 U724 ( .Y(n674), .A0(B[25]), .A1(A[25]) );
  inv01 U725 ( .Y(n663), .A(n674) );
  nor02 U726 ( .Y(n675), .A0(n655), .A1(n656) );
  inv01 U727 ( .Y(n665), .A(n675) );
  nor02 U728 ( .Y(n676), .A0(n658), .A1(n660) );
  inv01 U729 ( .Y(n666), .A(n676) );
  nor02 U730 ( .Y(n677), .A0(n662), .A1(n664) );
  inv01 U731 ( .Y(n667), .A(n677) );
  nor02 U732 ( .Y(n678), .A0(n668), .A1(n669) );
  inv01 U733 ( .Y(n671), .A(n678) );
  inv01 U734 ( .Y(SUM[24]), .A(n679) );
  inv02 U735 ( .Y(carry_25_), .A(n680) );
  inv02 U736 ( .Y(n681), .A(B[24]) );
  inv02 U737 ( .Y(n682), .A(A[24]) );
  inv02 U738 ( .Y(n683), .A(carry_24_) );
  nor02 U739 ( .Y(n684), .A0(n681), .A1(n685) );
  nor02 U740 ( .Y(n686), .A0(n682), .A1(n687) );
  nor02 U741 ( .Y(n688), .A0(n683), .A1(n689) );
  nor02 U742 ( .Y(n690), .A0(n683), .A1(n691) );
  nor02 U743 ( .Y(n679), .A0(n692), .A1(n693) );
  nor02 U744 ( .Y(n694), .A0(n682), .A1(n683) );
  nor02 U745 ( .Y(n695), .A0(n681), .A1(n683) );
  nor02 U746 ( .Y(n696), .A0(n681), .A1(n682) );
  nor02 U747 ( .Y(n680), .A0(n696), .A1(n697) );
  nor02 U748 ( .Y(n698), .A0(A[24]), .A1(carry_24_) );
  inv01 U749 ( .Y(n685), .A(n698) );
  nor02 U750 ( .Y(n699), .A0(B[24]), .A1(carry_24_) );
  inv01 U751 ( .Y(n687), .A(n699) );
  nor02 U752 ( .Y(n700), .A0(B[24]), .A1(A[24]) );
  inv01 U753 ( .Y(n689), .A(n700) );
  nor02 U754 ( .Y(n701), .A0(n681), .A1(n682) );
  inv01 U755 ( .Y(n691), .A(n701) );
  nor02 U756 ( .Y(n702), .A0(n684), .A1(n686) );
  inv01 U757 ( .Y(n692), .A(n702) );
  nor02 U758 ( .Y(n703), .A0(n688), .A1(n690) );
  inv01 U759 ( .Y(n693), .A(n703) );
  nor02 U760 ( .Y(n704), .A0(n694), .A1(n695) );
  inv01 U761 ( .Y(n697), .A(n704) );
  inv01 U762 ( .Y(SUM[23]), .A(n705) );
  inv02 U763 ( .Y(carry_24_), .A(n706) );
  inv02 U764 ( .Y(n707), .A(B[23]) );
  inv02 U765 ( .Y(n708), .A(A[23]) );
  inv02 U766 ( .Y(n709), .A(carry_23_) );
  nor02 U767 ( .Y(n710), .A0(n707), .A1(n711) );
  nor02 U768 ( .Y(n712), .A0(n708), .A1(n713) );
  nor02 U769 ( .Y(n714), .A0(n709), .A1(n715) );
  nor02 U770 ( .Y(n716), .A0(n709), .A1(n717) );
  nor02 U771 ( .Y(n705), .A0(n718), .A1(n719) );
  nor02 U772 ( .Y(n720), .A0(n708), .A1(n709) );
  nor02 U773 ( .Y(n721), .A0(n707), .A1(n709) );
  nor02 U774 ( .Y(n722), .A0(n707), .A1(n708) );
  nor02 U775 ( .Y(n706), .A0(n722), .A1(n723) );
  nor02 U776 ( .Y(n724), .A0(A[23]), .A1(carry_23_) );
  inv01 U777 ( .Y(n711), .A(n724) );
  nor02 U778 ( .Y(n725), .A0(B[23]), .A1(carry_23_) );
  inv01 U779 ( .Y(n713), .A(n725) );
  nor02 U780 ( .Y(n726), .A0(B[23]), .A1(A[23]) );
  inv01 U781 ( .Y(n715), .A(n726) );
  nor02 U782 ( .Y(n727), .A0(n707), .A1(n708) );
  inv01 U783 ( .Y(n717), .A(n727) );
  nor02 U784 ( .Y(n728), .A0(n710), .A1(n712) );
  inv01 U785 ( .Y(n718), .A(n728) );
  nor02 U786 ( .Y(n729), .A0(n714), .A1(n716) );
  inv01 U787 ( .Y(n719), .A(n729) );
  nor02 U788 ( .Y(n730), .A0(n720), .A1(n721) );
  inv01 U789 ( .Y(n723), .A(n730) );
  inv01 U790 ( .Y(SUM[22]), .A(n731) );
  inv02 U791 ( .Y(carry_23_), .A(n732) );
  inv02 U792 ( .Y(n733), .A(B[22]) );
  inv02 U793 ( .Y(n734), .A(A[22]) );
  inv02 U794 ( .Y(n735), .A(carry_22_) );
  nor02 U795 ( .Y(n736), .A0(n733), .A1(n737) );
  nor02 U796 ( .Y(n738), .A0(n734), .A1(n739) );
  nor02 U797 ( .Y(n740), .A0(n735), .A1(n741) );
  nor02 U798 ( .Y(n742), .A0(n735), .A1(n743) );
  nor02 U799 ( .Y(n731), .A0(n744), .A1(n745) );
  nor02 U800 ( .Y(n746), .A0(n734), .A1(n735) );
  nor02 U801 ( .Y(n747), .A0(n733), .A1(n735) );
  nor02 U802 ( .Y(n748), .A0(n733), .A1(n734) );
  nor02 U803 ( .Y(n732), .A0(n748), .A1(n749) );
  nor02 U804 ( .Y(n750), .A0(A[22]), .A1(carry_22_) );
  inv01 U805 ( .Y(n737), .A(n750) );
  nor02 U806 ( .Y(n751), .A0(B[22]), .A1(carry_22_) );
  inv01 U807 ( .Y(n739), .A(n751) );
  nor02 U808 ( .Y(n752), .A0(B[22]), .A1(A[22]) );
  inv01 U809 ( .Y(n741), .A(n752) );
  nor02 U810 ( .Y(n753), .A0(n733), .A1(n734) );
  inv01 U811 ( .Y(n743), .A(n753) );
  nor02 U812 ( .Y(n754), .A0(n736), .A1(n738) );
  inv01 U813 ( .Y(n744), .A(n754) );
  nor02 U814 ( .Y(n755), .A0(n740), .A1(n742) );
  inv01 U815 ( .Y(n745), .A(n755) );
  nor02 U816 ( .Y(n756), .A0(n746), .A1(n747) );
  inv01 U817 ( .Y(n749), .A(n756) );
  inv01 U818 ( .Y(SUM[21]), .A(n757) );
  inv02 U819 ( .Y(carry_22_), .A(n758) );
  inv02 U820 ( .Y(n759), .A(B[21]) );
  inv02 U821 ( .Y(n760), .A(A[21]) );
  inv02 U822 ( .Y(n761), .A(carry_21_) );
  nor02 U823 ( .Y(n762), .A0(n759), .A1(n763) );
  nor02 U824 ( .Y(n764), .A0(n760), .A1(n765) );
  nor02 U825 ( .Y(n766), .A0(n761), .A1(n767) );
  nor02 U826 ( .Y(n768), .A0(n761), .A1(n769) );
  nor02 U827 ( .Y(n757), .A0(n770), .A1(n771) );
  nor02 U828 ( .Y(n772), .A0(n760), .A1(n761) );
  nor02 U829 ( .Y(n773), .A0(n759), .A1(n761) );
  nor02 U830 ( .Y(n774), .A0(n759), .A1(n760) );
  nor02 U831 ( .Y(n758), .A0(n774), .A1(n775) );
  nor02 U832 ( .Y(n776), .A0(A[21]), .A1(carry_21_) );
  inv01 U833 ( .Y(n763), .A(n776) );
  nor02 U834 ( .Y(n777), .A0(B[21]), .A1(carry_21_) );
  inv01 U835 ( .Y(n765), .A(n777) );
  nor02 U836 ( .Y(n778), .A0(B[21]), .A1(A[21]) );
  inv01 U837 ( .Y(n767), .A(n778) );
  nor02 U838 ( .Y(n779), .A0(n759), .A1(n760) );
  inv01 U839 ( .Y(n769), .A(n779) );
  nor02 U840 ( .Y(n780), .A0(n762), .A1(n764) );
  inv01 U841 ( .Y(n770), .A(n780) );
  nor02 U842 ( .Y(n781), .A0(n766), .A1(n768) );
  inv01 U843 ( .Y(n771), .A(n781) );
  nor02 U844 ( .Y(n782), .A0(n772), .A1(n773) );
  inv01 U845 ( .Y(n775), .A(n782) );
  inv01 U846 ( .Y(SUM[20]), .A(n783) );
  inv02 U847 ( .Y(carry_21_), .A(n784) );
  inv02 U848 ( .Y(n785), .A(B[20]) );
  inv02 U849 ( .Y(n786), .A(A[20]) );
  inv02 U850 ( .Y(n787), .A(carry_20_) );
  nor02 U851 ( .Y(n788), .A0(n785), .A1(n789) );
  nor02 U852 ( .Y(n790), .A0(n786), .A1(n791) );
  nor02 U853 ( .Y(n792), .A0(n787), .A1(n793) );
  nor02 U854 ( .Y(n794), .A0(n787), .A1(n795) );
  nor02 U855 ( .Y(n783), .A0(n796), .A1(n797) );
  nor02 U856 ( .Y(n798), .A0(n786), .A1(n787) );
  nor02 U857 ( .Y(n799), .A0(n785), .A1(n787) );
  nor02 U858 ( .Y(n800), .A0(n785), .A1(n786) );
  nor02 U859 ( .Y(n784), .A0(n800), .A1(n801) );
  nor02 U860 ( .Y(n802), .A0(A[20]), .A1(carry_20_) );
  inv01 U861 ( .Y(n789), .A(n802) );
  nor02 U862 ( .Y(n803), .A0(B[20]), .A1(carry_20_) );
  inv01 U863 ( .Y(n791), .A(n803) );
  nor02 U864 ( .Y(n804), .A0(B[20]), .A1(A[20]) );
  inv01 U865 ( .Y(n793), .A(n804) );
  nor02 U866 ( .Y(n805), .A0(n785), .A1(n786) );
  inv01 U867 ( .Y(n795), .A(n805) );
  nor02 U868 ( .Y(n806), .A0(n788), .A1(n790) );
  inv01 U869 ( .Y(n796), .A(n806) );
  nor02 U870 ( .Y(n807), .A0(n792), .A1(n794) );
  inv01 U871 ( .Y(n797), .A(n807) );
  nor02 U872 ( .Y(n808), .A0(n798), .A1(n799) );
  inv01 U873 ( .Y(n801), .A(n808) );
  inv01 U874 ( .Y(SUM[19]), .A(n809) );
  inv02 U875 ( .Y(carry_20_), .A(n810) );
  inv02 U876 ( .Y(n811), .A(B[19]) );
  inv02 U877 ( .Y(n812), .A(A[19]) );
  inv02 U878 ( .Y(n813), .A(carry_19_) );
  nor02 U879 ( .Y(n814), .A0(n811), .A1(n815) );
  nor02 U880 ( .Y(n816), .A0(n812), .A1(n817) );
  nor02 U881 ( .Y(n818), .A0(n813), .A1(n819) );
  nor02 U882 ( .Y(n820), .A0(n813), .A1(n821) );
  nor02 U883 ( .Y(n809), .A0(n822), .A1(n823) );
  nor02 U884 ( .Y(n824), .A0(n812), .A1(n813) );
  nor02 U885 ( .Y(n825), .A0(n811), .A1(n813) );
  nor02 U886 ( .Y(n826), .A0(n811), .A1(n812) );
  nor02 U887 ( .Y(n810), .A0(n826), .A1(n827) );
  nor02 U888 ( .Y(n828), .A0(A[19]), .A1(carry_19_) );
  inv01 U889 ( .Y(n815), .A(n828) );
  nor02 U890 ( .Y(n829), .A0(B[19]), .A1(carry_19_) );
  inv01 U891 ( .Y(n817), .A(n829) );
  nor02 U892 ( .Y(n830), .A0(B[19]), .A1(A[19]) );
  inv01 U893 ( .Y(n819), .A(n830) );
  nor02 U894 ( .Y(n831), .A0(n811), .A1(n812) );
  inv01 U895 ( .Y(n821), .A(n831) );
  nor02 U896 ( .Y(n832), .A0(n814), .A1(n816) );
  inv01 U897 ( .Y(n822), .A(n832) );
  nor02 U898 ( .Y(n833), .A0(n818), .A1(n820) );
  inv01 U899 ( .Y(n823), .A(n833) );
  nor02 U900 ( .Y(n834), .A0(n824), .A1(n825) );
  inv01 U901 ( .Y(n827), .A(n834) );
  inv01 U902 ( .Y(SUM[18]), .A(n835) );
  inv02 U903 ( .Y(carry_19_), .A(n836) );
  inv02 U904 ( .Y(n837), .A(B[18]) );
  inv02 U905 ( .Y(n838), .A(A[18]) );
  inv02 U906 ( .Y(n839), .A(carry_18_) );
  nor02 U907 ( .Y(n840), .A0(n837), .A1(n841) );
  nor02 U908 ( .Y(n842), .A0(n838), .A1(n843) );
  nor02 U909 ( .Y(n844), .A0(n839), .A1(n845) );
  nor02 U910 ( .Y(n846), .A0(n839), .A1(n847) );
  nor02 U911 ( .Y(n835), .A0(n848), .A1(n849) );
  nor02 U912 ( .Y(n850), .A0(n838), .A1(n839) );
  nor02 U913 ( .Y(n851), .A0(n837), .A1(n839) );
  nor02 U914 ( .Y(n852), .A0(n837), .A1(n838) );
  nor02 U915 ( .Y(n836), .A0(n852), .A1(n853) );
  nor02 U916 ( .Y(n854), .A0(A[18]), .A1(carry_18_) );
  inv01 U917 ( .Y(n841), .A(n854) );
  nor02 U918 ( .Y(n855), .A0(B[18]), .A1(carry_18_) );
  inv01 U919 ( .Y(n843), .A(n855) );
  nor02 U920 ( .Y(n856), .A0(B[18]), .A1(A[18]) );
  inv01 U921 ( .Y(n845), .A(n856) );
  nor02 U922 ( .Y(n857), .A0(n837), .A1(n838) );
  inv01 U923 ( .Y(n847), .A(n857) );
  nor02 U924 ( .Y(n858), .A0(n840), .A1(n842) );
  inv01 U925 ( .Y(n848), .A(n858) );
  nor02 U926 ( .Y(n859), .A0(n844), .A1(n846) );
  inv01 U927 ( .Y(n849), .A(n859) );
  nor02 U928 ( .Y(n860), .A0(n850), .A1(n851) );
  inv01 U929 ( .Y(n853), .A(n860) );
  inv01 U930 ( .Y(SUM[17]), .A(n861) );
  inv02 U931 ( .Y(carry_18_), .A(n862) );
  inv02 U932 ( .Y(n863), .A(B[17]) );
  inv02 U933 ( .Y(n864), .A(A[17]) );
  inv02 U934 ( .Y(n865), .A(carry_17_) );
  nor02 U935 ( .Y(n866), .A0(n863), .A1(n867) );
  nor02 U936 ( .Y(n868), .A0(n864), .A1(n869) );
  nor02 U937 ( .Y(n870), .A0(n865), .A1(n871) );
  nor02 U938 ( .Y(n872), .A0(n865), .A1(n873) );
  nor02 U939 ( .Y(n861), .A0(n874), .A1(n875) );
  nor02 U940 ( .Y(n876), .A0(n864), .A1(n865) );
  nor02 U941 ( .Y(n877), .A0(n863), .A1(n865) );
  nor02 U942 ( .Y(n878), .A0(n863), .A1(n864) );
  nor02 U943 ( .Y(n862), .A0(n878), .A1(n879) );
  nor02 U944 ( .Y(n880), .A0(A[17]), .A1(carry_17_) );
  inv01 U945 ( .Y(n867), .A(n880) );
  nor02 U946 ( .Y(n881), .A0(B[17]), .A1(carry_17_) );
  inv01 U947 ( .Y(n869), .A(n881) );
  nor02 U948 ( .Y(n882), .A0(B[17]), .A1(A[17]) );
  inv01 U949 ( .Y(n871), .A(n882) );
  nor02 U950 ( .Y(n883), .A0(n863), .A1(n864) );
  inv01 U951 ( .Y(n873), .A(n883) );
  nor02 U952 ( .Y(n884), .A0(n866), .A1(n868) );
  inv01 U953 ( .Y(n874), .A(n884) );
  nor02 U954 ( .Y(n885), .A0(n870), .A1(n872) );
  inv01 U955 ( .Y(n875), .A(n885) );
  nor02 U956 ( .Y(n886), .A0(n876), .A1(n877) );
  inv01 U957 ( .Y(n879), .A(n886) );
  inv01 U958 ( .Y(SUM[16]), .A(n887) );
  inv02 U959 ( .Y(carry_17_), .A(n888) );
  inv02 U960 ( .Y(n889), .A(B[16]) );
  inv02 U961 ( .Y(n890), .A(A[16]) );
  inv02 U962 ( .Y(n891), .A(carry_16_) );
  nor02 U963 ( .Y(n892), .A0(n889), .A1(n893) );
  nor02 U964 ( .Y(n894), .A0(n890), .A1(n895) );
  nor02 U965 ( .Y(n896), .A0(n891), .A1(n897) );
  nor02 U966 ( .Y(n898), .A0(n891), .A1(n899) );
  nor02 U967 ( .Y(n887), .A0(n900), .A1(n901) );
  nor02 U968 ( .Y(n902), .A0(n890), .A1(n891) );
  nor02 U969 ( .Y(n903), .A0(n889), .A1(n891) );
  nor02 U970 ( .Y(n904), .A0(n889), .A1(n890) );
  nor02 U971 ( .Y(n888), .A0(n904), .A1(n905) );
  nor02 U972 ( .Y(n906), .A0(A[16]), .A1(carry_16_) );
  inv01 U973 ( .Y(n893), .A(n906) );
  nor02 U974 ( .Y(n907), .A0(B[16]), .A1(carry_16_) );
  inv01 U975 ( .Y(n895), .A(n907) );
  nor02 U976 ( .Y(n908), .A0(B[16]), .A1(A[16]) );
  inv01 U977 ( .Y(n897), .A(n908) );
  nor02 U978 ( .Y(n909), .A0(n889), .A1(n890) );
  inv01 U979 ( .Y(n899), .A(n909) );
  nor02 U980 ( .Y(n910), .A0(n892), .A1(n894) );
  inv01 U981 ( .Y(n900), .A(n910) );
  nor02 U982 ( .Y(n911), .A0(n896), .A1(n898) );
  inv01 U983 ( .Y(n901), .A(n911) );
  nor02 U984 ( .Y(n912), .A0(n902), .A1(n903) );
  inv01 U985 ( .Y(n905), .A(n912) );
  inv01 U986 ( .Y(SUM[15]), .A(n913) );
  inv02 U987 ( .Y(carry_16_), .A(n914) );
  inv02 U988 ( .Y(n915), .A(B[15]) );
  inv02 U989 ( .Y(n916), .A(A[15]) );
  inv02 U990 ( .Y(n917), .A(carry_15_) );
  nor02 U991 ( .Y(n918), .A0(n915), .A1(n919) );
  nor02 U992 ( .Y(n920), .A0(n916), .A1(n921) );
  nor02 U993 ( .Y(n922), .A0(n917), .A1(n923) );
  nor02 U994 ( .Y(n924), .A0(n917), .A1(n925) );
  nor02 U995 ( .Y(n913), .A0(n926), .A1(n927) );
  nor02 U996 ( .Y(n928), .A0(n916), .A1(n917) );
  nor02 U997 ( .Y(n929), .A0(n915), .A1(n917) );
  nor02 U998 ( .Y(n930), .A0(n915), .A1(n916) );
  nor02 U999 ( .Y(n914), .A0(n930), .A1(n931) );
  nor02 U1000 ( .Y(n932), .A0(A[15]), .A1(carry_15_) );
  inv01 U1001 ( .Y(n919), .A(n932) );
  nor02 U1002 ( .Y(n933), .A0(B[15]), .A1(carry_15_) );
  inv01 U1003 ( .Y(n921), .A(n933) );
  nor02 U1004 ( .Y(n934), .A0(B[15]), .A1(A[15]) );
  inv01 U1005 ( .Y(n923), .A(n934) );
  nor02 U1006 ( .Y(n935), .A0(n915), .A1(n916) );
  inv01 U1007 ( .Y(n925), .A(n935) );
  nor02 U1008 ( .Y(n936), .A0(n918), .A1(n920) );
  inv01 U1009 ( .Y(n926), .A(n936) );
  nor02 U1010 ( .Y(n937), .A0(n922), .A1(n924) );
  inv01 U1011 ( .Y(n927), .A(n937) );
  nor02 U1012 ( .Y(n938), .A0(n928), .A1(n929) );
  inv01 U1013 ( .Y(n931), .A(n938) );
  inv01 U1014 ( .Y(SUM[14]), .A(n939) );
  inv02 U1015 ( .Y(carry_15_), .A(n940) );
  inv02 U1016 ( .Y(n941), .A(B[14]) );
  inv02 U1017 ( .Y(n942), .A(A[14]) );
  inv02 U1018 ( .Y(n943), .A(carry_14_) );
  nor02 U1019 ( .Y(n944), .A0(n941), .A1(n945) );
  nor02 U1020 ( .Y(n946), .A0(n942), .A1(n947) );
  nor02 U1021 ( .Y(n948), .A0(n943), .A1(n949) );
  nor02 U1022 ( .Y(n950), .A0(n943), .A1(n951) );
  nor02 U1023 ( .Y(n939), .A0(n952), .A1(n953) );
  nor02 U1024 ( .Y(n954), .A0(n942), .A1(n943) );
  nor02 U1025 ( .Y(n955), .A0(n941), .A1(n943) );
  nor02 U1026 ( .Y(n956), .A0(n941), .A1(n942) );
  nor02 U1027 ( .Y(n940), .A0(n956), .A1(n957) );
  nor02 U1028 ( .Y(n958), .A0(A[14]), .A1(carry_14_) );
  inv01 U1029 ( .Y(n945), .A(n958) );
  nor02 U1030 ( .Y(n959), .A0(B[14]), .A1(carry_14_) );
  inv01 U1031 ( .Y(n947), .A(n959) );
  nor02 U1032 ( .Y(n960), .A0(B[14]), .A1(A[14]) );
  inv01 U1033 ( .Y(n949), .A(n960) );
  nor02 U1034 ( .Y(n961), .A0(n941), .A1(n942) );
  inv01 U1035 ( .Y(n951), .A(n961) );
  nor02 U1036 ( .Y(n962), .A0(n944), .A1(n946) );
  inv01 U1037 ( .Y(n952), .A(n962) );
  nor02 U1038 ( .Y(n963), .A0(n948), .A1(n950) );
  inv01 U1039 ( .Y(n953), .A(n963) );
  nor02 U1040 ( .Y(n964), .A0(n954), .A1(n955) );
  inv01 U1041 ( .Y(n957), .A(n964) );
  inv01 U1042 ( .Y(SUM[13]), .A(n965) );
  inv02 U1043 ( .Y(carry_14_), .A(n966) );
  inv02 U1044 ( .Y(n967), .A(B[13]) );
  inv02 U1045 ( .Y(n968), .A(A[13]) );
  inv02 U1046 ( .Y(n969), .A(carry_13_) );
  nor02 U1047 ( .Y(n970), .A0(n967), .A1(n971) );
  nor02 U1048 ( .Y(n972), .A0(n968), .A1(n973) );
  nor02 U1049 ( .Y(n974), .A0(n969), .A1(n975) );
  nor02 U1050 ( .Y(n976), .A0(n969), .A1(n977) );
  nor02 U1051 ( .Y(n965), .A0(n978), .A1(n979) );
  nor02 U1052 ( .Y(n980), .A0(n968), .A1(n969) );
  nor02 U1053 ( .Y(n981), .A0(n967), .A1(n969) );
  nor02 U1054 ( .Y(n982), .A0(n967), .A1(n968) );
  nor02 U1055 ( .Y(n966), .A0(n982), .A1(n983) );
  nor02 U1056 ( .Y(n984), .A0(A[13]), .A1(carry_13_) );
  inv01 U1057 ( .Y(n971), .A(n984) );
  nor02 U1058 ( .Y(n985), .A0(B[13]), .A1(carry_13_) );
  inv01 U1059 ( .Y(n973), .A(n985) );
  nor02 U1060 ( .Y(n986), .A0(B[13]), .A1(A[13]) );
  inv01 U1061 ( .Y(n975), .A(n986) );
  nor02 U1062 ( .Y(n987), .A0(n967), .A1(n968) );
  inv01 U1063 ( .Y(n977), .A(n987) );
  nor02 U1064 ( .Y(n988), .A0(n970), .A1(n972) );
  inv01 U1065 ( .Y(n978), .A(n988) );
  nor02 U1066 ( .Y(n989), .A0(n974), .A1(n976) );
  inv01 U1067 ( .Y(n979), .A(n989) );
  nor02 U1068 ( .Y(n990), .A0(n980), .A1(n981) );
  inv01 U1069 ( .Y(n983), .A(n990) );
  inv01 U1070 ( .Y(SUM[12]), .A(n991) );
  inv02 U1071 ( .Y(carry_13_), .A(n992) );
  inv02 U1072 ( .Y(n993), .A(B[12]) );
  inv02 U1073 ( .Y(n994), .A(A[12]) );
  inv02 U1074 ( .Y(n995), .A(carry_12_) );
  nor02 U1075 ( .Y(n996), .A0(n993), .A1(n997) );
  nor02 U1076 ( .Y(n998), .A0(n994), .A1(n999) );
  nor02 U1077 ( .Y(n1000), .A0(n995), .A1(n1001) );
  nor02 U1078 ( .Y(n1002), .A0(n995), .A1(n1003) );
  nor02 U1079 ( .Y(n991), .A0(n1004), .A1(n1005) );
  nor02 U1080 ( .Y(n1006), .A0(n994), .A1(n995) );
  nor02 U1081 ( .Y(n1007), .A0(n993), .A1(n995) );
  nor02 U1082 ( .Y(n1008), .A0(n993), .A1(n994) );
  nor02 U1083 ( .Y(n992), .A0(n1008), .A1(n1009) );
  nor02 U1084 ( .Y(n1010), .A0(A[12]), .A1(carry_12_) );
  inv01 U1085 ( .Y(n997), .A(n1010) );
  nor02 U1086 ( .Y(n1011), .A0(B[12]), .A1(carry_12_) );
  inv01 U1087 ( .Y(n999), .A(n1011) );
  nor02 U1088 ( .Y(n1012), .A0(B[12]), .A1(A[12]) );
  inv01 U1089 ( .Y(n1001), .A(n1012) );
  nor02 U1090 ( .Y(n1013), .A0(n993), .A1(n994) );
  inv01 U1091 ( .Y(n1003), .A(n1013) );
  nor02 U1092 ( .Y(n1014), .A0(n996), .A1(n998) );
  inv01 U1093 ( .Y(n1004), .A(n1014) );
  nor02 U1094 ( .Y(n1015), .A0(n1000), .A1(n1002) );
  inv01 U1095 ( .Y(n1005), .A(n1015) );
  nor02 U1096 ( .Y(n1016), .A0(n1006), .A1(n1007) );
  inv01 U1097 ( .Y(n1009), .A(n1016) );
  inv01 U1098 ( .Y(SUM[11]), .A(n1017) );
  inv02 U1099 ( .Y(carry_12_), .A(n1018) );
  inv02 U1100 ( .Y(n1019), .A(B[11]) );
  inv02 U1101 ( .Y(n1020), .A(A[11]) );
  inv02 U1102 ( .Y(n1021), .A(carry_11_) );
  nor02 U1103 ( .Y(n1022), .A0(n1019), .A1(n1023) );
  nor02 U1104 ( .Y(n1024), .A0(n1020), .A1(n1025) );
  nor02 U1105 ( .Y(n1026), .A0(n1021), .A1(n1027) );
  nor02 U1106 ( .Y(n1028), .A0(n1021), .A1(n1029) );
  nor02 U1107 ( .Y(n1017), .A0(n1030), .A1(n1031) );
  nor02 U1108 ( .Y(n1032), .A0(n1020), .A1(n1021) );
  nor02 U1109 ( .Y(n1033), .A0(n1019), .A1(n1021) );
  nor02 U1110 ( .Y(n1034), .A0(n1019), .A1(n1020) );
  nor02 U1111 ( .Y(n1018), .A0(n1034), .A1(n1035) );
  nor02 U1112 ( .Y(n1036), .A0(A[11]), .A1(carry_11_) );
  inv01 U1113 ( .Y(n1023), .A(n1036) );
  nor02 U1114 ( .Y(n1037), .A0(B[11]), .A1(carry_11_) );
  inv01 U1115 ( .Y(n1025), .A(n1037) );
  nor02 U1116 ( .Y(n1038), .A0(B[11]), .A1(A[11]) );
  inv01 U1117 ( .Y(n1027), .A(n1038) );
  nor02 U1118 ( .Y(n1039), .A0(n1019), .A1(n1020) );
  inv01 U1119 ( .Y(n1029), .A(n1039) );
  nor02 U1120 ( .Y(n1040), .A0(n1022), .A1(n1024) );
  inv01 U1121 ( .Y(n1030), .A(n1040) );
  nor02 U1122 ( .Y(n1041), .A0(n1026), .A1(n1028) );
  inv01 U1123 ( .Y(n1031), .A(n1041) );
  nor02 U1124 ( .Y(n1042), .A0(n1032), .A1(n1033) );
  inv01 U1125 ( .Y(n1035), .A(n1042) );
  inv01 U1126 ( .Y(SUM[10]), .A(n1043) );
  inv02 U1127 ( .Y(carry_11_), .A(n1044) );
  inv02 U1128 ( .Y(n1045), .A(B[10]) );
  inv02 U1129 ( .Y(n1046), .A(A[10]) );
  inv02 U1130 ( .Y(n1047), .A(carry_10_) );
  nor02 U1131 ( .Y(n1048), .A0(n1045), .A1(n1049) );
  nor02 U1132 ( .Y(n1050), .A0(n1046), .A1(n1051) );
  nor02 U1133 ( .Y(n1052), .A0(n1047), .A1(n1053) );
  nor02 U1134 ( .Y(n1054), .A0(n1047), .A1(n1055) );
  nor02 U1135 ( .Y(n1043), .A0(n1056), .A1(n1057) );
  nor02 U1136 ( .Y(n1058), .A0(n1046), .A1(n1047) );
  nor02 U1137 ( .Y(n1059), .A0(n1045), .A1(n1047) );
  nor02 U1138 ( .Y(n1060), .A0(n1045), .A1(n1046) );
  nor02 U1139 ( .Y(n1044), .A0(n1060), .A1(n1061) );
  nor02 U1140 ( .Y(n1062), .A0(A[10]), .A1(carry_10_) );
  inv01 U1141 ( .Y(n1049), .A(n1062) );
  nor02 U1142 ( .Y(n1063), .A0(B[10]), .A1(carry_10_) );
  inv01 U1143 ( .Y(n1051), .A(n1063) );
  nor02 U1144 ( .Y(n1064), .A0(B[10]), .A1(A[10]) );
  inv01 U1145 ( .Y(n1053), .A(n1064) );
  nor02 U1146 ( .Y(n1065), .A0(n1045), .A1(n1046) );
  inv01 U1147 ( .Y(n1055), .A(n1065) );
  nor02 U1148 ( .Y(n1066), .A0(n1048), .A1(n1050) );
  inv01 U1149 ( .Y(n1056), .A(n1066) );
  nor02 U1150 ( .Y(n1067), .A0(n1052), .A1(n1054) );
  inv01 U1151 ( .Y(n1057), .A(n1067) );
  nor02 U1152 ( .Y(n1068), .A0(n1058), .A1(n1059) );
  inv01 U1153 ( .Y(n1061), .A(n1068) );
  inv01 U1154 ( .Y(SUM[9]), .A(n1069) );
  inv02 U1155 ( .Y(carry_10_), .A(n1070) );
  inv02 U1156 ( .Y(n1071), .A(B[9]) );
  inv02 U1157 ( .Y(n1072), .A(A[9]) );
  inv02 U1158 ( .Y(n1073), .A(carry_9_) );
  nor02 U1159 ( .Y(n1074), .A0(n1071), .A1(n1075) );
  nor02 U1160 ( .Y(n1076), .A0(n1072), .A1(n1077) );
  nor02 U1161 ( .Y(n1078), .A0(n1073), .A1(n1079) );
  nor02 U1162 ( .Y(n1080), .A0(n1073), .A1(n1081) );
  nor02 U1163 ( .Y(n1069), .A0(n1082), .A1(n1083) );
  nor02 U1164 ( .Y(n1084), .A0(n1072), .A1(n1073) );
  nor02 U1165 ( .Y(n1085), .A0(n1071), .A1(n1073) );
  nor02 U1166 ( .Y(n1086), .A0(n1071), .A1(n1072) );
  nor02 U1167 ( .Y(n1070), .A0(n1086), .A1(n1087) );
  nor02 U1168 ( .Y(n1088), .A0(A[9]), .A1(carry_9_) );
  inv01 U1169 ( .Y(n1075), .A(n1088) );
  nor02 U1170 ( .Y(n1089), .A0(B[9]), .A1(carry_9_) );
  inv01 U1171 ( .Y(n1077), .A(n1089) );
  nor02 U1172 ( .Y(n1090), .A0(B[9]), .A1(A[9]) );
  inv01 U1173 ( .Y(n1079), .A(n1090) );
  nor02 U1174 ( .Y(n1091), .A0(n1071), .A1(n1072) );
  inv01 U1175 ( .Y(n1081), .A(n1091) );
  nor02 U1176 ( .Y(n1092), .A0(n1074), .A1(n1076) );
  inv01 U1177 ( .Y(n1082), .A(n1092) );
  nor02 U1178 ( .Y(n1093), .A0(n1078), .A1(n1080) );
  inv01 U1179 ( .Y(n1083), .A(n1093) );
  nor02 U1180 ( .Y(n1094), .A0(n1084), .A1(n1085) );
  inv01 U1181 ( .Y(n1087), .A(n1094) );
  inv01 U1182 ( .Y(SUM[8]), .A(n1095) );
  inv02 U1183 ( .Y(carry_9_), .A(n1096) );
  inv02 U1184 ( .Y(n1097), .A(B[8]) );
  inv02 U1185 ( .Y(n1098), .A(A[8]) );
  inv02 U1186 ( .Y(n1099), .A(carry_8_) );
  nor02 U1187 ( .Y(n1100), .A0(n1097), .A1(n1101) );
  nor02 U1188 ( .Y(n1102), .A0(n1098), .A1(n1103) );
  nor02 U1189 ( .Y(n1104), .A0(n1099), .A1(n1105) );
  nor02 U1190 ( .Y(n1106), .A0(n1099), .A1(n1107) );
  nor02 U1191 ( .Y(n1095), .A0(n1108), .A1(n1109) );
  nor02 U1192 ( .Y(n1110), .A0(n1098), .A1(n1099) );
  nor02 U1193 ( .Y(n1111), .A0(n1097), .A1(n1099) );
  nor02 U1194 ( .Y(n1112), .A0(n1097), .A1(n1098) );
  nor02 U1195 ( .Y(n1096), .A0(n1112), .A1(n1113) );
  nor02 U1196 ( .Y(n1114), .A0(A[8]), .A1(carry_8_) );
  inv01 U1197 ( .Y(n1101), .A(n1114) );
  nor02 U1198 ( .Y(n1115), .A0(B[8]), .A1(carry_8_) );
  inv01 U1199 ( .Y(n1103), .A(n1115) );
  nor02 U1200 ( .Y(n1116), .A0(B[8]), .A1(A[8]) );
  inv01 U1201 ( .Y(n1105), .A(n1116) );
  nor02 U1202 ( .Y(n1117), .A0(n1097), .A1(n1098) );
  inv01 U1203 ( .Y(n1107), .A(n1117) );
  nor02 U1204 ( .Y(n1118), .A0(n1100), .A1(n1102) );
  inv01 U1205 ( .Y(n1108), .A(n1118) );
  nor02 U1206 ( .Y(n1119), .A0(n1104), .A1(n1106) );
  inv01 U1207 ( .Y(n1109), .A(n1119) );
  nor02 U1208 ( .Y(n1120), .A0(n1110), .A1(n1111) );
  inv01 U1209 ( .Y(n1113), .A(n1120) );
  inv01 U1210 ( .Y(SUM[7]), .A(n1121) );
  inv02 U1211 ( .Y(carry_8_), .A(n1122) );
  inv02 U1212 ( .Y(n1123), .A(B[7]) );
  inv02 U1213 ( .Y(n1124), .A(A[7]) );
  inv02 U1214 ( .Y(n1125), .A(carry_7_) );
  nor02 U1215 ( .Y(n1126), .A0(n1123), .A1(n1127) );
  nor02 U1216 ( .Y(n1128), .A0(n1124), .A1(n1129) );
  nor02 U1217 ( .Y(n1130), .A0(n1125), .A1(n1131) );
  nor02 U1218 ( .Y(n1132), .A0(n1125), .A1(n1133) );
  nor02 U1219 ( .Y(n1121), .A0(n1134), .A1(n1135) );
  nor02 U1220 ( .Y(n1136), .A0(n1124), .A1(n1125) );
  nor02 U1221 ( .Y(n1137), .A0(n1123), .A1(n1125) );
  nor02 U1222 ( .Y(n1138), .A0(n1123), .A1(n1124) );
  nor02 U1223 ( .Y(n1122), .A0(n1138), .A1(n1139) );
  nor02 U1224 ( .Y(n1140), .A0(A[7]), .A1(carry_7_) );
  inv01 U1225 ( .Y(n1127), .A(n1140) );
  nor02 U1226 ( .Y(n1141), .A0(B[7]), .A1(carry_7_) );
  inv01 U1227 ( .Y(n1129), .A(n1141) );
  nor02 U1228 ( .Y(n1142), .A0(B[7]), .A1(A[7]) );
  inv01 U1229 ( .Y(n1131), .A(n1142) );
  nor02 U1230 ( .Y(n1143), .A0(n1123), .A1(n1124) );
  inv01 U1231 ( .Y(n1133), .A(n1143) );
  nor02 U1232 ( .Y(n1144), .A0(n1126), .A1(n1128) );
  inv01 U1233 ( .Y(n1134), .A(n1144) );
  nor02 U1234 ( .Y(n1145), .A0(n1130), .A1(n1132) );
  inv01 U1235 ( .Y(n1135), .A(n1145) );
  nor02 U1236 ( .Y(n1146), .A0(n1136), .A1(n1137) );
  inv01 U1237 ( .Y(n1139), .A(n1146) );
  inv01 U1238 ( .Y(SUM[6]), .A(n1147) );
  inv02 U1239 ( .Y(carry_7_), .A(n1148) );
  inv02 U1240 ( .Y(n1149), .A(B[6]) );
  inv02 U1241 ( .Y(n1150), .A(A[6]) );
  inv02 U1242 ( .Y(n1151), .A(carry_6_) );
  nor02 U1243 ( .Y(n1152), .A0(n1149), .A1(n1153) );
  nor02 U1244 ( .Y(n1154), .A0(n1150), .A1(n1155) );
  nor02 U1245 ( .Y(n1156), .A0(n1151), .A1(n1157) );
  nor02 U1246 ( .Y(n1158), .A0(n1151), .A1(n1159) );
  nor02 U1247 ( .Y(n1147), .A0(n1160), .A1(n1161) );
  nor02 U1248 ( .Y(n1162), .A0(n1150), .A1(n1151) );
  nor02 U1249 ( .Y(n1163), .A0(n1149), .A1(n1151) );
  nor02 U1250 ( .Y(n1164), .A0(n1149), .A1(n1150) );
  nor02 U1251 ( .Y(n1148), .A0(n1164), .A1(n1165) );
  nor02 U1252 ( .Y(n1166), .A0(A[6]), .A1(carry_6_) );
  inv01 U1253 ( .Y(n1153), .A(n1166) );
  nor02 U1254 ( .Y(n1167), .A0(B[6]), .A1(carry_6_) );
  inv01 U1255 ( .Y(n1155), .A(n1167) );
  nor02 U1256 ( .Y(n1168), .A0(B[6]), .A1(A[6]) );
  inv01 U1257 ( .Y(n1157), .A(n1168) );
  nor02 U1258 ( .Y(n1169), .A0(n1149), .A1(n1150) );
  inv01 U1259 ( .Y(n1159), .A(n1169) );
  nor02 U1260 ( .Y(n1170), .A0(n1152), .A1(n1154) );
  inv01 U1261 ( .Y(n1160), .A(n1170) );
  nor02 U1262 ( .Y(n1171), .A0(n1156), .A1(n1158) );
  inv01 U1263 ( .Y(n1161), .A(n1171) );
  nor02 U1264 ( .Y(n1172), .A0(n1162), .A1(n1163) );
  inv01 U1265 ( .Y(n1165), .A(n1172) );
  inv01 U1266 ( .Y(SUM[5]), .A(n1173) );
  inv02 U1267 ( .Y(carry_6_), .A(n1174) );
  inv02 U1268 ( .Y(n1175), .A(B[5]) );
  inv02 U1269 ( .Y(n1176), .A(A[5]) );
  inv02 U1270 ( .Y(n1177), .A(carry_5_) );
  nor02 U1271 ( .Y(n1178), .A0(n1175), .A1(n1179) );
  nor02 U1272 ( .Y(n1180), .A0(n1176), .A1(n1181) );
  nor02 U1273 ( .Y(n1182), .A0(n1177), .A1(n1183) );
  nor02 U1274 ( .Y(n1184), .A0(n1177), .A1(n1185) );
  nor02 U1275 ( .Y(n1173), .A0(n1186), .A1(n1187) );
  nor02 U1276 ( .Y(n1188), .A0(n1176), .A1(n1177) );
  nor02 U1277 ( .Y(n1189), .A0(n1175), .A1(n1177) );
  nor02 U1278 ( .Y(n1190), .A0(n1175), .A1(n1176) );
  nor02 U1279 ( .Y(n1174), .A0(n1190), .A1(n1191) );
  nor02 U1280 ( .Y(n1192), .A0(A[5]), .A1(carry_5_) );
  inv01 U1281 ( .Y(n1179), .A(n1192) );
  nor02 U1282 ( .Y(n1193), .A0(B[5]), .A1(carry_5_) );
  inv01 U1283 ( .Y(n1181), .A(n1193) );
  nor02 U1284 ( .Y(n1194), .A0(B[5]), .A1(A[5]) );
  inv01 U1285 ( .Y(n1183), .A(n1194) );
  nor02 U1286 ( .Y(n1195), .A0(n1175), .A1(n1176) );
  inv01 U1287 ( .Y(n1185), .A(n1195) );
  nor02 U1288 ( .Y(n1196), .A0(n1178), .A1(n1180) );
  inv01 U1289 ( .Y(n1186), .A(n1196) );
  nor02 U1290 ( .Y(n1197), .A0(n1182), .A1(n1184) );
  inv01 U1291 ( .Y(n1187), .A(n1197) );
  nor02 U1292 ( .Y(n1198), .A0(n1188), .A1(n1189) );
  inv01 U1293 ( .Y(n1191), .A(n1198) );
  inv01 U1294 ( .Y(SUM[4]), .A(n1199) );
  inv02 U1295 ( .Y(carry_5_), .A(n1200) );
  inv02 U1296 ( .Y(n1201), .A(B[4]) );
  inv02 U1297 ( .Y(n1202), .A(A[4]) );
  inv02 U1298 ( .Y(n1203), .A(carry_4_) );
  nor02 U1299 ( .Y(n1204), .A0(n1201), .A1(n1205) );
  nor02 U1300 ( .Y(n1206), .A0(n1202), .A1(n1207) );
  nor02 U1301 ( .Y(n1208), .A0(n1203), .A1(n1209) );
  nor02 U1302 ( .Y(n1210), .A0(n1203), .A1(n1211) );
  nor02 U1303 ( .Y(n1199), .A0(n1212), .A1(n1213) );
  nor02 U1304 ( .Y(n1214), .A0(n1202), .A1(n1203) );
  nor02 U1305 ( .Y(n1215), .A0(n1201), .A1(n1203) );
  nor02 U1306 ( .Y(n1216), .A0(n1201), .A1(n1202) );
  nor02 U1307 ( .Y(n1200), .A0(n1216), .A1(n1217) );
  nor02 U1308 ( .Y(n1218), .A0(A[4]), .A1(carry_4_) );
  inv01 U1309 ( .Y(n1205), .A(n1218) );
  nor02 U1310 ( .Y(n1219), .A0(B[4]), .A1(carry_4_) );
  inv01 U1311 ( .Y(n1207), .A(n1219) );
  nor02 U1312 ( .Y(n1220), .A0(B[4]), .A1(A[4]) );
  inv01 U1313 ( .Y(n1209), .A(n1220) );
  nor02 U1314 ( .Y(n1221), .A0(n1201), .A1(n1202) );
  inv01 U1315 ( .Y(n1211), .A(n1221) );
  nor02 U1316 ( .Y(n1222), .A0(n1204), .A1(n1206) );
  inv01 U1317 ( .Y(n1212), .A(n1222) );
  nor02 U1318 ( .Y(n1223), .A0(n1208), .A1(n1210) );
  inv01 U1319 ( .Y(n1213), .A(n1223) );
  nor02 U1320 ( .Y(n1224), .A0(n1214), .A1(n1215) );
  inv01 U1321 ( .Y(n1217), .A(n1224) );
  inv01 U1322 ( .Y(SUM[3]), .A(n1225) );
  inv02 U1323 ( .Y(carry_4_), .A(n1226) );
  inv02 U1324 ( .Y(n1227), .A(n1303) );
  inv02 U1325 ( .Y(n1228), .A(A[3]) );
  inv02 U1326 ( .Y(n1229), .A(carry_3_) );
  nor02 U1327 ( .Y(n1230), .A0(n1227), .A1(n1231) );
  nor02 U1328 ( .Y(n1232), .A0(n1228), .A1(n1233) );
  nor02 U1329 ( .Y(n1234), .A0(n1229), .A1(n1235) );
  nor02 U1330 ( .Y(n1236), .A0(n1229), .A1(n1237) );
  nor02 U1331 ( .Y(n1225), .A0(n1238), .A1(n1239) );
  nor02 U1332 ( .Y(n1240), .A0(n1228), .A1(n1229) );
  nor02 U1333 ( .Y(n1241), .A0(n1227), .A1(n1229) );
  nor02 U1334 ( .Y(n1242), .A0(n1227), .A1(n1228) );
  nor02 U1335 ( .Y(n1226), .A0(n1242), .A1(n1243) );
  nor02 U1336 ( .Y(n1244), .A0(A[3]), .A1(carry_3_) );
  inv01 U1337 ( .Y(n1231), .A(n1244) );
  nor02 U1338 ( .Y(n1245), .A0(n1303), .A1(carry_3_) );
  inv01 U1339 ( .Y(n1233), .A(n1245) );
  nor02 U1340 ( .Y(n1246), .A0(n1303), .A1(A[3]) );
  inv01 U1341 ( .Y(n1235), .A(n1246) );
  nor02 U1342 ( .Y(n1247), .A0(n1227), .A1(n1228) );
  inv01 U1343 ( .Y(n1237), .A(n1247) );
  nor02 U1344 ( .Y(n1248), .A0(n1230), .A1(n1232) );
  inv01 U1345 ( .Y(n1238), .A(n1248) );
  nor02 U1346 ( .Y(n1249), .A0(n1234), .A1(n1236) );
  inv01 U1347 ( .Y(n1239), .A(n1249) );
  nor02 U1348 ( .Y(n1250), .A0(n1240), .A1(n1241) );
  inv01 U1349 ( .Y(n1243), .A(n1250) );
  inv01 U1350 ( .Y(SUM[2]), .A(n1251) );
  inv02 U1351 ( .Y(carry_3_), .A(n1252) );
  inv02 U1352 ( .Y(n1253), .A(B[2]) );
  inv02 U1353 ( .Y(n1254), .A(A[2]) );
  inv02 U1354 ( .Y(n1255), .A(carry_2_) );
  nor02 U1355 ( .Y(n1256), .A0(n1253), .A1(n1257) );
  nor02 U1356 ( .Y(n1258), .A0(n1254), .A1(n1259) );
  nor02 U1357 ( .Y(n1260), .A0(n1255), .A1(n1261) );
  nor02 U1358 ( .Y(n1262), .A0(n1255), .A1(n1263) );
  nor02 U1359 ( .Y(n1251), .A0(n1264), .A1(n1265) );
  nor02 U1360 ( .Y(n1266), .A0(n1254), .A1(n1255) );
  nor02 U1361 ( .Y(n1267), .A0(n1253), .A1(n1255) );
  nor02 U1362 ( .Y(n1268), .A0(n1253), .A1(n1254) );
  nor02 U1363 ( .Y(n1252), .A0(n1268), .A1(n1269) );
  nor02 U1364 ( .Y(n1270), .A0(A[2]), .A1(carry_2_) );
  inv01 U1365 ( .Y(n1257), .A(n1270) );
  nor02 U1366 ( .Y(n1271), .A0(B[2]), .A1(carry_2_) );
  inv01 U1367 ( .Y(n1259), .A(n1271) );
  nor02 U1368 ( .Y(n1272), .A0(B[2]), .A1(A[2]) );
  inv01 U1369 ( .Y(n1261), .A(n1272) );
  nor02 U1370 ( .Y(n1273), .A0(n1253), .A1(n1254) );
  inv01 U1371 ( .Y(n1263), .A(n1273) );
  nor02 U1372 ( .Y(n1274), .A0(n1256), .A1(n1258) );
  inv01 U1373 ( .Y(n1264), .A(n1274) );
  nor02 U1374 ( .Y(n1275), .A0(n1260), .A1(n1262) );
  inv01 U1375 ( .Y(n1265), .A(n1275) );
  nor02 U1376 ( .Y(n1276), .A0(n1266), .A1(n1267) );
  inv01 U1377 ( .Y(n1269), .A(n1276) );
  inv01 U1378 ( .Y(SUM[1]), .A(n1277) );
  inv02 U1379 ( .Y(carry_2_), .A(n1278) );
  inv02 U1380 ( .Y(n1279), .A(B[1]) );
  inv02 U1381 ( .Y(n1280), .A(A[1]) );
  inv02 U1382 ( .Y(n1281), .A(n2) );
  nor02 U1383 ( .Y(n1282), .A0(n1279), .A1(n1283) );
  nor02 U1384 ( .Y(n1284), .A0(n1280), .A1(n1285) );
  nor02 U1385 ( .Y(n1286), .A0(n1281), .A1(n1287) );
  nor02 U1386 ( .Y(n1288), .A0(n1281), .A1(n1289) );
  nor02 U1387 ( .Y(n1277), .A0(n1290), .A1(n1291) );
  nor02 U1388 ( .Y(n1292), .A0(n1280), .A1(n1281) );
  nor02 U1389 ( .Y(n1293), .A0(n1279), .A1(n1281) );
  nor02 U1390 ( .Y(n1294), .A0(n1279), .A1(n1280) );
  nor02 U1391 ( .Y(n1278), .A0(n1294), .A1(n1295) );
  nor02 U1392 ( .Y(n1296), .A0(A[1]), .A1(n2) );
  inv01 U1393 ( .Y(n1283), .A(n1296) );
  nor02 U1394 ( .Y(n1297), .A0(B[1]), .A1(n2) );
  inv01 U1395 ( .Y(n1285), .A(n1297) );
  nor02 U1396 ( .Y(n1298), .A0(B[1]), .A1(A[1]) );
  inv01 U1397 ( .Y(n1287), .A(n1298) );
  nor02 U1398 ( .Y(n1299), .A0(n1279), .A1(n1280) );
  inv01 U1399 ( .Y(n1289), .A(n1299) );
  nor02 U1400 ( .Y(n1300), .A0(n1282), .A1(n1284) );
  inv01 U1401 ( .Y(n1290), .A(n1300) );
  nor02 U1402 ( .Y(n1301), .A0(n1286), .A1(n1288) );
  inv01 U1403 ( .Y(n1291), .A(n1301) );
  nor02 U1404 ( .Y(n1302), .A0(n1292), .A1(n1293) );
  inv01 U1405 ( .Y(n1295), .A(n1302) );
  buf02 U1406 ( .Y(n1303), .A(B[3]) );
  xor2 U1407 ( .Y(SUM[0]), .A0(B[0]), .A1(A[0]) );
  fadd1 U1_51 ( .S(SUM[51]), .A(A[51]), .B(B[51]), .CI(carry_51_) );
endmodule


module sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_sub_52_0 ( A, B, CI, DIFF, CO );
  input [51:0] A;
  input [51:0] B;
  output [51:0] DIFF;
  input CI;
  output CO;
  wire   carry_51_, carry_50_, carry_49_, carry_48_, carry_47_, carry_46_,
         carry_45_, carry_44_, carry_43_, carry_42_, carry_41_, carry_40_,
         carry_39_, carry_38_, carry_37_, carry_36_, carry_35_, carry_34_,
         carry_33_, carry_32_, carry_31_, carry_30_, carry_29_, carry_28_,
         carry_27_, carry_26_, carry_25_, carry_24_, carry_23_, carry_22_,
         carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, carry_6_, carry_5_, carry_4_, carry_3_,
         carry_2_, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314;
  wire   [51:0] B_not;

  xor2 U6 ( .Y(n5), .A0(B_not[0]), .A1(A[0]) );
  inv01 U7 ( .Y(DIFF[0]), .A(n5) );
  inv01 U8 ( .Y(DIFF[50]), .A(n7) );
  inv02 U9 ( .Y(carry_51_), .A(n8) );
  inv02 U10 ( .Y(n9), .A(B_not[50]) );
  inv02 U11 ( .Y(n10), .A(A[50]) );
  inv02 U12 ( .Y(n11), .A(carry_50_) );
  nor02 U13 ( .Y(n12), .A0(n9), .A1(n13) );
  nor02 U14 ( .Y(n14), .A0(n10), .A1(n15) );
  nor02 U15 ( .Y(n16), .A0(n11), .A1(n17) );
  nor02 U16 ( .Y(n18), .A0(n11), .A1(n19) );
  nor02 U17 ( .Y(n7), .A0(n20), .A1(n21) );
  nor02 U18 ( .Y(n22), .A0(n10), .A1(n11) );
  nor02 U19 ( .Y(n23), .A0(n9), .A1(n11) );
  nor02 U20 ( .Y(n24), .A0(n9), .A1(n10) );
  nor02 U21 ( .Y(n8), .A0(n24), .A1(n25) );
  nor02 U22 ( .Y(n26), .A0(A[50]), .A1(carry_50_) );
  inv01 U23 ( .Y(n13), .A(n26) );
  nor02 U24 ( .Y(n27), .A0(B_not[50]), .A1(carry_50_) );
  inv01 U25 ( .Y(n15), .A(n27) );
  nor02 U26 ( .Y(n28), .A0(B_not[50]), .A1(A[50]) );
  inv01 U27 ( .Y(n17), .A(n28) );
  nor02 U28 ( .Y(n29), .A0(n9), .A1(n10) );
  inv01 U29 ( .Y(n19), .A(n29) );
  nor02 U30 ( .Y(n30), .A0(n12), .A1(n14) );
  inv01 U31 ( .Y(n20), .A(n30) );
  nor02 U32 ( .Y(n31), .A0(n16), .A1(n18) );
  inv01 U33 ( .Y(n21), .A(n31) );
  nor02 U34 ( .Y(n32), .A0(n22), .A1(n23) );
  inv01 U35 ( .Y(n25), .A(n32) );
  inv02 U36 ( .Y(B_not[50]), .A(B[50]) );
  inv01 U37 ( .Y(DIFF[49]), .A(n33) );
  inv02 U38 ( .Y(carry_50_), .A(n34) );
  inv02 U39 ( .Y(n35), .A(B_not[49]) );
  inv02 U40 ( .Y(n36), .A(A[49]) );
  inv02 U41 ( .Y(n37), .A(carry_49_) );
  nor02 U42 ( .Y(n38), .A0(n35), .A1(n39) );
  nor02 U43 ( .Y(n40), .A0(n36), .A1(n41) );
  nor02 U44 ( .Y(n42), .A0(n37), .A1(n43) );
  nor02 U45 ( .Y(n44), .A0(n37), .A1(n45) );
  nor02 U46 ( .Y(n33), .A0(n46), .A1(n47) );
  nor02 U47 ( .Y(n48), .A0(n36), .A1(n37) );
  nor02 U48 ( .Y(n49), .A0(n35), .A1(n37) );
  nor02 U49 ( .Y(n50), .A0(n35), .A1(n36) );
  nor02 U50 ( .Y(n34), .A0(n50), .A1(n51) );
  nor02 U51 ( .Y(n52), .A0(A[49]), .A1(carry_49_) );
  inv01 U52 ( .Y(n39), .A(n52) );
  nor02 U53 ( .Y(n53), .A0(B_not[49]), .A1(carry_49_) );
  inv01 U54 ( .Y(n41), .A(n53) );
  nor02 U55 ( .Y(n54), .A0(B_not[49]), .A1(A[49]) );
  inv01 U56 ( .Y(n43), .A(n54) );
  nor02 U57 ( .Y(n55), .A0(n35), .A1(n36) );
  inv01 U58 ( .Y(n45), .A(n55) );
  nor02 U59 ( .Y(n56), .A0(n38), .A1(n40) );
  inv01 U60 ( .Y(n46), .A(n56) );
  nor02 U61 ( .Y(n57), .A0(n42), .A1(n44) );
  inv01 U62 ( .Y(n47), .A(n57) );
  nor02 U63 ( .Y(n58), .A0(n48), .A1(n49) );
  inv01 U64 ( .Y(n51), .A(n58) );
  inv02 U65 ( .Y(B_not[49]), .A(B[49]) );
  inv01 U66 ( .Y(DIFF[48]), .A(n59) );
  inv02 U67 ( .Y(carry_49_), .A(n60) );
  inv02 U68 ( .Y(n61), .A(B_not[48]) );
  inv02 U69 ( .Y(n62), .A(A[48]) );
  inv02 U70 ( .Y(n63), .A(carry_48_) );
  nor02 U71 ( .Y(n64), .A0(n61), .A1(n65) );
  nor02 U72 ( .Y(n66), .A0(n62), .A1(n67) );
  nor02 U73 ( .Y(n68), .A0(n63), .A1(n69) );
  nor02 U74 ( .Y(n70), .A0(n63), .A1(n71) );
  nor02 U75 ( .Y(n59), .A0(n72), .A1(n73) );
  nor02 U76 ( .Y(n74), .A0(n62), .A1(n63) );
  nor02 U77 ( .Y(n75), .A0(n61), .A1(n63) );
  nor02 U78 ( .Y(n76), .A0(n61), .A1(n62) );
  nor02 U79 ( .Y(n60), .A0(n76), .A1(n77) );
  nor02 U80 ( .Y(n78), .A0(A[48]), .A1(carry_48_) );
  inv01 U81 ( .Y(n65), .A(n78) );
  nor02 U82 ( .Y(n79), .A0(B_not[48]), .A1(carry_48_) );
  inv01 U83 ( .Y(n67), .A(n79) );
  nor02 U84 ( .Y(n80), .A0(B_not[48]), .A1(A[48]) );
  inv01 U85 ( .Y(n69), .A(n80) );
  nor02 U86 ( .Y(n81), .A0(n61), .A1(n62) );
  inv01 U87 ( .Y(n71), .A(n81) );
  nor02 U88 ( .Y(n82), .A0(n64), .A1(n66) );
  inv01 U89 ( .Y(n72), .A(n82) );
  nor02 U90 ( .Y(n83), .A0(n68), .A1(n70) );
  inv01 U91 ( .Y(n73), .A(n83) );
  nor02 U92 ( .Y(n84), .A0(n74), .A1(n75) );
  inv01 U93 ( .Y(n77), .A(n84) );
  inv01 U94 ( .Y(DIFF[47]), .A(n85) );
  inv02 U95 ( .Y(carry_48_), .A(n86) );
  inv02 U96 ( .Y(n87), .A(B_not[47]) );
  inv02 U97 ( .Y(n88), .A(A[47]) );
  inv02 U98 ( .Y(n89), .A(carry_47_) );
  nor02 U99 ( .Y(n90), .A0(n87), .A1(n91) );
  nor02 U100 ( .Y(n92), .A0(n88), .A1(n93) );
  nor02 U101 ( .Y(n94), .A0(n89), .A1(n95) );
  nor02 U102 ( .Y(n96), .A0(n89), .A1(n97) );
  nor02 U103 ( .Y(n85), .A0(n98), .A1(n99) );
  nor02 U104 ( .Y(n100), .A0(n88), .A1(n89) );
  nor02 U105 ( .Y(n101), .A0(n87), .A1(n89) );
  nor02 U106 ( .Y(n102), .A0(n87), .A1(n88) );
  nor02 U107 ( .Y(n86), .A0(n102), .A1(n103) );
  nor02 U108 ( .Y(n104), .A0(A[47]), .A1(carry_47_) );
  inv01 U109 ( .Y(n91), .A(n104) );
  nor02 U110 ( .Y(n105), .A0(B_not[47]), .A1(carry_47_) );
  inv01 U111 ( .Y(n93), .A(n105) );
  nor02 U112 ( .Y(n106), .A0(B_not[47]), .A1(A[47]) );
  inv01 U113 ( .Y(n95), .A(n106) );
  nor02 U114 ( .Y(n107), .A0(n87), .A1(n88) );
  inv01 U115 ( .Y(n97), .A(n107) );
  nor02 U116 ( .Y(n108), .A0(n90), .A1(n92) );
  inv01 U117 ( .Y(n98), .A(n108) );
  nor02 U118 ( .Y(n109), .A0(n94), .A1(n96) );
  inv01 U119 ( .Y(n99), .A(n109) );
  nor02 U120 ( .Y(n110), .A0(n100), .A1(n101) );
  inv01 U121 ( .Y(n103), .A(n110) );
  inv01 U122 ( .Y(DIFF[46]), .A(n111) );
  inv02 U123 ( .Y(carry_47_), .A(n112) );
  inv02 U124 ( .Y(n113), .A(B_not[46]) );
  inv02 U125 ( .Y(n114), .A(A[46]) );
  inv02 U126 ( .Y(n115), .A(carry_46_) );
  nor02 U127 ( .Y(n116), .A0(n113), .A1(n117) );
  nor02 U128 ( .Y(n118), .A0(n114), .A1(n119) );
  nor02 U129 ( .Y(n120), .A0(n115), .A1(n121) );
  nor02 U130 ( .Y(n122), .A0(n115), .A1(n123) );
  nor02 U131 ( .Y(n111), .A0(n124), .A1(n125) );
  nor02 U132 ( .Y(n126), .A0(n114), .A1(n115) );
  nor02 U133 ( .Y(n127), .A0(n113), .A1(n115) );
  nor02 U134 ( .Y(n128), .A0(n113), .A1(n114) );
  nor02 U135 ( .Y(n112), .A0(n128), .A1(n129) );
  nor02 U136 ( .Y(n130), .A0(A[46]), .A1(carry_46_) );
  inv01 U137 ( .Y(n117), .A(n130) );
  nor02 U138 ( .Y(n131), .A0(B_not[46]), .A1(carry_46_) );
  inv01 U139 ( .Y(n119), .A(n131) );
  nor02 U140 ( .Y(n132), .A0(B_not[46]), .A1(A[46]) );
  inv01 U141 ( .Y(n121), .A(n132) );
  nor02 U142 ( .Y(n133), .A0(n113), .A1(n114) );
  inv01 U143 ( .Y(n123), .A(n133) );
  nor02 U144 ( .Y(n134), .A0(n116), .A1(n118) );
  inv01 U145 ( .Y(n124), .A(n134) );
  nor02 U146 ( .Y(n135), .A0(n120), .A1(n122) );
  inv01 U147 ( .Y(n125), .A(n135) );
  nor02 U148 ( .Y(n136), .A0(n126), .A1(n127) );
  inv01 U149 ( .Y(n129), .A(n136) );
  inv02 U150 ( .Y(B_not[46]), .A(B[46]) );
  inv01 U151 ( .Y(DIFF[45]), .A(n137) );
  inv02 U152 ( .Y(carry_46_), .A(n138) );
  inv02 U153 ( .Y(n139), .A(B_not[45]) );
  inv02 U154 ( .Y(n140), .A(A[45]) );
  inv02 U155 ( .Y(n141), .A(carry_45_) );
  nor02 U156 ( .Y(n142), .A0(n139), .A1(n143) );
  nor02 U157 ( .Y(n144), .A0(n140), .A1(n145) );
  nor02 U158 ( .Y(n146), .A0(n141), .A1(n147) );
  nor02 U159 ( .Y(n148), .A0(n141), .A1(n149) );
  nor02 U160 ( .Y(n137), .A0(n150), .A1(n151) );
  nor02 U161 ( .Y(n152), .A0(n140), .A1(n141) );
  nor02 U162 ( .Y(n153), .A0(n139), .A1(n141) );
  nor02 U163 ( .Y(n154), .A0(n139), .A1(n140) );
  nor02 U164 ( .Y(n138), .A0(n154), .A1(n155) );
  nor02 U165 ( .Y(n156), .A0(A[45]), .A1(carry_45_) );
  inv01 U166 ( .Y(n143), .A(n156) );
  nor02 U167 ( .Y(n157), .A0(B_not[45]), .A1(carry_45_) );
  inv01 U168 ( .Y(n145), .A(n157) );
  nor02 U169 ( .Y(n158), .A0(B_not[45]), .A1(A[45]) );
  inv01 U170 ( .Y(n147), .A(n158) );
  nor02 U171 ( .Y(n159), .A0(n139), .A1(n140) );
  inv01 U172 ( .Y(n149), .A(n159) );
  nor02 U173 ( .Y(n160), .A0(n142), .A1(n144) );
  inv01 U174 ( .Y(n150), .A(n160) );
  nor02 U175 ( .Y(n161), .A0(n146), .A1(n148) );
  inv01 U176 ( .Y(n151), .A(n161) );
  nor02 U177 ( .Y(n162), .A0(n152), .A1(n153) );
  inv01 U178 ( .Y(n155), .A(n162) );
  inv01 U179 ( .Y(DIFF[44]), .A(n163) );
  inv02 U180 ( .Y(carry_45_), .A(n164) );
  inv02 U181 ( .Y(n165), .A(B_not[44]) );
  inv02 U182 ( .Y(n166), .A(A[44]) );
  inv02 U183 ( .Y(n167), .A(carry_44_) );
  nor02 U184 ( .Y(n168), .A0(n165), .A1(n169) );
  nor02 U185 ( .Y(n170), .A0(n166), .A1(n171) );
  nor02 U186 ( .Y(n172), .A0(n167), .A1(n173) );
  nor02 U187 ( .Y(n174), .A0(n167), .A1(n175) );
  nor02 U188 ( .Y(n163), .A0(n176), .A1(n177) );
  nor02 U189 ( .Y(n178), .A0(n166), .A1(n167) );
  nor02 U190 ( .Y(n179), .A0(n165), .A1(n167) );
  nor02 U191 ( .Y(n180), .A0(n165), .A1(n166) );
  nor02 U192 ( .Y(n164), .A0(n180), .A1(n181) );
  nor02 U193 ( .Y(n182), .A0(A[44]), .A1(carry_44_) );
  inv01 U194 ( .Y(n169), .A(n182) );
  nor02 U195 ( .Y(n183), .A0(B_not[44]), .A1(carry_44_) );
  inv01 U196 ( .Y(n171), .A(n183) );
  nor02 U197 ( .Y(n184), .A0(B_not[44]), .A1(A[44]) );
  inv01 U198 ( .Y(n173), .A(n184) );
  nor02 U199 ( .Y(n185), .A0(n165), .A1(n166) );
  inv01 U200 ( .Y(n175), .A(n185) );
  nor02 U201 ( .Y(n186), .A0(n168), .A1(n170) );
  inv01 U202 ( .Y(n176), .A(n186) );
  nor02 U203 ( .Y(n187), .A0(n172), .A1(n174) );
  inv01 U204 ( .Y(n177), .A(n187) );
  nor02 U205 ( .Y(n188), .A0(n178), .A1(n179) );
  inv01 U206 ( .Y(n181), .A(n188) );
  inv01 U207 ( .Y(DIFF[43]), .A(n189) );
  inv02 U208 ( .Y(carry_44_), .A(n190) );
  inv02 U209 ( .Y(n191), .A(B_not[43]) );
  inv02 U210 ( .Y(n192), .A(A[43]) );
  inv02 U211 ( .Y(n193), .A(carry_43_) );
  nor02 U212 ( .Y(n194), .A0(n191), .A1(n195) );
  nor02 U213 ( .Y(n196), .A0(n192), .A1(n197) );
  nor02 U214 ( .Y(n198), .A0(n193), .A1(n199) );
  nor02 U215 ( .Y(n200), .A0(n193), .A1(n201) );
  nor02 U216 ( .Y(n189), .A0(n202), .A1(n203) );
  nor02 U217 ( .Y(n204), .A0(n192), .A1(n193) );
  nor02 U218 ( .Y(n205), .A0(n191), .A1(n193) );
  nor02 U219 ( .Y(n206), .A0(n191), .A1(n192) );
  nor02 U220 ( .Y(n190), .A0(n206), .A1(n207) );
  nor02 U221 ( .Y(n208), .A0(A[43]), .A1(carry_43_) );
  inv01 U222 ( .Y(n195), .A(n208) );
  nor02 U223 ( .Y(n209), .A0(B_not[43]), .A1(carry_43_) );
  inv01 U224 ( .Y(n197), .A(n209) );
  nor02 U225 ( .Y(n210), .A0(B_not[43]), .A1(A[43]) );
  inv01 U226 ( .Y(n199), .A(n210) );
  nor02 U227 ( .Y(n211), .A0(n191), .A1(n192) );
  inv01 U228 ( .Y(n201), .A(n211) );
  nor02 U229 ( .Y(n212), .A0(n194), .A1(n196) );
  inv01 U230 ( .Y(n202), .A(n212) );
  nor02 U231 ( .Y(n213), .A0(n198), .A1(n200) );
  inv01 U232 ( .Y(n203), .A(n213) );
  nor02 U233 ( .Y(n214), .A0(n204), .A1(n205) );
  inv01 U234 ( .Y(n207), .A(n214) );
  inv02 U235 ( .Y(B_not[43]), .A(B[43]) );
  inv01 U236 ( .Y(DIFF[22]), .A(n215) );
  inv02 U237 ( .Y(carry_23_), .A(n216) );
  inv02 U238 ( .Y(n217), .A(B_not[22]) );
  inv02 U239 ( .Y(n218), .A(A[22]) );
  inv02 U240 ( .Y(n219), .A(carry_22_) );
  nor02 U241 ( .Y(n220), .A0(n217), .A1(n221) );
  nor02 U242 ( .Y(n222), .A0(n218), .A1(n223) );
  nor02 U243 ( .Y(n224), .A0(n219), .A1(n225) );
  nor02 U244 ( .Y(n226), .A0(n219), .A1(n227) );
  nor02 U245 ( .Y(n215), .A0(n228), .A1(n229) );
  nor02 U246 ( .Y(n230), .A0(n218), .A1(n219) );
  nor02 U247 ( .Y(n231), .A0(n217), .A1(n219) );
  nor02 U248 ( .Y(n232), .A0(n217), .A1(n218) );
  nor02 U249 ( .Y(n216), .A0(n232), .A1(n233) );
  nor02 U250 ( .Y(n234), .A0(A[22]), .A1(carry_22_) );
  inv01 U251 ( .Y(n221), .A(n234) );
  nor02 U252 ( .Y(n235), .A0(B_not[22]), .A1(carry_22_) );
  inv01 U253 ( .Y(n223), .A(n235) );
  nor02 U254 ( .Y(n236), .A0(B_not[22]), .A1(A[22]) );
  inv01 U255 ( .Y(n225), .A(n236) );
  nor02 U256 ( .Y(n237), .A0(n217), .A1(n218) );
  inv01 U257 ( .Y(n227), .A(n237) );
  nor02 U258 ( .Y(n238), .A0(n220), .A1(n222) );
  inv01 U259 ( .Y(n228), .A(n238) );
  nor02 U260 ( .Y(n239), .A0(n224), .A1(n226) );
  inv01 U261 ( .Y(n229), .A(n239) );
  nor02 U262 ( .Y(n240), .A0(n230), .A1(n231) );
  inv01 U263 ( .Y(n233), .A(n240) );
  inv01 U264 ( .Y(DIFF[42]), .A(n241) );
  inv02 U265 ( .Y(carry_43_), .A(n242) );
  inv02 U266 ( .Y(n243), .A(B_not[42]) );
  inv02 U267 ( .Y(n244), .A(A[42]) );
  inv02 U268 ( .Y(n245), .A(carry_42_) );
  nor02 U269 ( .Y(n246), .A0(n243), .A1(n247) );
  nor02 U270 ( .Y(n248), .A0(n244), .A1(n249) );
  nor02 U271 ( .Y(n250), .A0(n245), .A1(n251) );
  nor02 U272 ( .Y(n252), .A0(n245), .A1(n253) );
  nor02 U273 ( .Y(n241), .A0(n254), .A1(n255) );
  nor02 U274 ( .Y(n256), .A0(n244), .A1(n245) );
  nor02 U275 ( .Y(n257), .A0(n243), .A1(n245) );
  nor02 U276 ( .Y(n258), .A0(n243), .A1(n244) );
  nor02 U277 ( .Y(n242), .A0(n258), .A1(n259) );
  nor02 U278 ( .Y(n260), .A0(A[42]), .A1(carry_42_) );
  inv01 U279 ( .Y(n247), .A(n260) );
  nor02 U280 ( .Y(n261), .A0(B_not[42]), .A1(carry_42_) );
  inv01 U281 ( .Y(n249), .A(n261) );
  nor02 U282 ( .Y(n262), .A0(B_not[42]), .A1(A[42]) );
  inv01 U283 ( .Y(n251), .A(n262) );
  nor02 U284 ( .Y(n263), .A0(n243), .A1(n244) );
  inv01 U285 ( .Y(n253), .A(n263) );
  nor02 U286 ( .Y(n264), .A0(n246), .A1(n248) );
  inv01 U287 ( .Y(n254), .A(n264) );
  nor02 U288 ( .Y(n265), .A0(n250), .A1(n252) );
  inv01 U289 ( .Y(n255), .A(n265) );
  nor02 U290 ( .Y(n266), .A0(n256), .A1(n257) );
  inv01 U291 ( .Y(n259), .A(n266) );
  inv02 U292 ( .Y(B_not[42]), .A(B[42]) );
  inv01 U293 ( .Y(DIFF[23]), .A(n267) );
  inv02 U294 ( .Y(carry_24_), .A(n268) );
  inv02 U295 ( .Y(n269), .A(B_not[23]) );
  inv02 U296 ( .Y(n270), .A(A[23]) );
  inv02 U297 ( .Y(n271), .A(carry_23_) );
  nor02 U298 ( .Y(n272), .A0(n269), .A1(n273) );
  nor02 U299 ( .Y(n274), .A0(n270), .A1(n275) );
  nor02 U300 ( .Y(n276), .A0(n271), .A1(n277) );
  nor02 U301 ( .Y(n278), .A0(n271), .A1(n279) );
  nor02 U302 ( .Y(n267), .A0(n280), .A1(n281) );
  nor02 U303 ( .Y(n282), .A0(n270), .A1(n271) );
  nor02 U304 ( .Y(n283), .A0(n269), .A1(n271) );
  nor02 U305 ( .Y(n284), .A0(n269), .A1(n270) );
  nor02 U306 ( .Y(n268), .A0(n284), .A1(n285) );
  nor02 U307 ( .Y(n286), .A0(A[23]), .A1(carry_23_) );
  inv01 U308 ( .Y(n273), .A(n286) );
  nor02 U309 ( .Y(n287), .A0(B_not[23]), .A1(carry_23_) );
  inv01 U310 ( .Y(n275), .A(n287) );
  nor02 U311 ( .Y(n288), .A0(B_not[23]), .A1(A[23]) );
  inv01 U312 ( .Y(n277), .A(n288) );
  nor02 U313 ( .Y(n289), .A0(n269), .A1(n270) );
  inv01 U314 ( .Y(n279), .A(n289) );
  nor02 U315 ( .Y(n290), .A0(n272), .A1(n274) );
  inv01 U316 ( .Y(n280), .A(n290) );
  nor02 U317 ( .Y(n291), .A0(n276), .A1(n278) );
  inv01 U318 ( .Y(n281), .A(n291) );
  nor02 U319 ( .Y(n292), .A0(n282), .A1(n283) );
  inv01 U320 ( .Y(n285), .A(n292) );
  inv01 U321 ( .Y(DIFF[41]), .A(n293) );
  inv02 U322 ( .Y(carry_42_), .A(n294) );
  inv02 U323 ( .Y(n295), .A(B_not[41]) );
  inv02 U324 ( .Y(n296), .A(A[41]) );
  inv02 U325 ( .Y(n297), .A(carry_41_) );
  nor02 U326 ( .Y(n298), .A0(n295), .A1(n299) );
  nor02 U327 ( .Y(n300), .A0(n296), .A1(n301) );
  nor02 U328 ( .Y(n302), .A0(n297), .A1(n303) );
  nor02 U329 ( .Y(n304), .A0(n297), .A1(n305) );
  nor02 U330 ( .Y(n293), .A0(n306), .A1(n307) );
  nor02 U331 ( .Y(n308), .A0(n296), .A1(n297) );
  nor02 U332 ( .Y(n309), .A0(n295), .A1(n297) );
  nor02 U333 ( .Y(n310), .A0(n295), .A1(n296) );
  nor02 U334 ( .Y(n294), .A0(n310), .A1(n311) );
  nor02 U335 ( .Y(n312), .A0(A[41]), .A1(carry_41_) );
  inv01 U336 ( .Y(n299), .A(n312) );
  nor02 U337 ( .Y(n313), .A0(B_not[41]), .A1(carry_41_) );
  inv01 U338 ( .Y(n301), .A(n313) );
  nor02 U339 ( .Y(n314), .A0(B_not[41]), .A1(A[41]) );
  inv01 U340 ( .Y(n303), .A(n314) );
  nor02 U341 ( .Y(n315), .A0(n295), .A1(n296) );
  inv01 U342 ( .Y(n305), .A(n315) );
  nor02 U343 ( .Y(n316), .A0(n298), .A1(n300) );
  inv01 U344 ( .Y(n306), .A(n316) );
  nor02 U345 ( .Y(n317), .A0(n302), .A1(n304) );
  inv01 U346 ( .Y(n307), .A(n317) );
  nor02 U347 ( .Y(n318), .A0(n308), .A1(n309) );
  inv01 U348 ( .Y(n311), .A(n318) );
  inv01 U349 ( .Y(DIFF[21]), .A(n319) );
  inv02 U350 ( .Y(carry_22_), .A(n320) );
  inv02 U351 ( .Y(n321), .A(B_not[21]) );
  inv02 U352 ( .Y(n322), .A(A[21]) );
  inv02 U353 ( .Y(n323), .A(carry_21_) );
  nor02 U354 ( .Y(n324), .A0(n321), .A1(n325) );
  nor02 U355 ( .Y(n326), .A0(n322), .A1(n327) );
  nor02 U356 ( .Y(n328), .A0(n323), .A1(n329) );
  nor02 U357 ( .Y(n330), .A0(n323), .A1(n331) );
  nor02 U358 ( .Y(n319), .A0(n332), .A1(n333) );
  nor02 U359 ( .Y(n334), .A0(n322), .A1(n323) );
  nor02 U360 ( .Y(n335), .A0(n321), .A1(n323) );
  nor02 U361 ( .Y(n336), .A0(n321), .A1(n322) );
  nor02 U362 ( .Y(n320), .A0(n336), .A1(n337) );
  nor02 U363 ( .Y(n338), .A0(A[21]), .A1(carry_21_) );
  inv01 U364 ( .Y(n325), .A(n338) );
  nor02 U365 ( .Y(n339), .A0(B_not[21]), .A1(carry_21_) );
  inv01 U366 ( .Y(n327), .A(n339) );
  nor02 U367 ( .Y(n340), .A0(B_not[21]), .A1(A[21]) );
  inv01 U368 ( .Y(n329), .A(n340) );
  nor02 U369 ( .Y(n341), .A0(n321), .A1(n322) );
  inv01 U370 ( .Y(n331), .A(n341) );
  nor02 U371 ( .Y(n342), .A0(n324), .A1(n326) );
  inv01 U372 ( .Y(n332), .A(n342) );
  nor02 U373 ( .Y(n343), .A0(n328), .A1(n330) );
  inv01 U374 ( .Y(n333), .A(n343) );
  nor02 U375 ( .Y(n344), .A0(n334), .A1(n335) );
  inv01 U376 ( .Y(n337), .A(n344) );
  inv02 U377 ( .Y(B_not[23]), .A(B[23]) );
  inv02 U378 ( .Y(B_not[21]), .A(B[21]) );
  inv01 U379 ( .Y(DIFF[24]), .A(n345) );
  inv02 U380 ( .Y(carry_25_), .A(n346) );
  inv02 U381 ( .Y(n347), .A(B_not[24]) );
  inv02 U382 ( .Y(n348), .A(A[24]) );
  inv02 U383 ( .Y(n349), .A(carry_24_) );
  nor02 U384 ( .Y(n350), .A0(n347), .A1(n351) );
  nor02 U385 ( .Y(n352), .A0(n348), .A1(n353) );
  nor02 U386 ( .Y(n354), .A0(n349), .A1(n355) );
  nor02 U387 ( .Y(n356), .A0(n349), .A1(n357) );
  nor02 U388 ( .Y(n345), .A0(n358), .A1(n359) );
  nor02 U389 ( .Y(n360), .A0(n348), .A1(n349) );
  nor02 U390 ( .Y(n361), .A0(n347), .A1(n349) );
  nor02 U391 ( .Y(n362), .A0(n347), .A1(n348) );
  nor02 U392 ( .Y(n346), .A0(n362), .A1(n363) );
  nor02 U393 ( .Y(n364), .A0(A[24]), .A1(carry_24_) );
  inv01 U394 ( .Y(n351), .A(n364) );
  nor02 U395 ( .Y(n365), .A0(B_not[24]), .A1(carry_24_) );
  inv01 U396 ( .Y(n353), .A(n365) );
  nor02 U397 ( .Y(n366), .A0(B_not[24]), .A1(A[24]) );
  inv01 U398 ( .Y(n355), .A(n366) );
  nor02 U399 ( .Y(n367), .A0(n347), .A1(n348) );
  inv01 U400 ( .Y(n357), .A(n367) );
  nor02 U401 ( .Y(n368), .A0(n350), .A1(n352) );
  inv01 U402 ( .Y(n358), .A(n368) );
  nor02 U403 ( .Y(n369), .A0(n354), .A1(n356) );
  inv01 U404 ( .Y(n359), .A(n369) );
  nor02 U405 ( .Y(n370), .A0(n360), .A1(n361) );
  inv01 U406 ( .Y(n363), .A(n370) );
  inv01 U407 ( .Y(DIFF[40]), .A(n371) );
  inv02 U408 ( .Y(carry_41_), .A(n372) );
  inv02 U409 ( .Y(n373), .A(B_not[40]) );
  inv02 U410 ( .Y(n374), .A(A[40]) );
  inv02 U411 ( .Y(n375), .A(carry_40_) );
  nor02 U412 ( .Y(n376), .A0(n373), .A1(n377) );
  nor02 U413 ( .Y(n378), .A0(n374), .A1(n379) );
  nor02 U414 ( .Y(n380), .A0(n375), .A1(n381) );
  nor02 U415 ( .Y(n382), .A0(n375), .A1(n383) );
  nor02 U416 ( .Y(n371), .A0(n384), .A1(n385) );
  nor02 U417 ( .Y(n386), .A0(n374), .A1(n375) );
  nor02 U418 ( .Y(n387), .A0(n373), .A1(n375) );
  nor02 U419 ( .Y(n388), .A0(n373), .A1(n374) );
  nor02 U420 ( .Y(n372), .A0(n388), .A1(n389) );
  nor02 U421 ( .Y(n390), .A0(A[40]), .A1(carry_40_) );
  inv01 U422 ( .Y(n377), .A(n390) );
  nor02 U423 ( .Y(n391), .A0(B_not[40]), .A1(carry_40_) );
  inv01 U424 ( .Y(n379), .A(n391) );
  nor02 U425 ( .Y(n392), .A0(B_not[40]), .A1(A[40]) );
  inv01 U426 ( .Y(n381), .A(n392) );
  nor02 U427 ( .Y(n393), .A0(n373), .A1(n374) );
  inv01 U428 ( .Y(n383), .A(n393) );
  nor02 U429 ( .Y(n394), .A0(n376), .A1(n378) );
  inv01 U430 ( .Y(n384), .A(n394) );
  nor02 U431 ( .Y(n395), .A0(n380), .A1(n382) );
  inv01 U432 ( .Y(n385), .A(n395) );
  nor02 U433 ( .Y(n396), .A0(n386), .A1(n387) );
  inv01 U434 ( .Y(n389), .A(n396) );
  inv01 U435 ( .Y(DIFF[20]), .A(n397) );
  inv02 U436 ( .Y(carry_21_), .A(n398) );
  inv02 U437 ( .Y(n399), .A(B_not[20]) );
  inv02 U438 ( .Y(n400), .A(A[20]) );
  inv02 U439 ( .Y(n401), .A(carry_20_) );
  nor02 U440 ( .Y(n402), .A0(n399), .A1(n403) );
  nor02 U441 ( .Y(n404), .A0(n400), .A1(n405) );
  nor02 U442 ( .Y(n406), .A0(n401), .A1(n407) );
  nor02 U443 ( .Y(n408), .A0(n401), .A1(n409) );
  nor02 U444 ( .Y(n397), .A0(n410), .A1(n411) );
  nor02 U445 ( .Y(n412), .A0(n400), .A1(n401) );
  nor02 U446 ( .Y(n413), .A0(n399), .A1(n401) );
  nor02 U447 ( .Y(n414), .A0(n399), .A1(n400) );
  nor02 U448 ( .Y(n398), .A0(n414), .A1(n415) );
  nor02 U449 ( .Y(n416), .A0(A[20]), .A1(carry_20_) );
  inv01 U450 ( .Y(n403), .A(n416) );
  nor02 U451 ( .Y(n417), .A0(B_not[20]), .A1(carry_20_) );
  inv01 U452 ( .Y(n405), .A(n417) );
  nor02 U453 ( .Y(n418), .A0(B_not[20]), .A1(A[20]) );
  inv01 U454 ( .Y(n407), .A(n418) );
  nor02 U455 ( .Y(n419), .A0(n399), .A1(n400) );
  inv01 U456 ( .Y(n409), .A(n419) );
  nor02 U457 ( .Y(n420), .A0(n402), .A1(n404) );
  inv01 U458 ( .Y(n410), .A(n420) );
  nor02 U459 ( .Y(n421), .A0(n406), .A1(n408) );
  inv01 U460 ( .Y(n411), .A(n421) );
  nor02 U461 ( .Y(n422), .A0(n412), .A1(n413) );
  inv01 U462 ( .Y(n415), .A(n422) );
  inv02 U463 ( .Y(B_not[24]), .A(n1313) );
  inv01 U464 ( .Y(DIFF[25]), .A(n423) );
  inv02 U465 ( .Y(carry_26_), .A(n424) );
  inv02 U466 ( .Y(n425), .A(B_not[25]) );
  inv02 U467 ( .Y(n426), .A(A[25]) );
  inv02 U468 ( .Y(n427), .A(carry_25_) );
  nor02 U469 ( .Y(n428), .A0(n425), .A1(n429) );
  nor02 U470 ( .Y(n430), .A0(n426), .A1(n431) );
  nor02 U471 ( .Y(n432), .A0(n427), .A1(n433) );
  nor02 U472 ( .Y(n434), .A0(n427), .A1(n435) );
  nor02 U473 ( .Y(n423), .A0(n436), .A1(n437) );
  nor02 U474 ( .Y(n438), .A0(n426), .A1(n427) );
  nor02 U475 ( .Y(n439), .A0(n425), .A1(n427) );
  nor02 U476 ( .Y(n440), .A0(n425), .A1(n426) );
  nor02 U477 ( .Y(n424), .A0(n440), .A1(n441) );
  nor02 U478 ( .Y(n442), .A0(A[25]), .A1(carry_25_) );
  inv01 U479 ( .Y(n429), .A(n442) );
  nor02 U480 ( .Y(n443), .A0(B_not[25]), .A1(carry_25_) );
  inv01 U481 ( .Y(n431), .A(n443) );
  nor02 U482 ( .Y(n444), .A0(B_not[25]), .A1(A[25]) );
  inv01 U483 ( .Y(n433), .A(n444) );
  nor02 U484 ( .Y(n445), .A0(n425), .A1(n426) );
  inv01 U485 ( .Y(n435), .A(n445) );
  nor02 U486 ( .Y(n446), .A0(n428), .A1(n430) );
  inv01 U487 ( .Y(n436), .A(n446) );
  nor02 U488 ( .Y(n447), .A0(n432), .A1(n434) );
  inv01 U489 ( .Y(n437), .A(n447) );
  nor02 U490 ( .Y(n448), .A0(n438), .A1(n439) );
  inv01 U491 ( .Y(n441), .A(n448) );
  inv01 U492 ( .Y(DIFF[19]), .A(n449) );
  inv02 U493 ( .Y(carry_20_), .A(n450) );
  inv02 U494 ( .Y(n451), .A(B_not[19]) );
  inv02 U495 ( .Y(n452), .A(A[19]) );
  inv02 U496 ( .Y(n453), .A(carry_19_) );
  nor02 U497 ( .Y(n454), .A0(n451), .A1(n455) );
  nor02 U498 ( .Y(n456), .A0(n452), .A1(n457) );
  nor02 U499 ( .Y(n458), .A0(n453), .A1(n459) );
  nor02 U500 ( .Y(n460), .A0(n453), .A1(n461) );
  nor02 U501 ( .Y(n449), .A0(n462), .A1(n463) );
  nor02 U502 ( .Y(n464), .A0(n452), .A1(n453) );
  nor02 U503 ( .Y(n465), .A0(n451), .A1(n453) );
  nor02 U504 ( .Y(n466), .A0(n451), .A1(n452) );
  nor02 U505 ( .Y(n450), .A0(n466), .A1(n467) );
  nor02 U506 ( .Y(n468), .A0(A[19]), .A1(carry_19_) );
  inv01 U507 ( .Y(n455), .A(n468) );
  nor02 U508 ( .Y(n469), .A0(B_not[19]), .A1(carry_19_) );
  inv01 U509 ( .Y(n457), .A(n469) );
  nor02 U510 ( .Y(n470), .A0(B_not[19]), .A1(A[19]) );
  inv01 U511 ( .Y(n459), .A(n470) );
  nor02 U512 ( .Y(n471), .A0(n451), .A1(n452) );
  inv01 U513 ( .Y(n461), .A(n471) );
  nor02 U514 ( .Y(n472), .A0(n454), .A1(n456) );
  inv01 U515 ( .Y(n462), .A(n472) );
  nor02 U516 ( .Y(n473), .A0(n458), .A1(n460) );
  inv01 U517 ( .Y(n463), .A(n473) );
  nor02 U518 ( .Y(n474), .A0(n464), .A1(n465) );
  inv01 U519 ( .Y(n467), .A(n474) );
  inv01 U520 ( .Y(DIFF[39]), .A(n475) );
  inv02 U521 ( .Y(carry_40_), .A(n476) );
  inv02 U522 ( .Y(n477), .A(B_not[39]) );
  inv02 U523 ( .Y(n478), .A(A[39]) );
  inv02 U524 ( .Y(n479), .A(carry_39_) );
  nor02 U525 ( .Y(n480), .A0(n477), .A1(n481) );
  nor02 U526 ( .Y(n482), .A0(n478), .A1(n483) );
  nor02 U527 ( .Y(n484), .A0(n479), .A1(n485) );
  nor02 U528 ( .Y(n486), .A0(n479), .A1(n487) );
  nor02 U529 ( .Y(n475), .A0(n488), .A1(n489) );
  nor02 U530 ( .Y(n490), .A0(n478), .A1(n479) );
  nor02 U531 ( .Y(n491), .A0(n477), .A1(n479) );
  nor02 U532 ( .Y(n492), .A0(n477), .A1(n478) );
  nor02 U533 ( .Y(n476), .A0(n492), .A1(n493) );
  nor02 U534 ( .Y(n494), .A0(A[39]), .A1(carry_39_) );
  inv01 U535 ( .Y(n481), .A(n494) );
  nor02 U536 ( .Y(n495), .A0(B_not[39]), .A1(carry_39_) );
  inv01 U537 ( .Y(n483), .A(n495) );
  nor02 U538 ( .Y(n496), .A0(B_not[39]), .A1(A[39]) );
  inv01 U539 ( .Y(n485), .A(n496) );
  nor02 U540 ( .Y(n497), .A0(n477), .A1(n478) );
  inv01 U541 ( .Y(n487), .A(n497) );
  nor02 U542 ( .Y(n498), .A0(n480), .A1(n482) );
  inv01 U543 ( .Y(n488), .A(n498) );
  nor02 U544 ( .Y(n499), .A0(n484), .A1(n486) );
  inv01 U545 ( .Y(n489), .A(n499) );
  nor02 U546 ( .Y(n500), .A0(n490), .A1(n491) );
  inv01 U547 ( .Y(n493), .A(n500) );
  inv01 U548 ( .Y(DIFF[26]), .A(n501) );
  inv02 U549 ( .Y(carry_27_), .A(n502) );
  inv02 U550 ( .Y(n503), .A(B_not[26]) );
  inv02 U551 ( .Y(n504), .A(A[26]) );
  inv02 U552 ( .Y(n505), .A(carry_26_) );
  nor02 U553 ( .Y(n506), .A0(n503), .A1(n507) );
  nor02 U554 ( .Y(n508), .A0(n504), .A1(n509) );
  nor02 U555 ( .Y(n510), .A0(n505), .A1(n511) );
  nor02 U556 ( .Y(n512), .A0(n505), .A1(n513) );
  nor02 U557 ( .Y(n501), .A0(n514), .A1(n515) );
  nor02 U558 ( .Y(n516), .A0(n504), .A1(n505) );
  nor02 U559 ( .Y(n517), .A0(n503), .A1(n505) );
  nor02 U560 ( .Y(n518), .A0(n503), .A1(n504) );
  nor02 U561 ( .Y(n502), .A0(n518), .A1(n519) );
  nor02 U562 ( .Y(n520), .A0(A[26]), .A1(carry_26_) );
  inv01 U563 ( .Y(n507), .A(n520) );
  nor02 U564 ( .Y(n521), .A0(B_not[26]), .A1(carry_26_) );
  inv01 U565 ( .Y(n509), .A(n521) );
  nor02 U566 ( .Y(n522), .A0(B_not[26]), .A1(A[26]) );
  inv01 U567 ( .Y(n511), .A(n522) );
  nor02 U568 ( .Y(n523), .A0(n503), .A1(n504) );
  inv01 U569 ( .Y(n513), .A(n523) );
  nor02 U570 ( .Y(n524), .A0(n506), .A1(n508) );
  inv01 U571 ( .Y(n514), .A(n524) );
  nor02 U572 ( .Y(n525), .A0(n510), .A1(n512) );
  inv01 U573 ( .Y(n515), .A(n525) );
  nor02 U574 ( .Y(n526), .A0(n516), .A1(n517) );
  inv01 U575 ( .Y(n519), .A(n526) );
  inv01 U576 ( .Y(DIFF[18]), .A(n527) );
  inv02 U577 ( .Y(carry_19_), .A(n528) );
  inv02 U578 ( .Y(n529), .A(B_not[18]) );
  inv02 U579 ( .Y(n530), .A(A[18]) );
  inv02 U580 ( .Y(n531), .A(carry_18_) );
  nor02 U581 ( .Y(n532), .A0(n529), .A1(n533) );
  nor02 U582 ( .Y(n534), .A0(n530), .A1(n535) );
  nor02 U583 ( .Y(n536), .A0(n531), .A1(n537) );
  nor02 U584 ( .Y(n538), .A0(n531), .A1(n539) );
  nor02 U585 ( .Y(n527), .A0(n540), .A1(n541) );
  nor02 U586 ( .Y(n542), .A0(n530), .A1(n531) );
  nor02 U587 ( .Y(n543), .A0(n529), .A1(n531) );
  nor02 U588 ( .Y(n544), .A0(n529), .A1(n530) );
  nor02 U589 ( .Y(n528), .A0(n544), .A1(n545) );
  nor02 U590 ( .Y(n546), .A0(A[18]), .A1(carry_18_) );
  inv01 U591 ( .Y(n533), .A(n546) );
  nor02 U592 ( .Y(n547), .A0(B_not[18]), .A1(carry_18_) );
  inv01 U593 ( .Y(n535), .A(n547) );
  nor02 U594 ( .Y(n548), .A0(B_not[18]), .A1(A[18]) );
  inv01 U595 ( .Y(n537), .A(n548) );
  nor02 U596 ( .Y(n549), .A0(n529), .A1(n530) );
  inv01 U597 ( .Y(n539), .A(n549) );
  nor02 U598 ( .Y(n550), .A0(n532), .A1(n534) );
  inv01 U599 ( .Y(n540), .A(n550) );
  nor02 U600 ( .Y(n551), .A0(n536), .A1(n538) );
  inv01 U601 ( .Y(n541), .A(n551) );
  nor02 U602 ( .Y(n552), .A0(n542), .A1(n543) );
  inv01 U603 ( .Y(n545), .A(n552) );
  inv01 U604 ( .Y(DIFF[38]), .A(n553) );
  inv02 U605 ( .Y(carry_39_), .A(n554) );
  inv02 U606 ( .Y(n555), .A(B_not[38]) );
  inv02 U607 ( .Y(n556), .A(A[38]) );
  inv02 U608 ( .Y(n557), .A(carry_38_) );
  nor02 U609 ( .Y(n558), .A0(n555), .A1(n559) );
  nor02 U610 ( .Y(n560), .A0(n556), .A1(n561) );
  nor02 U611 ( .Y(n562), .A0(n557), .A1(n563) );
  nor02 U612 ( .Y(n564), .A0(n557), .A1(n565) );
  nor02 U613 ( .Y(n553), .A0(n566), .A1(n567) );
  nor02 U614 ( .Y(n568), .A0(n556), .A1(n557) );
  nor02 U615 ( .Y(n569), .A0(n555), .A1(n557) );
  nor02 U616 ( .Y(n570), .A0(n555), .A1(n556) );
  nor02 U617 ( .Y(n554), .A0(n570), .A1(n571) );
  nor02 U618 ( .Y(n572), .A0(A[38]), .A1(carry_38_) );
  inv01 U619 ( .Y(n559), .A(n572) );
  nor02 U620 ( .Y(n573), .A0(B_not[38]), .A1(carry_38_) );
  inv01 U621 ( .Y(n561), .A(n573) );
  nor02 U622 ( .Y(n574), .A0(B_not[38]), .A1(A[38]) );
  inv01 U623 ( .Y(n563), .A(n574) );
  nor02 U624 ( .Y(n575), .A0(n555), .A1(n556) );
  inv01 U625 ( .Y(n565), .A(n575) );
  nor02 U626 ( .Y(n576), .A0(n558), .A1(n560) );
  inv01 U627 ( .Y(n566), .A(n576) );
  nor02 U628 ( .Y(n577), .A0(n562), .A1(n564) );
  inv01 U629 ( .Y(n567), .A(n577) );
  nor02 U630 ( .Y(n578), .A0(n568), .A1(n569) );
  inv01 U631 ( .Y(n571), .A(n578) );
  inv01 U632 ( .Y(DIFF[27]), .A(n579) );
  inv02 U633 ( .Y(carry_28_), .A(n580) );
  inv02 U634 ( .Y(n581), .A(B_not[27]) );
  inv02 U635 ( .Y(n582), .A(A[27]) );
  inv02 U636 ( .Y(n583), .A(carry_27_) );
  nor02 U637 ( .Y(n584), .A0(n581), .A1(n585) );
  nor02 U638 ( .Y(n586), .A0(n582), .A1(n587) );
  nor02 U639 ( .Y(n588), .A0(n583), .A1(n589) );
  nor02 U640 ( .Y(n590), .A0(n583), .A1(n591) );
  nor02 U641 ( .Y(n579), .A0(n592), .A1(n593) );
  nor02 U642 ( .Y(n594), .A0(n582), .A1(n583) );
  nor02 U643 ( .Y(n595), .A0(n581), .A1(n583) );
  nor02 U644 ( .Y(n596), .A0(n581), .A1(n582) );
  nor02 U645 ( .Y(n580), .A0(n596), .A1(n597) );
  nor02 U646 ( .Y(n598), .A0(A[27]), .A1(carry_27_) );
  inv01 U647 ( .Y(n585), .A(n598) );
  nor02 U648 ( .Y(n599), .A0(B_not[27]), .A1(carry_27_) );
  inv01 U649 ( .Y(n587), .A(n599) );
  nor02 U650 ( .Y(n600), .A0(B_not[27]), .A1(A[27]) );
  inv01 U651 ( .Y(n589), .A(n600) );
  nor02 U652 ( .Y(n601), .A0(n581), .A1(n582) );
  inv01 U653 ( .Y(n591), .A(n601) );
  nor02 U654 ( .Y(n602), .A0(n584), .A1(n586) );
  inv01 U655 ( .Y(n592), .A(n602) );
  nor02 U656 ( .Y(n603), .A0(n588), .A1(n590) );
  inv01 U657 ( .Y(n593), .A(n603) );
  nor02 U658 ( .Y(n604), .A0(n594), .A1(n595) );
  inv01 U659 ( .Y(n597), .A(n604) );
  inv01 U660 ( .Y(DIFF[37]), .A(n605) );
  inv02 U661 ( .Y(carry_38_), .A(n606) );
  inv02 U662 ( .Y(n607), .A(B_not[37]) );
  inv02 U663 ( .Y(n608), .A(A[37]) );
  inv02 U664 ( .Y(n609), .A(carry_37_) );
  nor02 U665 ( .Y(n610), .A0(n607), .A1(n611) );
  nor02 U666 ( .Y(n612), .A0(n608), .A1(n613) );
  nor02 U667 ( .Y(n614), .A0(n609), .A1(n615) );
  nor02 U668 ( .Y(n616), .A0(n609), .A1(n617) );
  nor02 U669 ( .Y(n605), .A0(n618), .A1(n619) );
  nor02 U670 ( .Y(n620), .A0(n608), .A1(n609) );
  nor02 U671 ( .Y(n621), .A0(n607), .A1(n609) );
  nor02 U672 ( .Y(n622), .A0(n607), .A1(n608) );
  nor02 U673 ( .Y(n606), .A0(n622), .A1(n623) );
  nor02 U674 ( .Y(n624), .A0(A[37]), .A1(carry_37_) );
  inv01 U675 ( .Y(n611), .A(n624) );
  nor02 U676 ( .Y(n625), .A0(B_not[37]), .A1(carry_37_) );
  inv01 U677 ( .Y(n613), .A(n625) );
  nor02 U678 ( .Y(n626), .A0(B_not[37]), .A1(A[37]) );
  inv01 U679 ( .Y(n615), .A(n626) );
  nor02 U680 ( .Y(n627), .A0(n607), .A1(n608) );
  inv01 U681 ( .Y(n617), .A(n627) );
  nor02 U682 ( .Y(n628), .A0(n610), .A1(n612) );
  inv01 U683 ( .Y(n618), .A(n628) );
  nor02 U684 ( .Y(n629), .A0(n614), .A1(n616) );
  inv01 U685 ( .Y(n619), .A(n629) );
  nor02 U686 ( .Y(n630), .A0(n620), .A1(n621) );
  inv01 U687 ( .Y(n623), .A(n630) );
  inv01 U688 ( .Y(DIFF[17]), .A(n631) );
  inv02 U689 ( .Y(carry_18_), .A(n632) );
  inv02 U690 ( .Y(n633), .A(B_not[17]) );
  inv02 U691 ( .Y(n634), .A(A[17]) );
  inv02 U692 ( .Y(n635), .A(carry_17_) );
  nor02 U693 ( .Y(n636), .A0(n633), .A1(n637) );
  nor02 U694 ( .Y(n638), .A0(n634), .A1(n639) );
  nor02 U695 ( .Y(n640), .A0(n635), .A1(n641) );
  nor02 U696 ( .Y(n642), .A0(n635), .A1(n643) );
  nor02 U697 ( .Y(n631), .A0(n644), .A1(n645) );
  nor02 U698 ( .Y(n646), .A0(n634), .A1(n635) );
  nor02 U699 ( .Y(n647), .A0(n633), .A1(n635) );
  nor02 U700 ( .Y(n648), .A0(n633), .A1(n634) );
  nor02 U701 ( .Y(n632), .A0(n648), .A1(n649) );
  nor02 U702 ( .Y(n650), .A0(A[17]), .A1(carry_17_) );
  inv01 U703 ( .Y(n637), .A(n650) );
  nor02 U704 ( .Y(n651), .A0(B_not[17]), .A1(carry_17_) );
  inv01 U705 ( .Y(n639), .A(n651) );
  nor02 U706 ( .Y(n652), .A0(B_not[17]), .A1(A[17]) );
  inv01 U707 ( .Y(n641), .A(n652) );
  nor02 U708 ( .Y(n653), .A0(n633), .A1(n634) );
  inv01 U709 ( .Y(n643), .A(n653) );
  nor02 U710 ( .Y(n654), .A0(n636), .A1(n638) );
  inv01 U711 ( .Y(n644), .A(n654) );
  nor02 U712 ( .Y(n655), .A0(n640), .A1(n642) );
  inv01 U713 ( .Y(n645), .A(n655) );
  nor02 U714 ( .Y(n656), .A0(n646), .A1(n647) );
  inv01 U715 ( .Y(n649), .A(n656) );
  inv01 U716 ( .Y(DIFF[28]), .A(n657) );
  inv02 U717 ( .Y(carry_29_), .A(n658) );
  inv02 U718 ( .Y(n659), .A(B_not[28]) );
  inv02 U719 ( .Y(n660), .A(A[28]) );
  inv02 U720 ( .Y(n661), .A(carry_28_) );
  nor02 U721 ( .Y(n662), .A0(n659), .A1(n663) );
  nor02 U722 ( .Y(n664), .A0(n660), .A1(n665) );
  nor02 U723 ( .Y(n666), .A0(n661), .A1(n667) );
  nor02 U724 ( .Y(n668), .A0(n661), .A1(n669) );
  nor02 U725 ( .Y(n657), .A0(n670), .A1(n671) );
  nor02 U726 ( .Y(n672), .A0(n660), .A1(n661) );
  nor02 U727 ( .Y(n673), .A0(n659), .A1(n661) );
  nor02 U728 ( .Y(n674), .A0(n659), .A1(n660) );
  nor02 U729 ( .Y(n658), .A0(n674), .A1(n675) );
  nor02 U730 ( .Y(n676), .A0(A[28]), .A1(carry_28_) );
  inv01 U731 ( .Y(n663), .A(n676) );
  nor02 U732 ( .Y(n677), .A0(B_not[28]), .A1(carry_28_) );
  inv01 U733 ( .Y(n665), .A(n677) );
  nor02 U734 ( .Y(n678), .A0(B_not[28]), .A1(A[28]) );
  inv01 U735 ( .Y(n667), .A(n678) );
  nor02 U736 ( .Y(n679), .A0(n659), .A1(n660) );
  inv01 U737 ( .Y(n669), .A(n679) );
  nor02 U738 ( .Y(n680), .A0(n662), .A1(n664) );
  inv01 U739 ( .Y(n670), .A(n680) );
  nor02 U740 ( .Y(n681), .A0(n666), .A1(n668) );
  inv01 U741 ( .Y(n671), .A(n681) );
  nor02 U742 ( .Y(n682), .A0(n672), .A1(n673) );
  inv01 U743 ( .Y(n675), .A(n682) );
  inv01 U744 ( .Y(DIFF[36]), .A(n683) );
  inv02 U745 ( .Y(carry_37_), .A(n684) );
  inv02 U746 ( .Y(n685), .A(B_not[36]) );
  inv02 U747 ( .Y(n686), .A(A[36]) );
  inv02 U748 ( .Y(n687), .A(carry_36_) );
  nor02 U749 ( .Y(n688), .A0(n685), .A1(n689) );
  nor02 U750 ( .Y(n690), .A0(n686), .A1(n691) );
  nor02 U751 ( .Y(n692), .A0(n687), .A1(n693) );
  nor02 U752 ( .Y(n694), .A0(n687), .A1(n695) );
  nor02 U753 ( .Y(n683), .A0(n696), .A1(n697) );
  nor02 U754 ( .Y(n698), .A0(n686), .A1(n687) );
  nor02 U755 ( .Y(n699), .A0(n685), .A1(n687) );
  nor02 U756 ( .Y(n700), .A0(n685), .A1(n686) );
  nor02 U757 ( .Y(n684), .A0(n700), .A1(n701) );
  nor02 U758 ( .Y(n702), .A0(A[36]), .A1(carry_36_) );
  inv01 U759 ( .Y(n689), .A(n702) );
  nor02 U760 ( .Y(n703), .A0(B_not[36]), .A1(carry_36_) );
  inv01 U761 ( .Y(n691), .A(n703) );
  nor02 U762 ( .Y(n704), .A0(B_not[36]), .A1(A[36]) );
  inv01 U763 ( .Y(n693), .A(n704) );
  nor02 U764 ( .Y(n705), .A0(n685), .A1(n686) );
  inv01 U765 ( .Y(n695), .A(n705) );
  nor02 U766 ( .Y(n706), .A0(n688), .A1(n690) );
  inv01 U767 ( .Y(n696), .A(n706) );
  nor02 U768 ( .Y(n707), .A0(n692), .A1(n694) );
  inv01 U769 ( .Y(n697), .A(n707) );
  nor02 U770 ( .Y(n708), .A0(n698), .A1(n699) );
  inv01 U771 ( .Y(n701), .A(n708) );
  inv01 U772 ( .Y(DIFF[16]), .A(n709) );
  inv02 U773 ( .Y(carry_17_), .A(n710) );
  inv02 U774 ( .Y(n711), .A(B_not[16]) );
  inv02 U775 ( .Y(n712), .A(A[16]) );
  inv02 U776 ( .Y(n713), .A(carry_16_) );
  nor02 U777 ( .Y(n714), .A0(n711), .A1(n715) );
  nor02 U778 ( .Y(n716), .A0(n712), .A1(n717) );
  nor02 U779 ( .Y(n718), .A0(n713), .A1(n719) );
  nor02 U780 ( .Y(n720), .A0(n713), .A1(n721) );
  nor02 U781 ( .Y(n709), .A0(n722), .A1(n723) );
  nor02 U782 ( .Y(n724), .A0(n712), .A1(n713) );
  nor02 U783 ( .Y(n725), .A0(n711), .A1(n713) );
  nor02 U784 ( .Y(n726), .A0(n711), .A1(n712) );
  nor02 U785 ( .Y(n710), .A0(n726), .A1(n727) );
  nor02 U786 ( .Y(n728), .A0(A[16]), .A1(carry_16_) );
  inv01 U787 ( .Y(n715), .A(n728) );
  nor02 U788 ( .Y(n729), .A0(B_not[16]), .A1(carry_16_) );
  inv01 U789 ( .Y(n717), .A(n729) );
  nor02 U790 ( .Y(n730), .A0(B_not[16]), .A1(A[16]) );
  inv01 U791 ( .Y(n719), .A(n730) );
  nor02 U792 ( .Y(n731), .A0(n711), .A1(n712) );
  inv01 U793 ( .Y(n721), .A(n731) );
  nor02 U794 ( .Y(n732), .A0(n714), .A1(n716) );
  inv01 U795 ( .Y(n722), .A(n732) );
  nor02 U796 ( .Y(n733), .A0(n718), .A1(n720) );
  inv01 U797 ( .Y(n723), .A(n733) );
  nor02 U798 ( .Y(n734), .A0(n724), .A1(n725) );
  inv01 U799 ( .Y(n727), .A(n734) );
  inv01 U800 ( .Y(DIFF[29]), .A(n735) );
  inv02 U801 ( .Y(carry_30_), .A(n736) );
  inv02 U802 ( .Y(n737), .A(B_not[29]) );
  inv02 U803 ( .Y(n738), .A(A[29]) );
  inv02 U804 ( .Y(n739), .A(carry_29_) );
  nor02 U805 ( .Y(n740), .A0(n737), .A1(n741) );
  nor02 U806 ( .Y(n742), .A0(n738), .A1(n743) );
  nor02 U807 ( .Y(n744), .A0(n739), .A1(n745) );
  nor02 U808 ( .Y(n746), .A0(n739), .A1(n747) );
  nor02 U809 ( .Y(n735), .A0(n748), .A1(n749) );
  nor02 U810 ( .Y(n750), .A0(n738), .A1(n739) );
  nor02 U811 ( .Y(n751), .A0(n737), .A1(n739) );
  nor02 U812 ( .Y(n752), .A0(n737), .A1(n738) );
  nor02 U813 ( .Y(n736), .A0(n752), .A1(n753) );
  nor02 U814 ( .Y(n754), .A0(A[29]), .A1(carry_29_) );
  inv01 U815 ( .Y(n741), .A(n754) );
  nor02 U816 ( .Y(n755), .A0(B_not[29]), .A1(carry_29_) );
  inv01 U817 ( .Y(n743), .A(n755) );
  nor02 U818 ( .Y(n756), .A0(B_not[29]), .A1(A[29]) );
  inv01 U819 ( .Y(n745), .A(n756) );
  nor02 U820 ( .Y(n757), .A0(n737), .A1(n738) );
  inv01 U821 ( .Y(n747), .A(n757) );
  nor02 U822 ( .Y(n758), .A0(n740), .A1(n742) );
  inv01 U823 ( .Y(n748), .A(n758) );
  nor02 U824 ( .Y(n759), .A0(n744), .A1(n746) );
  inv01 U825 ( .Y(n749), .A(n759) );
  nor02 U826 ( .Y(n760), .A0(n750), .A1(n751) );
  inv01 U827 ( .Y(n753), .A(n760) );
  inv01 U828 ( .Y(DIFF[35]), .A(n761) );
  inv02 U829 ( .Y(carry_36_), .A(n762) );
  inv02 U830 ( .Y(n763), .A(B_not[35]) );
  inv02 U831 ( .Y(n764), .A(A[35]) );
  inv02 U832 ( .Y(n765), .A(carry_35_) );
  nor02 U833 ( .Y(n766), .A0(n763), .A1(n767) );
  nor02 U834 ( .Y(n768), .A0(n764), .A1(n769) );
  nor02 U835 ( .Y(n770), .A0(n765), .A1(n771) );
  nor02 U836 ( .Y(n772), .A0(n765), .A1(n773) );
  nor02 U837 ( .Y(n761), .A0(n774), .A1(n775) );
  nor02 U838 ( .Y(n776), .A0(n764), .A1(n765) );
  nor02 U839 ( .Y(n777), .A0(n763), .A1(n765) );
  nor02 U840 ( .Y(n778), .A0(n763), .A1(n764) );
  nor02 U841 ( .Y(n762), .A0(n778), .A1(n779) );
  nor02 U842 ( .Y(n780), .A0(A[35]), .A1(carry_35_) );
  inv01 U843 ( .Y(n767), .A(n780) );
  nor02 U844 ( .Y(n781), .A0(B_not[35]), .A1(carry_35_) );
  inv01 U845 ( .Y(n769), .A(n781) );
  nor02 U846 ( .Y(n782), .A0(B_not[35]), .A1(A[35]) );
  inv01 U847 ( .Y(n771), .A(n782) );
  nor02 U848 ( .Y(n783), .A0(n763), .A1(n764) );
  inv01 U849 ( .Y(n773), .A(n783) );
  nor02 U850 ( .Y(n784), .A0(n766), .A1(n768) );
  inv01 U851 ( .Y(n774), .A(n784) );
  nor02 U852 ( .Y(n785), .A0(n770), .A1(n772) );
  inv01 U853 ( .Y(n775), .A(n785) );
  nor02 U854 ( .Y(n786), .A0(n776), .A1(n777) );
  inv01 U855 ( .Y(n779), .A(n786) );
  inv01 U856 ( .Y(DIFF[15]), .A(n787) );
  inv02 U857 ( .Y(carry_16_), .A(n788) );
  inv02 U858 ( .Y(n789), .A(B_not[15]) );
  inv02 U859 ( .Y(n790), .A(A[15]) );
  inv02 U860 ( .Y(n791), .A(carry_15_) );
  nor02 U861 ( .Y(n792), .A0(n789), .A1(n793) );
  nor02 U862 ( .Y(n794), .A0(n790), .A1(n795) );
  nor02 U863 ( .Y(n796), .A0(n791), .A1(n797) );
  nor02 U864 ( .Y(n798), .A0(n791), .A1(n799) );
  nor02 U865 ( .Y(n787), .A0(n800), .A1(n801) );
  nor02 U866 ( .Y(n802), .A0(n790), .A1(n791) );
  nor02 U867 ( .Y(n803), .A0(n789), .A1(n791) );
  nor02 U868 ( .Y(n804), .A0(n789), .A1(n790) );
  nor02 U869 ( .Y(n788), .A0(n804), .A1(n805) );
  nor02 U870 ( .Y(n806), .A0(A[15]), .A1(carry_15_) );
  inv01 U871 ( .Y(n793), .A(n806) );
  nor02 U872 ( .Y(n807), .A0(B_not[15]), .A1(carry_15_) );
  inv01 U873 ( .Y(n795), .A(n807) );
  nor02 U874 ( .Y(n808), .A0(B_not[15]), .A1(A[15]) );
  inv01 U875 ( .Y(n797), .A(n808) );
  nor02 U876 ( .Y(n809), .A0(n789), .A1(n790) );
  inv01 U877 ( .Y(n799), .A(n809) );
  nor02 U878 ( .Y(n810), .A0(n792), .A1(n794) );
  inv01 U879 ( .Y(n800), .A(n810) );
  nor02 U880 ( .Y(n811), .A0(n796), .A1(n798) );
  inv01 U881 ( .Y(n801), .A(n811) );
  nor02 U882 ( .Y(n812), .A0(n802), .A1(n803) );
  inv01 U883 ( .Y(n805), .A(n812) );
  inv01 U884 ( .Y(DIFF[30]), .A(n813) );
  inv02 U885 ( .Y(carry_31_), .A(n814) );
  inv02 U886 ( .Y(n815), .A(B_not[30]) );
  inv02 U887 ( .Y(n816), .A(A[30]) );
  inv02 U888 ( .Y(n817), .A(carry_30_) );
  nor02 U889 ( .Y(n818), .A0(n815), .A1(n819) );
  nor02 U890 ( .Y(n820), .A0(n816), .A1(n821) );
  nor02 U891 ( .Y(n822), .A0(n817), .A1(n823) );
  nor02 U892 ( .Y(n824), .A0(n817), .A1(n825) );
  nor02 U893 ( .Y(n813), .A0(n826), .A1(n827) );
  nor02 U894 ( .Y(n828), .A0(n816), .A1(n817) );
  nor02 U895 ( .Y(n829), .A0(n815), .A1(n817) );
  nor02 U896 ( .Y(n830), .A0(n815), .A1(n816) );
  nor02 U897 ( .Y(n814), .A0(n830), .A1(n831) );
  nor02 U898 ( .Y(n832), .A0(A[30]), .A1(carry_30_) );
  inv01 U899 ( .Y(n819), .A(n832) );
  nor02 U900 ( .Y(n833), .A0(B_not[30]), .A1(carry_30_) );
  inv01 U901 ( .Y(n821), .A(n833) );
  nor02 U902 ( .Y(n834), .A0(B_not[30]), .A1(A[30]) );
  inv01 U903 ( .Y(n823), .A(n834) );
  nor02 U904 ( .Y(n835), .A0(n815), .A1(n816) );
  inv01 U905 ( .Y(n825), .A(n835) );
  nor02 U906 ( .Y(n836), .A0(n818), .A1(n820) );
  inv01 U907 ( .Y(n826), .A(n836) );
  nor02 U908 ( .Y(n837), .A0(n822), .A1(n824) );
  inv01 U909 ( .Y(n827), .A(n837) );
  nor02 U910 ( .Y(n838), .A0(n828), .A1(n829) );
  inv01 U911 ( .Y(n831), .A(n838) );
  inv01 U912 ( .Y(DIFF[14]), .A(n839) );
  inv02 U913 ( .Y(carry_15_), .A(n840) );
  inv02 U914 ( .Y(n841), .A(B_not[14]) );
  inv02 U915 ( .Y(n842), .A(A[14]) );
  inv02 U916 ( .Y(n843), .A(carry_14_) );
  nor02 U917 ( .Y(n844), .A0(n841), .A1(n845) );
  nor02 U918 ( .Y(n846), .A0(n842), .A1(n847) );
  nor02 U919 ( .Y(n848), .A0(n843), .A1(n849) );
  nor02 U920 ( .Y(n850), .A0(n843), .A1(n851) );
  nor02 U921 ( .Y(n839), .A0(n852), .A1(n853) );
  nor02 U922 ( .Y(n854), .A0(n842), .A1(n843) );
  nor02 U923 ( .Y(n855), .A0(n841), .A1(n843) );
  nor02 U924 ( .Y(n856), .A0(n841), .A1(n842) );
  nor02 U925 ( .Y(n840), .A0(n856), .A1(n857) );
  nor02 U926 ( .Y(n858), .A0(A[14]), .A1(carry_14_) );
  inv01 U927 ( .Y(n845), .A(n858) );
  nor02 U928 ( .Y(n859), .A0(B_not[14]), .A1(carry_14_) );
  inv01 U929 ( .Y(n847), .A(n859) );
  nor02 U930 ( .Y(n860), .A0(B_not[14]), .A1(A[14]) );
  inv01 U931 ( .Y(n849), .A(n860) );
  nor02 U932 ( .Y(n861), .A0(n841), .A1(n842) );
  inv01 U933 ( .Y(n851), .A(n861) );
  nor02 U934 ( .Y(n862), .A0(n844), .A1(n846) );
  inv01 U935 ( .Y(n852), .A(n862) );
  nor02 U936 ( .Y(n863), .A0(n848), .A1(n850) );
  inv01 U937 ( .Y(n853), .A(n863) );
  nor02 U938 ( .Y(n864), .A0(n854), .A1(n855) );
  inv01 U939 ( .Y(n857), .A(n864) );
  inv01 U940 ( .Y(DIFF[34]), .A(n865) );
  inv02 U941 ( .Y(carry_35_), .A(n866) );
  inv02 U942 ( .Y(n867), .A(B_not[34]) );
  inv02 U943 ( .Y(n868), .A(A[34]) );
  inv02 U944 ( .Y(n869), .A(carry_34_) );
  nor02 U945 ( .Y(n870), .A0(n867), .A1(n871) );
  nor02 U946 ( .Y(n872), .A0(n868), .A1(n873) );
  nor02 U947 ( .Y(n874), .A0(n869), .A1(n875) );
  nor02 U948 ( .Y(n876), .A0(n869), .A1(n877) );
  nor02 U949 ( .Y(n865), .A0(n878), .A1(n879) );
  nor02 U950 ( .Y(n880), .A0(n868), .A1(n869) );
  nor02 U951 ( .Y(n881), .A0(n867), .A1(n869) );
  nor02 U952 ( .Y(n882), .A0(n867), .A1(n868) );
  nor02 U953 ( .Y(n866), .A0(n882), .A1(n883) );
  nor02 U954 ( .Y(n884), .A0(A[34]), .A1(carry_34_) );
  inv01 U955 ( .Y(n871), .A(n884) );
  nor02 U956 ( .Y(n885), .A0(B_not[34]), .A1(carry_34_) );
  inv01 U957 ( .Y(n873), .A(n885) );
  nor02 U958 ( .Y(n886), .A0(B_not[34]), .A1(A[34]) );
  inv01 U959 ( .Y(n875), .A(n886) );
  nor02 U960 ( .Y(n887), .A0(n867), .A1(n868) );
  inv01 U961 ( .Y(n877), .A(n887) );
  nor02 U962 ( .Y(n888), .A0(n870), .A1(n872) );
  inv01 U963 ( .Y(n878), .A(n888) );
  nor02 U964 ( .Y(n889), .A0(n874), .A1(n876) );
  inv01 U965 ( .Y(n879), .A(n889) );
  nor02 U966 ( .Y(n890), .A0(n880), .A1(n881) );
  inv01 U967 ( .Y(n883), .A(n890) );
  inv02 U968 ( .Y(B_not[30]), .A(n1312) );
  inv02 U969 ( .Y(B_not[34]), .A(n1311) );
  inv01 U970 ( .Y(DIFF[31]), .A(n891) );
  inv02 U971 ( .Y(carry_32_), .A(n892) );
  inv02 U972 ( .Y(n893), .A(B_not[31]) );
  inv02 U973 ( .Y(n894), .A(A[31]) );
  inv02 U974 ( .Y(n895), .A(carry_31_) );
  nor02 U975 ( .Y(n896), .A0(n893), .A1(n897) );
  nor02 U976 ( .Y(n898), .A0(n894), .A1(n899) );
  nor02 U977 ( .Y(n900), .A0(n895), .A1(n901) );
  nor02 U978 ( .Y(n902), .A0(n895), .A1(n903) );
  nor02 U979 ( .Y(n891), .A0(n904), .A1(n905) );
  nor02 U980 ( .Y(n906), .A0(n894), .A1(n895) );
  nor02 U981 ( .Y(n907), .A0(n893), .A1(n895) );
  nor02 U982 ( .Y(n908), .A0(n893), .A1(n894) );
  nor02 U983 ( .Y(n892), .A0(n908), .A1(n909) );
  nor02 U984 ( .Y(n910), .A0(A[31]), .A1(carry_31_) );
  inv01 U985 ( .Y(n897), .A(n910) );
  nor02 U986 ( .Y(n911), .A0(B_not[31]), .A1(carry_31_) );
  inv01 U987 ( .Y(n899), .A(n911) );
  nor02 U988 ( .Y(n912), .A0(B_not[31]), .A1(A[31]) );
  inv01 U989 ( .Y(n901), .A(n912) );
  nor02 U990 ( .Y(n913), .A0(n893), .A1(n894) );
  inv01 U991 ( .Y(n903), .A(n913) );
  nor02 U992 ( .Y(n914), .A0(n896), .A1(n898) );
  inv01 U993 ( .Y(n904), .A(n914) );
  nor02 U994 ( .Y(n915), .A0(n900), .A1(n902) );
  inv01 U995 ( .Y(n905), .A(n915) );
  nor02 U996 ( .Y(n916), .A0(n906), .A1(n907) );
  inv01 U997 ( .Y(n909), .A(n916) );
  inv01 U998 ( .Y(DIFF[33]), .A(n917) );
  inv02 U999 ( .Y(carry_34_), .A(n918) );
  inv02 U1000 ( .Y(n919), .A(B_not[33]) );
  inv02 U1001 ( .Y(n920), .A(A[33]) );
  inv02 U1002 ( .Y(n921), .A(carry_33_) );
  nor02 U1003 ( .Y(n922), .A0(n919), .A1(n923) );
  nor02 U1004 ( .Y(n924), .A0(n920), .A1(n925) );
  nor02 U1005 ( .Y(n926), .A0(n921), .A1(n927) );
  nor02 U1006 ( .Y(n928), .A0(n921), .A1(n929) );
  nor02 U1007 ( .Y(n917), .A0(n930), .A1(n931) );
  nor02 U1008 ( .Y(n932), .A0(n920), .A1(n921) );
  nor02 U1009 ( .Y(n933), .A0(n919), .A1(n921) );
  nor02 U1010 ( .Y(n934), .A0(n919), .A1(n920) );
  nor02 U1011 ( .Y(n918), .A0(n934), .A1(n935) );
  nor02 U1012 ( .Y(n936), .A0(A[33]), .A1(carry_33_) );
  inv01 U1013 ( .Y(n923), .A(n936) );
  nor02 U1014 ( .Y(n937), .A0(B_not[33]), .A1(carry_33_) );
  inv01 U1015 ( .Y(n925), .A(n937) );
  nor02 U1016 ( .Y(n938), .A0(B_not[33]), .A1(A[33]) );
  inv01 U1017 ( .Y(n927), .A(n938) );
  nor02 U1018 ( .Y(n939), .A0(n919), .A1(n920) );
  inv01 U1019 ( .Y(n929), .A(n939) );
  nor02 U1020 ( .Y(n940), .A0(n922), .A1(n924) );
  inv01 U1021 ( .Y(n930), .A(n940) );
  nor02 U1022 ( .Y(n941), .A0(n926), .A1(n928) );
  inv01 U1023 ( .Y(n931), .A(n941) );
  nor02 U1024 ( .Y(n942), .A0(n932), .A1(n933) );
  inv01 U1025 ( .Y(n935), .A(n942) );
  inv01 U1026 ( .Y(DIFF[13]), .A(n943) );
  inv02 U1027 ( .Y(carry_14_), .A(n944) );
  inv02 U1028 ( .Y(n945), .A(B_not[13]) );
  inv02 U1029 ( .Y(n946), .A(A[13]) );
  inv02 U1030 ( .Y(n947), .A(carry_13_) );
  nor02 U1031 ( .Y(n948), .A0(n945), .A1(n949) );
  nor02 U1032 ( .Y(n950), .A0(n946), .A1(n951) );
  nor02 U1033 ( .Y(n952), .A0(n947), .A1(n953) );
  nor02 U1034 ( .Y(n954), .A0(n947), .A1(n955) );
  nor02 U1035 ( .Y(n943), .A0(n956), .A1(n957) );
  nor02 U1036 ( .Y(n958), .A0(n946), .A1(n947) );
  nor02 U1037 ( .Y(n959), .A0(n945), .A1(n947) );
  nor02 U1038 ( .Y(n960), .A0(n945), .A1(n946) );
  nor02 U1039 ( .Y(n944), .A0(n960), .A1(n961) );
  nor02 U1040 ( .Y(n962), .A0(A[13]), .A1(carry_13_) );
  inv01 U1041 ( .Y(n949), .A(n962) );
  nor02 U1042 ( .Y(n963), .A0(B_not[13]), .A1(carry_13_) );
  inv01 U1043 ( .Y(n951), .A(n963) );
  nor02 U1044 ( .Y(n964), .A0(B_not[13]), .A1(A[13]) );
  inv01 U1045 ( .Y(n953), .A(n964) );
  nor02 U1046 ( .Y(n965), .A0(n945), .A1(n946) );
  inv01 U1047 ( .Y(n955), .A(n965) );
  nor02 U1048 ( .Y(n966), .A0(n948), .A1(n950) );
  inv01 U1049 ( .Y(n956), .A(n966) );
  nor02 U1050 ( .Y(n967), .A0(n952), .A1(n954) );
  inv01 U1051 ( .Y(n957), .A(n967) );
  nor02 U1052 ( .Y(n968), .A0(n958), .A1(n959) );
  inv01 U1053 ( .Y(n961), .A(n968) );
  inv01 U1054 ( .Y(DIFF[32]), .A(n969) );
  inv02 U1055 ( .Y(carry_33_), .A(n970) );
  inv02 U1056 ( .Y(n971), .A(B_not[32]) );
  inv02 U1057 ( .Y(n972), .A(A[32]) );
  inv02 U1058 ( .Y(n973), .A(carry_32_) );
  nor02 U1059 ( .Y(n974), .A0(n971), .A1(n975) );
  nor02 U1060 ( .Y(n976), .A0(n972), .A1(n977) );
  nor02 U1061 ( .Y(n978), .A0(n973), .A1(n979) );
  nor02 U1062 ( .Y(n980), .A0(n973), .A1(n981) );
  nor02 U1063 ( .Y(n969), .A0(n982), .A1(n983) );
  nor02 U1064 ( .Y(n984), .A0(n972), .A1(n973) );
  nor02 U1065 ( .Y(n985), .A0(n971), .A1(n973) );
  nor02 U1066 ( .Y(n986), .A0(n971), .A1(n972) );
  nor02 U1067 ( .Y(n970), .A0(n986), .A1(n987) );
  nor02 U1068 ( .Y(n988), .A0(A[32]), .A1(carry_32_) );
  inv01 U1069 ( .Y(n975), .A(n988) );
  nor02 U1070 ( .Y(n989), .A0(B_not[32]), .A1(carry_32_) );
  inv01 U1071 ( .Y(n977), .A(n989) );
  nor02 U1072 ( .Y(n990), .A0(B_not[32]), .A1(A[32]) );
  inv01 U1073 ( .Y(n979), .A(n990) );
  nor02 U1074 ( .Y(n991), .A0(n971), .A1(n972) );
  inv01 U1075 ( .Y(n981), .A(n991) );
  nor02 U1076 ( .Y(n992), .A0(n974), .A1(n976) );
  inv01 U1077 ( .Y(n982), .A(n992) );
  nor02 U1078 ( .Y(n993), .A0(n978), .A1(n980) );
  inv01 U1079 ( .Y(n983), .A(n993) );
  nor02 U1080 ( .Y(n994), .A0(n984), .A1(n985) );
  inv01 U1081 ( .Y(n987), .A(n994) );
  inv01 U1082 ( .Y(DIFF[12]), .A(n995) );
  inv02 U1083 ( .Y(carry_13_), .A(n996) );
  inv02 U1084 ( .Y(n997), .A(B_not[12]) );
  inv02 U1085 ( .Y(n998), .A(A[12]) );
  inv02 U1086 ( .Y(n999), .A(carry_12_) );
  nor02 U1087 ( .Y(n1000), .A0(n997), .A1(n1001) );
  nor02 U1088 ( .Y(n1002), .A0(n998), .A1(n1003) );
  nor02 U1089 ( .Y(n1004), .A0(n999), .A1(n1005) );
  nor02 U1090 ( .Y(n1006), .A0(n999), .A1(n1007) );
  nor02 U1091 ( .Y(n995), .A0(n1008), .A1(n1009) );
  nor02 U1092 ( .Y(n1010), .A0(n998), .A1(n999) );
  nor02 U1093 ( .Y(n1011), .A0(n997), .A1(n999) );
  nor02 U1094 ( .Y(n1012), .A0(n997), .A1(n998) );
  nor02 U1095 ( .Y(n996), .A0(n1012), .A1(n1013) );
  nor02 U1096 ( .Y(n1014), .A0(A[12]), .A1(carry_12_) );
  inv01 U1097 ( .Y(n1001), .A(n1014) );
  nor02 U1098 ( .Y(n1015), .A0(B_not[12]), .A1(carry_12_) );
  inv01 U1099 ( .Y(n1003), .A(n1015) );
  nor02 U1100 ( .Y(n1016), .A0(B_not[12]), .A1(A[12]) );
  inv01 U1101 ( .Y(n1005), .A(n1016) );
  nor02 U1102 ( .Y(n1017), .A0(n997), .A1(n998) );
  inv01 U1103 ( .Y(n1007), .A(n1017) );
  nor02 U1104 ( .Y(n1018), .A0(n1000), .A1(n1002) );
  inv01 U1105 ( .Y(n1008), .A(n1018) );
  nor02 U1106 ( .Y(n1019), .A0(n1004), .A1(n1006) );
  inv01 U1107 ( .Y(n1009), .A(n1019) );
  nor02 U1108 ( .Y(n1020), .A0(n1010), .A1(n1011) );
  inv01 U1109 ( .Y(n1013), .A(n1020) );
  inv01 U1110 ( .Y(DIFF[11]), .A(n1021) );
  inv02 U1111 ( .Y(carry_12_), .A(n1022) );
  inv02 U1112 ( .Y(n1023), .A(B_not[11]) );
  inv02 U1113 ( .Y(n1024), .A(A[11]) );
  inv02 U1114 ( .Y(n1025), .A(carry_11_) );
  nor02 U1115 ( .Y(n1026), .A0(n1023), .A1(n1027) );
  nor02 U1116 ( .Y(n1028), .A0(n1024), .A1(n1029) );
  nor02 U1117 ( .Y(n1030), .A0(n1025), .A1(n1031) );
  nor02 U1118 ( .Y(n1032), .A0(n1025), .A1(n1033) );
  nor02 U1119 ( .Y(n1021), .A0(n1034), .A1(n1035) );
  nor02 U1120 ( .Y(n1036), .A0(n1024), .A1(n1025) );
  nor02 U1121 ( .Y(n1037), .A0(n1023), .A1(n1025) );
  nor02 U1122 ( .Y(n1038), .A0(n1023), .A1(n1024) );
  nor02 U1123 ( .Y(n1022), .A0(n1038), .A1(n1039) );
  nor02 U1124 ( .Y(n1040), .A0(A[11]), .A1(carry_11_) );
  inv01 U1125 ( .Y(n1027), .A(n1040) );
  nor02 U1126 ( .Y(n1041), .A0(B_not[11]), .A1(carry_11_) );
  inv01 U1127 ( .Y(n1029), .A(n1041) );
  nor02 U1128 ( .Y(n1042), .A0(B_not[11]), .A1(A[11]) );
  inv01 U1129 ( .Y(n1031), .A(n1042) );
  nor02 U1130 ( .Y(n1043), .A0(n1023), .A1(n1024) );
  inv01 U1131 ( .Y(n1033), .A(n1043) );
  nor02 U1132 ( .Y(n1044), .A0(n1026), .A1(n1028) );
  inv01 U1133 ( .Y(n1034), .A(n1044) );
  nor02 U1134 ( .Y(n1045), .A0(n1030), .A1(n1032) );
  inv01 U1135 ( .Y(n1035), .A(n1045) );
  nor02 U1136 ( .Y(n1046), .A0(n1036), .A1(n1037) );
  inv01 U1137 ( .Y(n1039), .A(n1046) );
  inv01 U1138 ( .Y(DIFF[10]), .A(n1047) );
  inv02 U1139 ( .Y(carry_11_), .A(n1048) );
  inv02 U1140 ( .Y(n1049), .A(B_not[10]) );
  inv02 U1141 ( .Y(n1050), .A(A[10]) );
  inv02 U1142 ( .Y(n1051), .A(carry_10_) );
  nor02 U1143 ( .Y(n1052), .A0(n1049), .A1(n1053) );
  nor02 U1144 ( .Y(n1054), .A0(n1050), .A1(n1055) );
  nor02 U1145 ( .Y(n1056), .A0(n1051), .A1(n1057) );
  nor02 U1146 ( .Y(n1058), .A0(n1051), .A1(n1059) );
  nor02 U1147 ( .Y(n1047), .A0(n1060), .A1(n1061) );
  nor02 U1148 ( .Y(n1062), .A0(n1050), .A1(n1051) );
  nor02 U1149 ( .Y(n1063), .A0(n1049), .A1(n1051) );
  nor02 U1150 ( .Y(n1064), .A0(n1049), .A1(n1050) );
  nor02 U1151 ( .Y(n1048), .A0(n1064), .A1(n1065) );
  nor02 U1152 ( .Y(n1066), .A0(A[10]), .A1(carry_10_) );
  inv01 U1153 ( .Y(n1053), .A(n1066) );
  nor02 U1154 ( .Y(n1067), .A0(B_not[10]), .A1(carry_10_) );
  inv01 U1155 ( .Y(n1055), .A(n1067) );
  nor02 U1156 ( .Y(n1068), .A0(B_not[10]), .A1(A[10]) );
  inv01 U1157 ( .Y(n1057), .A(n1068) );
  nor02 U1158 ( .Y(n1069), .A0(n1049), .A1(n1050) );
  inv01 U1159 ( .Y(n1059), .A(n1069) );
  nor02 U1160 ( .Y(n1070), .A0(n1052), .A1(n1054) );
  inv01 U1161 ( .Y(n1060), .A(n1070) );
  nor02 U1162 ( .Y(n1071), .A0(n1056), .A1(n1058) );
  inv01 U1163 ( .Y(n1061), .A(n1071) );
  nor02 U1164 ( .Y(n1072), .A0(n1062), .A1(n1063) );
  inv01 U1165 ( .Y(n1065), .A(n1072) );
  inv02 U1166 ( .Y(B_not[10]), .A(n1314) );
  inv01 U1167 ( .Y(DIFF[9]), .A(n1073) );
  inv02 U1168 ( .Y(carry_10_), .A(n1074) );
  inv02 U1169 ( .Y(n1075), .A(B_not[9]) );
  inv02 U1170 ( .Y(n1076), .A(A[9]) );
  inv02 U1171 ( .Y(n1077), .A(carry_9_) );
  nor02 U1172 ( .Y(n1078), .A0(n1075), .A1(n1079) );
  nor02 U1173 ( .Y(n1080), .A0(n1076), .A1(n1081) );
  nor02 U1174 ( .Y(n1082), .A0(n1077), .A1(n1083) );
  nor02 U1175 ( .Y(n1084), .A0(n1077), .A1(n1085) );
  nor02 U1176 ( .Y(n1073), .A0(n1086), .A1(n1087) );
  nor02 U1177 ( .Y(n1088), .A0(n1076), .A1(n1077) );
  nor02 U1178 ( .Y(n1089), .A0(n1075), .A1(n1077) );
  nor02 U1179 ( .Y(n1090), .A0(n1075), .A1(n1076) );
  nor02 U1180 ( .Y(n1074), .A0(n1090), .A1(n1091) );
  nor02 U1181 ( .Y(n1092), .A0(A[9]), .A1(carry_9_) );
  inv01 U1182 ( .Y(n1079), .A(n1092) );
  nor02 U1183 ( .Y(n1093), .A0(B_not[9]), .A1(carry_9_) );
  inv01 U1184 ( .Y(n1081), .A(n1093) );
  nor02 U1185 ( .Y(n1094), .A0(B_not[9]), .A1(A[9]) );
  inv01 U1186 ( .Y(n1083), .A(n1094) );
  nor02 U1187 ( .Y(n1095), .A0(n1075), .A1(n1076) );
  inv01 U1188 ( .Y(n1085), .A(n1095) );
  nor02 U1189 ( .Y(n1096), .A0(n1078), .A1(n1080) );
  inv01 U1190 ( .Y(n1086), .A(n1096) );
  nor02 U1191 ( .Y(n1097), .A0(n1082), .A1(n1084) );
  inv01 U1192 ( .Y(n1087), .A(n1097) );
  nor02 U1193 ( .Y(n1098), .A0(n1088), .A1(n1089) );
  inv01 U1194 ( .Y(n1091), .A(n1098) );
  inv01 U1195 ( .Y(DIFF[8]), .A(n1099) );
  inv02 U1196 ( .Y(carry_9_), .A(n1100) );
  inv02 U1197 ( .Y(n1101), .A(B_not[8]) );
  inv02 U1198 ( .Y(n1102), .A(A[8]) );
  inv02 U1199 ( .Y(n1103), .A(carry_8_) );
  nor02 U1200 ( .Y(n1104), .A0(n1101), .A1(n1105) );
  nor02 U1201 ( .Y(n1106), .A0(n1102), .A1(n1107) );
  nor02 U1202 ( .Y(n1108), .A0(n1103), .A1(n1109) );
  nor02 U1203 ( .Y(n1110), .A0(n1103), .A1(n1111) );
  nor02 U1204 ( .Y(n1099), .A0(n1112), .A1(n1113) );
  nor02 U1205 ( .Y(n1114), .A0(n1102), .A1(n1103) );
  nor02 U1206 ( .Y(n1115), .A0(n1101), .A1(n1103) );
  nor02 U1207 ( .Y(n1116), .A0(n1101), .A1(n1102) );
  nor02 U1208 ( .Y(n1100), .A0(n1116), .A1(n1117) );
  nor02 U1209 ( .Y(n1118), .A0(A[8]), .A1(carry_8_) );
  inv01 U1210 ( .Y(n1105), .A(n1118) );
  nor02 U1211 ( .Y(n1119), .A0(B_not[8]), .A1(carry_8_) );
  inv01 U1212 ( .Y(n1107), .A(n1119) );
  nor02 U1213 ( .Y(n1120), .A0(B_not[8]), .A1(A[8]) );
  inv01 U1214 ( .Y(n1109), .A(n1120) );
  nor02 U1215 ( .Y(n1121), .A0(n1101), .A1(n1102) );
  inv01 U1216 ( .Y(n1111), .A(n1121) );
  nor02 U1217 ( .Y(n1122), .A0(n1104), .A1(n1106) );
  inv01 U1218 ( .Y(n1112), .A(n1122) );
  nor02 U1219 ( .Y(n1123), .A0(n1108), .A1(n1110) );
  inv01 U1220 ( .Y(n1113), .A(n1123) );
  nor02 U1221 ( .Y(n1124), .A0(n1114), .A1(n1115) );
  inv01 U1222 ( .Y(n1117), .A(n1124) );
  inv01 U1223 ( .Y(DIFF[7]), .A(n1125) );
  inv02 U1224 ( .Y(carry_8_), .A(n1126) );
  inv02 U1225 ( .Y(n1127), .A(B_not[7]) );
  inv02 U1226 ( .Y(n1128), .A(A[7]) );
  inv02 U1227 ( .Y(n1129), .A(carry_7_) );
  nor02 U1228 ( .Y(n1130), .A0(n1127), .A1(n1131) );
  nor02 U1229 ( .Y(n1132), .A0(n1128), .A1(n1133) );
  nor02 U1230 ( .Y(n1134), .A0(n1129), .A1(n1135) );
  nor02 U1231 ( .Y(n1136), .A0(n1129), .A1(n1137) );
  nor02 U1232 ( .Y(n1125), .A0(n1138), .A1(n1139) );
  nor02 U1233 ( .Y(n1140), .A0(n1128), .A1(n1129) );
  nor02 U1234 ( .Y(n1141), .A0(n1127), .A1(n1129) );
  nor02 U1235 ( .Y(n1142), .A0(n1127), .A1(n1128) );
  nor02 U1236 ( .Y(n1126), .A0(n1142), .A1(n1143) );
  nor02 U1237 ( .Y(n1144), .A0(A[7]), .A1(carry_7_) );
  inv01 U1238 ( .Y(n1131), .A(n1144) );
  nor02 U1239 ( .Y(n1145), .A0(B_not[7]), .A1(carry_7_) );
  inv01 U1240 ( .Y(n1133), .A(n1145) );
  nor02 U1241 ( .Y(n1146), .A0(B_not[7]), .A1(A[7]) );
  inv01 U1242 ( .Y(n1135), .A(n1146) );
  nor02 U1243 ( .Y(n1147), .A0(n1127), .A1(n1128) );
  inv01 U1244 ( .Y(n1137), .A(n1147) );
  nor02 U1245 ( .Y(n1148), .A0(n1130), .A1(n1132) );
  inv01 U1246 ( .Y(n1138), .A(n1148) );
  nor02 U1247 ( .Y(n1149), .A0(n1134), .A1(n1136) );
  inv01 U1248 ( .Y(n1139), .A(n1149) );
  nor02 U1249 ( .Y(n1150), .A0(n1140), .A1(n1141) );
  inv01 U1250 ( .Y(n1143), .A(n1150) );
  inv01 U1251 ( .Y(DIFF[6]), .A(n1151) );
  inv02 U1252 ( .Y(carry_7_), .A(n1152) );
  inv02 U1253 ( .Y(n1153), .A(B_not[6]) );
  inv02 U1254 ( .Y(n1154), .A(A[6]) );
  inv02 U1255 ( .Y(n1155), .A(carry_6_) );
  nor02 U1256 ( .Y(n1156), .A0(n1153), .A1(n1157) );
  nor02 U1257 ( .Y(n1158), .A0(n1154), .A1(n1159) );
  nor02 U1258 ( .Y(n1160), .A0(n1155), .A1(n1161) );
  nor02 U1259 ( .Y(n1162), .A0(n1155), .A1(n1163) );
  nor02 U1260 ( .Y(n1151), .A0(n1164), .A1(n1165) );
  nor02 U1261 ( .Y(n1166), .A0(n1154), .A1(n1155) );
  nor02 U1262 ( .Y(n1167), .A0(n1153), .A1(n1155) );
  nor02 U1263 ( .Y(n1168), .A0(n1153), .A1(n1154) );
  nor02 U1264 ( .Y(n1152), .A0(n1168), .A1(n1169) );
  nor02 U1265 ( .Y(n1170), .A0(A[6]), .A1(carry_6_) );
  inv01 U1266 ( .Y(n1157), .A(n1170) );
  nor02 U1267 ( .Y(n1171), .A0(B_not[6]), .A1(carry_6_) );
  inv01 U1268 ( .Y(n1159), .A(n1171) );
  nor02 U1269 ( .Y(n1172), .A0(B_not[6]), .A1(A[6]) );
  inv01 U1270 ( .Y(n1161), .A(n1172) );
  nor02 U1271 ( .Y(n1173), .A0(n1153), .A1(n1154) );
  inv01 U1272 ( .Y(n1163), .A(n1173) );
  nor02 U1273 ( .Y(n1174), .A0(n1156), .A1(n1158) );
  inv01 U1274 ( .Y(n1164), .A(n1174) );
  nor02 U1275 ( .Y(n1175), .A0(n1160), .A1(n1162) );
  inv01 U1276 ( .Y(n1165), .A(n1175) );
  nor02 U1277 ( .Y(n1176), .A0(n1166), .A1(n1167) );
  inv01 U1278 ( .Y(n1169), .A(n1176) );
  inv02 U1279 ( .Y(B_not[6]), .A(n1309) );
  inv01 U1280 ( .Y(DIFF[5]), .A(n1177) );
  inv02 U1281 ( .Y(carry_6_), .A(n1178) );
  inv02 U1282 ( .Y(n1179), .A(B_not[5]) );
  inv02 U1283 ( .Y(n1180), .A(A[5]) );
  inv02 U1284 ( .Y(n1181), .A(carry_5_) );
  nor02 U1285 ( .Y(n1182), .A0(n1179), .A1(n1183) );
  nor02 U1286 ( .Y(n1184), .A0(n1180), .A1(n1185) );
  nor02 U1287 ( .Y(n1186), .A0(n1181), .A1(n1187) );
  nor02 U1288 ( .Y(n1188), .A0(n1181), .A1(n1189) );
  nor02 U1289 ( .Y(n1177), .A0(n1190), .A1(n1191) );
  nor02 U1290 ( .Y(n1192), .A0(n1180), .A1(n1181) );
  nor02 U1291 ( .Y(n1193), .A0(n1179), .A1(n1181) );
  nor02 U1292 ( .Y(n1194), .A0(n1179), .A1(n1180) );
  nor02 U1293 ( .Y(n1178), .A0(n1194), .A1(n1195) );
  nor02 U1294 ( .Y(n1196), .A0(A[5]), .A1(carry_5_) );
  inv01 U1295 ( .Y(n1183), .A(n1196) );
  nor02 U1296 ( .Y(n1197), .A0(B_not[5]), .A1(carry_5_) );
  inv01 U1297 ( .Y(n1185), .A(n1197) );
  nor02 U1298 ( .Y(n1198), .A0(B_not[5]), .A1(A[5]) );
  inv01 U1299 ( .Y(n1187), .A(n1198) );
  nor02 U1300 ( .Y(n1199), .A0(n1179), .A1(n1180) );
  inv01 U1301 ( .Y(n1189), .A(n1199) );
  nor02 U1302 ( .Y(n1200), .A0(n1182), .A1(n1184) );
  inv01 U1303 ( .Y(n1190), .A(n1200) );
  nor02 U1304 ( .Y(n1201), .A0(n1186), .A1(n1188) );
  inv01 U1305 ( .Y(n1191), .A(n1201) );
  nor02 U1306 ( .Y(n1202), .A0(n1192), .A1(n1193) );
  inv01 U1307 ( .Y(n1195), .A(n1202) );
  inv02 U1308 ( .Y(B_not[5]), .A(n1310) );
  inv01 U1309 ( .Y(DIFF[4]), .A(n1203) );
  inv02 U1310 ( .Y(carry_5_), .A(n1204) );
  inv02 U1311 ( .Y(n1205), .A(B_not[4]) );
  inv02 U1312 ( .Y(n1206), .A(A[4]) );
  inv02 U1313 ( .Y(n1207), .A(carry_4_) );
  nor02 U1314 ( .Y(n1208), .A0(n1205), .A1(n1209) );
  nor02 U1315 ( .Y(n1210), .A0(n1206), .A1(n1211) );
  nor02 U1316 ( .Y(n1212), .A0(n1207), .A1(n1213) );
  nor02 U1317 ( .Y(n1214), .A0(n1207), .A1(n1215) );
  nor02 U1318 ( .Y(n1203), .A0(n1216), .A1(n1217) );
  nor02 U1319 ( .Y(n1218), .A0(n1206), .A1(n1207) );
  nor02 U1320 ( .Y(n1219), .A0(n1205), .A1(n1207) );
  nor02 U1321 ( .Y(n1220), .A0(n1205), .A1(n1206) );
  nor02 U1322 ( .Y(n1204), .A0(n1220), .A1(n1221) );
  nor02 U1323 ( .Y(n1222), .A0(A[4]), .A1(carry_4_) );
  inv01 U1324 ( .Y(n1209), .A(n1222) );
  nor02 U1325 ( .Y(n1223), .A0(B_not[4]), .A1(carry_4_) );
  inv01 U1326 ( .Y(n1211), .A(n1223) );
  nor02 U1327 ( .Y(n1224), .A0(B_not[4]), .A1(A[4]) );
  inv01 U1328 ( .Y(n1213), .A(n1224) );
  nor02 U1329 ( .Y(n1225), .A0(n1205), .A1(n1206) );
  inv01 U1330 ( .Y(n1215), .A(n1225) );
  nor02 U1331 ( .Y(n1226), .A0(n1208), .A1(n1210) );
  inv01 U1332 ( .Y(n1216), .A(n1226) );
  nor02 U1333 ( .Y(n1227), .A0(n1212), .A1(n1214) );
  inv01 U1334 ( .Y(n1217), .A(n1227) );
  nor02 U1335 ( .Y(n1228), .A0(n1218), .A1(n1219) );
  inv01 U1336 ( .Y(n1221), .A(n1228) );
  inv01 U1337 ( .Y(DIFF[3]), .A(n1229) );
  inv02 U1338 ( .Y(carry_4_), .A(n1230) );
  inv02 U1339 ( .Y(n1231), .A(B_not[3]) );
  inv02 U1340 ( .Y(n1232), .A(A[3]) );
  inv02 U1341 ( .Y(n1233), .A(carry_3_) );
  nor02 U1342 ( .Y(n1234), .A0(n1231), .A1(n1235) );
  nor02 U1343 ( .Y(n1236), .A0(n1232), .A1(n1237) );
  nor02 U1344 ( .Y(n1238), .A0(n1233), .A1(n1239) );
  nor02 U1345 ( .Y(n1240), .A0(n1233), .A1(n1241) );
  nor02 U1346 ( .Y(n1229), .A0(n1242), .A1(n1243) );
  nor02 U1347 ( .Y(n1244), .A0(n1232), .A1(n1233) );
  nor02 U1348 ( .Y(n1245), .A0(n1231), .A1(n1233) );
  nor02 U1349 ( .Y(n1246), .A0(n1231), .A1(n1232) );
  nor02 U1350 ( .Y(n1230), .A0(n1246), .A1(n1247) );
  nor02 U1351 ( .Y(n1248), .A0(A[3]), .A1(carry_3_) );
  inv01 U1352 ( .Y(n1235), .A(n1248) );
  nor02 U1353 ( .Y(n1249), .A0(B_not[3]), .A1(carry_3_) );
  inv01 U1354 ( .Y(n1237), .A(n1249) );
  nor02 U1355 ( .Y(n1250), .A0(B_not[3]), .A1(A[3]) );
  inv01 U1356 ( .Y(n1239), .A(n1250) );
  nor02 U1357 ( .Y(n1251), .A0(n1231), .A1(n1232) );
  inv01 U1358 ( .Y(n1241), .A(n1251) );
  nor02 U1359 ( .Y(n1252), .A0(n1234), .A1(n1236) );
  inv01 U1360 ( .Y(n1242), .A(n1252) );
  nor02 U1361 ( .Y(n1253), .A0(n1238), .A1(n1240) );
  inv01 U1362 ( .Y(n1243), .A(n1253) );
  nor02 U1363 ( .Y(n1254), .A0(n1244), .A1(n1245) );
  inv01 U1364 ( .Y(n1247), .A(n1254) );
  nor02 U1365 ( .Y(n1255), .A0(B_not[0]), .A1(A[0]) );
  inv02 U1366 ( .Y(n1256), .A(n1255) );
  inv01 U1367 ( .Y(DIFF[2]), .A(n1257) );
  inv02 U1368 ( .Y(carry_3_), .A(n1258) );
  inv02 U1369 ( .Y(n1259), .A(B_not[2]) );
  inv02 U1370 ( .Y(n1260), .A(A[2]) );
  inv02 U1371 ( .Y(n1261), .A(carry_2_) );
  nor02 U1372 ( .Y(n1262), .A0(n1259), .A1(n1263) );
  nor02 U1373 ( .Y(n1264), .A0(n1260), .A1(n1265) );
  nor02 U1374 ( .Y(n1266), .A0(n1261), .A1(n1267) );
  nor02 U1375 ( .Y(n1268), .A0(n1261), .A1(n1269) );
  nor02 U1376 ( .Y(n1257), .A0(n1270), .A1(n1271) );
  nor02 U1377 ( .Y(n1272), .A0(n1260), .A1(n1261) );
  nor02 U1378 ( .Y(n1273), .A0(n1259), .A1(n1261) );
  nor02 U1379 ( .Y(n1274), .A0(n1259), .A1(n1260) );
  nor02 U1380 ( .Y(n1258), .A0(n1274), .A1(n1275) );
  nor02 U1381 ( .Y(n1276), .A0(A[2]), .A1(carry_2_) );
  inv01 U1382 ( .Y(n1263), .A(n1276) );
  nor02 U1383 ( .Y(n1277), .A0(B_not[2]), .A1(carry_2_) );
  inv01 U1384 ( .Y(n1265), .A(n1277) );
  nor02 U1385 ( .Y(n1278), .A0(B_not[2]), .A1(A[2]) );
  inv01 U1386 ( .Y(n1267), .A(n1278) );
  nor02 U1387 ( .Y(n1279), .A0(n1259), .A1(n1260) );
  inv01 U1388 ( .Y(n1269), .A(n1279) );
  nor02 U1389 ( .Y(n1280), .A0(n1262), .A1(n1264) );
  inv01 U1390 ( .Y(n1270), .A(n1280) );
  nor02 U1391 ( .Y(n1281), .A0(n1266), .A1(n1268) );
  inv01 U1392 ( .Y(n1271), .A(n1281) );
  nor02 U1393 ( .Y(n1282), .A0(n1272), .A1(n1273) );
  inv01 U1394 ( .Y(n1275), .A(n1282) );
  inv01 U1395 ( .Y(DIFF[1]), .A(n1283) );
  inv02 U1396 ( .Y(carry_2_), .A(n1284) );
  inv02 U1397 ( .Y(n1285), .A(B_not[1]) );
  inv02 U1398 ( .Y(n1286), .A(A[1]) );
  inv02 U1399 ( .Y(n1287), .A(n1256) );
  nor02 U1400 ( .Y(n1288), .A0(n1285), .A1(n1289) );
  nor02 U1401 ( .Y(n1290), .A0(n1286), .A1(n1291) );
  nor02 U1402 ( .Y(n1292), .A0(n1287), .A1(n1293) );
  nor02 U1403 ( .Y(n1294), .A0(n1287), .A1(n1295) );
  nor02 U1404 ( .Y(n1283), .A0(n1296), .A1(n1297) );
  nor02 U1405 ( .Y(n1298), .A0(n1286), .A1(n1287) );
  nor02 U1406 ( .Y(n1299), .A0(n1285), .A1(n1287) );
  nor02 U1407 ( .Y(n1300), .A0(n1285), .A1(n1286) );
  nor02 U1408 ( .Y(n1284), .A0(n1300), .A1(n1301) );
  nor02 U1409 ( .Y(n1302), .A0(A[1]), .A1(n1256) );
  inv01 U1410 ( .Y(n1289), .A(n1302) );
  nor02 U1411 ( .Y(n1303), .A0(B_not[1]), .A1(n1256) );
  inv01 U1412 ( .Y(n1291), .A(n1303) );
  nor02 U1413 ( .Y(n1304), .A0(B_not[1]), .A1(A[1]) );
  inv01 U1414 ( .Y(n1293), .A(n1304) );
  nor02 U1415 ( .Y(n1305), .A0(n1285), .A1(n1286) );
  inv01 U1416 ( .Y(n1295), .A(n1305) );
  nor02 U1417 ( .Y(n1306), .A0(n1288), .A1(n1290) );
  inv01 U1418 ( .Y(n1296), .A(n1306) );
  nor02 U1419 ( .Y(n1307), .A0(n1292), .A1(n1294) );
  inv01 U1420 ( .Y(n1297), .A(n1307) );
  nor02 U1421 ( .Y(n1308), .A0(n1298), .A1(n1299) );
  inv01 U1422 ( .Y(n1301), .A(n1308) );
  buf02 U1423 ( .Y(n1309), .A(B[6]) );
  inv02 U1424 ( .Y(B_not[7]), .A(B[7]) );
  buf02 U1425 ( .Y(n1310), .A(B[5]) );
  inv02 U1426 ( .Y(B_not[18]), .A(B[18]) );
  inv02 U1427 ( .Y(B_not[16]), .A(B[16]) );
  inv02 U1428 ( .Y(B_not[19]), .A(B[19]) );
  inv02 U1429 ( .Y(B_not[17]), .A(B[17]) );
  inv02 U1430 ( .Y(B_not[40]), .A(B[40]) );
  inv02 U1431 ( .Y(B_not[51]), .A(B[51]) );
  inv02 U1432 ( .Y(B_not[44]), .A(B[44]) );
  inv02 U1433 ( .Y(B_not[45]), .A(B[45]) );
  inv02 U1434 ( .Y(B_not[47]), .A(B[47]) );
  inv02 U1435 ( .Y(B_not[36]), .A(B[36]) );
  inv02 U1436 ( .Y(B_not[48]), .A(B[48]) );
  inv02 U1437 ( .Y(B_not[41]), .A(B[41]) );
  inv02 U1438 ( .Y(B_not[39]), .A(B[39]) );
  inv02 U1439 ( .Y(B_not[37]), .A(B[37]) );
  inv02 U1440 ( .Y(B_not[38]), .A(B[38]) );
  inv02 U1441 ( .Y(B_not[22]), .A(B[22]) );
  buf02 U1442 ( .Y(n1311), .A(B[34]) );
  inv02 U1443 ( .Y(B_not[29]), .A(B[29]) );
  inv02 U1444 ( .Y(B_not[26]), .A(B[26]) );
  inv02 U1445 ( .Y(B_not[27]), .A(B[27]) );
  buf02 U1446 ( .Y(n1312), .A(B[30]) );
  inv02 U1447 ( .Y(B_not[35]), .A(B[35]) );
  inv02 U1448 ( .Y(B_not[20]), .A(B[20]) );
  inv02 U1449 ( .Y(B_not[32]), .A(B[32]) );
  buf02 U1450 ( .Y(n1313), .A(B[24]) );
  inv02 U1451 ( .Y(B_not[25]), .A(B[25]) );
  inv02 U1452 ( .Y(B_not[28]), .A(B[28]) );
  inv02 U1453 ( .Y(B_not[33]), .A(B[33]) );
  inv02 U1454 ( .Y(B_not[31]), .A(B[31]) );
  inv02 U1455 ( .Y(B_not[2]), .A(B[2]) );
  inv02 U1456 ( .Y(B_not[1]), .A(B[1]) );
  inv02 U1457 ( .Y(B_not[3]), .A(B[3]) );
  inv02 U1458 ( .Y(B_not[0]), .A(B[0]) );
  inv02 U1459 ( .Y(B_not[13]), .A(B[13]) );
  inv02 U1460 ( .Y(B_not[15]), .A(B[15]) );
  inv02 U1461 ( .Y(B_not[14]), .A(B[14]) );
  buf02 U1462 ( .Y(n1314), .A(B[10]) );
  inv02 U1463 ( .Y(B_not[8]), .A(B[8]) );
  inv02 U1464 ( .Y(B_not[9]), .A(B[9]) );
  inv02 U1465 ( .Y(B_not[12]), .A(B[12]) );
  inv02 U1466 ( .Y(B_not[11]), .A(B[11]) );
  inv02 U1467 ( .Y(B_not[4]), .A(B[4]) );
  fadd1 U2_51 ( .S(DIFF[51]), .A(A[51]), .B(B_not[51]), .CI(carry_51_) );
endmodule


module sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_add_26_0 ( A, B, CI, SUM, CO );
  input [25:0] A;
  input [25:0] B;
  output [25:0] SUM;
  input CI;
  output CO;
  wire   carry_25_, carry_24_, carry_23_, carry_22_, carry_21_, carry_20_,
         carry_19_, carry_18_, carry_17_, carry_16_, carry_15_, carry_14_,
         carry_13_, carry_12_, carry_11_, carry_10_, carry_9_, carry_8_,
         carry_7_, carry_6_, carry_5_, carry_4_, carry_3_, carry_2_, carry_1_,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625;

  and02 U4 ( .Y(n1), .A0(A[0]), .A1(B[0]) );
  inv01 U5 ( .Y(SUM[24]), .A(n2) );
  inv02 U6 ( .Y(carry_25_), .A(n3) );
  inv02 U7 ( .Y(n4), .A(B[24]) );
  inv02 U8 ( .Y(n5), .A(A[24]) );
  inv02 U9 ( .Y(n6), .A(carry_24_) );
  nor02 U10 ( .Y(n7), .A0(n4), .A1(n8) );
  nor02 U11 ( .Y(n9), .A0(n5), .A1(n10) );
  nor02 U12 ( .Y(n11), .A0(n6), .A1(n12) );
  nor02 U13 ( .Y(n13), .A0(n6), .A1(n14) );
  nor02 U14 ( .Y(n2), .A0(n15), .A1(n16) );
  nor02 U15 ( .Y(n17), .A0(n5), .A1(n6) );
  nor02 U16 ( .Y(n18), .A0(n4), .A1(n6) );
  nor02 U17 ( .Y(n19), .A0(n4), .A1(n5) );
  nor02 U18 ( .Y(n3), .A0(n19), .A1(n20) );
  nor02 U19 ( .Y(n21), .A0(A[24]), .A1(carry_24_) );
  inv01 U20 ( .Y(n8), .A(n21) );
  nor02 U21 ( .Y(n22), .A0(B[24]), .A1(carry_24_) );
  inv01 U22 ( .Y(n10), .A(n22) );
  nor02 U23 ( .Y(n23), .A0(B[24]), .A1(A[24]) );
  inv01 U24 ( .Y(n12), .A(n23) );
  nor02 U25 ( .Y(n24), .A0(n4), .A1(n5) );
  inv01 U26 ( .Y(n14), .A(n24) );
  nor02 U27 ( .Y(n25), .A0(n7), .A1(n9) );
  inv01 U28 ( .Y(n15), .A(n25) );
  nor02 U29 ( .Y(n26), .A0(n11), .A1(n13) );
  inv01 U30 ( .Y(n16), .A(n26) );
  nor02 U31 ( .Y(n27), .A0(n17), .A1(n18) );
  inv01 U32 ( .Y(n20), .A(n27) );
  inv01 U33 ( .Y(SUM[23]), .A(n28) );
  inv02 U34 ( .Y(carry_24_), .A(n29) );
  inv02 U35 ( .Y(n30), .A(B[23]) );
  inv02 U36 ( .Y(n31), .A(A[23]) );
  inv02 U37 ( .Y(n32), .A(carry_23_) );
  nor02 U38 ( .Y(n33), .A0(n30), .A1(n34) );
  nor02 U39 ( .Y(n35), .A0(n31), .A1(n36) );
  nor02 U40 ( .Y(n37), .A0(n32), .A1(n38) );
  nor02 U41 ( .Y(n39), .A0(n32), .A1(n40) );
  nor02 U42 ( .Y(n28), .A0(n41), .A1(n42) );
  nor02 U43 ( .Y(n43), .A0(n31), .A1(n32) );
  nor02 U44 ( .Y(n44), .A0(n30), .A1(n32) );
  nor02 U45 ( .Y(n45), .A0(n30), .A1(n31) );
  nor02 U46 ( .Y(n29), .A0(n45), .A1(n46) );
  nor02 U47 ( .Y(n47), .A0(A[23]), .A1(carry_23_) );
  inv01 U48 ( .Y(n34), .A(n47) );
  nor02 U49 ( .Y(n48), .A0(B[23]), .A1(carry_23_) );
  inv01 U50 ( .Y(n36), .A(n48) );
  nor02 U51 ( .Y(n49), .A0(B[23]), .A1(A[23]) );
  inv01 U52 ( .Y(n38), .A(n49) );
  nor02 U53 ( .Y(n50), .A0(n30), .A1(n31) );
  inv01 U54 ( .Y(n40), .A(n50) );
  nor02 U55 ( .Y(n51), .A0(n33), .A1(n35) );
  inv01 U56 ( .Y(n41), .A(n51) );
  nor02 U57 ( .Y(n52), .A0(n37), .A1(n39) );
  inv01 U58 ( .Y(n42), .A(n52) );
  nor02 U59 ( .Y(n53), .A0(n43), .A1(n44) );
  inv01 U60 ( .Y(n46), .A(n53) );
  inv01 U61 ( .Y(SUM[22]), .A(n54) );
  inv02 U62 ( .Y(carry_23_), .A(n55) );
  inv02 U63 ( .Y(n56), .A(B[22]) );
  inv02 U64 ( .Y(n57), .A(A[22]) );
  inv02 U65 ( .Y(n58), .A(carry_22_) );
  nor02 U66 ( .Y(n59), .A0(n56), .A1(n60) );
  nor02 U67 ( .Y(n61), .A0(n57), .A1(n62) );
  nor02 U68 ( .Y(n63), .A0(n58), .A1(n64) );
  nor02 U69 ( .Y(n65), .A0(n58), .A1(n66) );
  nor02 U70 ( .Y(n54), .A0(n67), .A1(n68) );
  nor02 U71 ( .Y(n69), .A0(n57), .A1(n58) );
  nor02 U72 ( .Y(n70), .A0(n56), .A1(n58) );
  nor02 U73 ( .Y(n71), .A0(n56), .A1(n57) );
  nor02 U74 ( .Y(n55), .A0(n71), .A1(n72) );
  nor02 U75 ( .Y(n73), .A0(A[22]), .A1(carry_22_) );
  inv01 U76 ( .Y(n60), .A(n73) );
  nor02 U77 ( .Y(n74), .A0(B[22]), .A1(carry_22_) );
  inv01 U78 ( .Y(n62), .A(n74) );
  nor02 U79 ( .Y(n75), .A0(B[22]), .A1(A[22]) );
  inv01 U80 ( .Y(n64), .A(n75) );
  nor02 U81 ( .Y(n76), .A0(n56), .A1(n57) );
  inv01 U82 ( .Y(n66), .A(n76) );
  nor02 U83 ( .Y(n77), .A0(n59), .A1(n61) );
  inv01 U84 ( .Y(n67), .A(n77) );
  nor02 U85 ( .Y(n78), .A0(n63), .A1(n65) );
  inv01 U86 ( .Y(n68), .A(n78) );
  nor02 U87 ( .Y(n79), .A0(n69), .A1(n70) );
  inv01 U88 ( .Y(n72), .A(n79) );
  inv01 U89 ( .Y(SUM[21]), .A(n80) );
  inv02 U90 ( .Y(carry_22_), .A(n81) );
  inv02 U91 ( .Y(n82), .A(B[21]) );
  inv02 U92 ( .Y(n83), .A(A[21]) );
  inv02 U93 ( .Y(n84), .A(carry_21_) );
  nor02 U94 ( .Y(n85), .A0(n82), .A1(n86) );
  nor02 U95 ( .Y(n87), .A0(n83), .A1(n88) );
  nor02 U96 ( .Y(n89), .A0(n84), .A1(n90) );
  nor02 U97 ( .Y(n91), .A0(n84), .A1(n92) );
  nor02 U98 ( .Y(n80), .A0(n93), .A1(n94) );
  nor02 U99 ( .Y(n95), .A0(n83), .A1(n84) );
  nor02 U100 ( .Y(n96), .A0(n82), .A1(n84) );
  nor02 U101 ( .Y(n97), .A0(n82), .A1(n83) );
  nor02 U102 ( .Y(n81), .A0(n97), .A1(n98) );
  nor02 U103 ( .Y(n99), .A0(A[21]), .A1(carry_21_) );
  inv01 U104 ( .Y(n86), .A(n99) );
  nor02 U105 ( .Y(n100), .A0(B[21]), .A1(carry_21_) );
  inv01 U106 ( .Y(n88), .A(n100) );
  nor02 U107 ( .Y(n101), .A0(B[21]), .A1(A[21]) );
  inv01 U108 ( .Y(n90), .A(n101) );
  nor02 U109 ( .Y(n102), .A0(n82), .A1(n83) );
  inv01 U110 ( .Y(n92), .A(n102) );
  nor02 U111 ( .Y(n103), .A0(n85), .A1(n87) );
  inv01 U112 ( .Y(n93), .A(n103) );
  nor02 U113 ( .Y(n104), .A0(n89), .A1(n91) );
  inv01 U114 ( .Y(n94), .A(n104) );
  nor02 U115 ( .Y(n105), .A0(n95), .A1(n96) );
  inv01 U116 ( .Y(n98), .A(n105) );
  inv01 U117 ( .Y(SUM[20]), .A(n106) );
  inv02 U118 ( .Y(carry_21_), .A(n107) );
  inv02 U119 ( .Y(n108), .A(B[20]) );
  inv02 U120 ( .Y(n109), .A(A[20]) );
  inv02 U121 ( .Y(n110), .A(carry_20_) );
  nor02 U122 ( .Y(n111), .A0(n108), .A1(n112) );
  nor02 U123 ( .Y(n113), .A0(n109), .A1(n114) );
  nor02 U124 ( .Y(n115), .A0(n110), .A1(n116) );
  nor02 U125 ( .Y(n117), .A0(n110), .A1(n118) );
  nor02 U126 ( .Y(n106), .A0(n119), .A1(n120) );
  nor02 U127 ( .Y(n121), .A0(n109), .A1(n110) );
  nor02 U128 ( .Y(n122), .A0(n108), .A1(n110) );
  nor02 U129 ( .Y(n123), .A0(n108), .A1(n109) );
  nor02 U130 ( .Y(n107), .A0(n123), .A1(n124) );
  nor02 U131 ( .Y(n125), .A0(A[20]), .A1(carry_20_) );
  inv01 U132 ( .Y(n112), .A(n125) );
  nor02 U133 ( .Y(n126), .A0(B[20]), .A1(carry_20_) );
  inv01 U134 ( .Y(n114), .A(n126) );
  nor02 U135 ( .Y(n127), .A0(B[20]), .A1(A[20]) );
  inv01 U136 ( .Y(n116), .A(n127) );
  nor02 U137 ( .Y(n128), .A0(n108), .A1(n109) );
  inv01 U138 ( .Y(n118), .A(n128) );
  nor02 U139 ( .Y(n129), .A0(n111), .A1(n113) );
  inv01 U140 ( .Y(n119), .A(n129) );
  nor02 U141 ( .Y(n130), .A0(n115), .A1(n117) );
  inv01 U142 ( .Y(n120), .A(n130) );
  nor02 U143 ( .Y(n131), .A0(n121), .A1(n122) );
  inv01 U144 ( .Y(n124), .A(n131) );
  inv01 U145 ( .Y(SUM[19]), .A(n132) );
  inv02 U146 ( .Y(carry_20_), .A(n133) );
  inv02 U147 ( .Y(n134), .A(B[19]) );
  inv02 U148 ( .Y(n135), .A(A[19]) );
  inv02 U149 ( .Y(n136), .A(carry_19_) );
  nor02 U150 ( .Y(n137), .A0(n134), .A1(n138) );
  nor02 U151 ( .Y(n139), .A0(n135), .A1(n140) );
  nor02 U152 ( .Y(n141), .A0(n136), .A1(n142) );
  nor02 U153 ( .Y(n143), .A0(n136), .A1(n144) );
  nor02 U154 ( .Y(n132), .A0(n145), .A1(n146) );
  nor02 U155 ( .Y(n147), .A0(n135), .A1(n136) );
  nor02 U156 ( .Y(n148), .A0(n134), .A1(n136) );
  nor02 U157 ( .Y(n149), .A0(n134), .A1(n135) );
  nor02 U158 ( .Y(n133), .A0(n149), .A1(n150) );
  nor02 U159 ( .Y(n151), .A0(A[19]), .A1(carry_19_) );
  inv01 U160 ( .Y(n138), .A(n151) );
  nor02 U161 ( .Y(n152), .A0(B[19]), .A1(carry_19_) );
  inv01 U162 ( .Y(n140), .A(n152) );
  nor02 U163 ( .Y(n153), .A0(B[19]), .A1(A[19]) );
  inv01 U164 ( .Y(n142), .A(n153) );
  nor02 U165 ( .Y(n154), .A0(n134), .A1(n135) );
  inv01 U166 ( .Y(n144), .A(n154) );
  nor02 U167 ( .Y(n155), .A0(n137), .A1(n139) );
  inv01 U168 ( .Y(n145), .A(n155) );
  nor02 U169 ( .Y(n156), .A0(n141), .A1(n143) );
  inv01 U170 ( .Y(n146), .A(n156) );
  nor02 U171 ( .Y(n157), .A0(n147), .A1(n148) );
  inv01 U172 ( .Y(n150), .A(n157) );
  inv01 U173 ( .Y(SUM[18]), .A(n158) );
  inv02 U174 ( .Y(carry_19_), .A(n159) );
  inv02 U175 ( .Y(n160), .A(B[18]) );
  inv02 U176 ( .Y(n161), .A(A[18]) );
  inv02 U177 ( .Y(n162), .A(carry_18_) );
  nor02 U178 ( .Y(n163), .A0(n160), .A1(n164) );
  nor02 U179 ( .Y(n165), .A0(n161), .A1(n166) );
  nor02 U180 ( .Y(n167), .A0(n162), .A1(n168) );
  nor02 U181 ( .Y(n169), .A0(n162), .A1(n170) );
  nor02 U182 ( .Y(n158), .A0(n171), .A1(n172) );
  nor02 U183 ( .Y(n173), .A0(n161), .A1(n162) );
  nor02 U184 ( .Y(n174), .A0(n160), .A1(n162) );
  nor02 U185 ( .Y(n175), .A0(n160), .A1(n161) );
  nor02 U186 ( .Y(n159), .A0(n175), .A1(n176) );
  nor02 U187 ( .Y(n177), .A0(A[18]), .A1(carry_18_) );
  inv01 U188 ( .Y(n164), .A(n177) );
  nor02 U189 ( .Y(n178), .A0(B[18]), .A1(carry_18_) );
  inv01 U190 ( .Y(n166), .A(n178) );
  nor02 U191 ( .Y(n179), .A0(B[18]), .A1(A[18]) );
  inv01 U192 ( .Y(n168), .A(n179) );
  nor02 U193 ( .Y(n180), .A0(n160), .A1(n161) );
  inv01 U194 ( .Y(n170), .A(n180) );
  nor02 U195 ( .Y(n181), .A0(n163), .A1(n165) );
  inv01 U196 ( .Y(n171), .A(n181) );
  nor02 U197 ( .Y(n182), .A0(n167), .A1(n169) );
  inv01 U198 ( .Y(n172), .A(n182) );
  nor02 U199 ( .Y(n183), .A0(n173), .A1(n174) );
  inv01 U200 ( .Y(n176), .A(n183) );
  inv01 U201 ( .Y(SUM[17]), .A(n184) );
  inv02 U202 ( .Y(carry_18_), .A(n185) );
  inv02 U203 ( .Y(n186), .A(B[17]) );
  inv02 U204 ( .Y(n187), .A(A[17]) );
  inv02 U205 ( .Y(n188), .A(carry_17_) );
  nor02 U206 ( .Y(n189), .A0(n186), .A1(n190) );
  nor02 U207 ( .Y(n191), .A0(n187), .A1(n192) );
  nor02 U208 ( .Y(n193), .A0(n188), .A1(n194) );
  nor02 U209 ( .Y(n195), .A0(n188), .A1(n196) );
  nor02 U210 ( .Y(n184), .A0(n197), .A1(n198) );
  nor02 U211 ( .Y(n199), .A0(n187), .A1(n188) );
  nor02 U212 ( .Y(n200), .A0(n186), .A1(n188) );
  nor02 U213 ( .Y(n201), .A0(n186), .A1(n187) );
  nor02 U214 ( .Y(n185), .A0(n201), .A1(n202) );
  nor02 U215 ( .Y(n203), .A0(A[17]), .A1(carry_17_) );
  inv01 U216 ( .Y(n190), .A(n203) );
  nor02 U217 ( .Y(n204), .A0(B[17]), .A1(carry_17_) );
  inv01 U218 ( .Y(n192), .A(n204) );
  nor02 U219 ( .Y(n205), .A0(B[17]), .A1(A[17]) );
  inv01 U220 ( .Y(n194), .A(n205) );
  nor02 U221 ( .Y(n206), .A0(n186), .A1(n187) );
  inv01 U222 ( .Y(n196), .A(n206) );
  nor02 U223 ( .Y(n207), .A0(n189), .A1(n191) );
  inv01 U224 ( .Y(n197), .A(n207) );
  nor02 U225 ( .Y(n208), .A0(n193), .A1(n195) );
  inv01 U226 ( .Y(n198), .A(n208) );
  nor02 U227 ( .Y(n209), .A0(n199), .A1(n200) );
  inv01 U228 ( .Y(n202), .A(n209) );
  inv01 U229 ( .Y(SUM[16]), .A(n210) );
  inv02 U230 ( .Y(carry_17_), .A(n211) );
  inv02 U231 ( .Y(n212), .A(B[16]) );
  inv02 U232 ( .Y(n213), .A(A[16]) );
  inv02 U233 ( .Y(n214), .A(carry_16_) );
  nor02 U234 ( .Y(n215), .A0(n212), .A1(n216) );
  nor02 U235 ( .Y(n217), .A0(n213), .A1(n218) );
  nor02 U236 ( .Y(n219), .A0(n214), .A1(n220) );
  nor02 U237 ( .Y(n221), .A0(n214), .A1(n222) );
  nor02 U238 ( .Y(n210), .A0(n223), .A1(n224) );
  nor02 U239 ( .Y(n225), .A0(n213), .A1(n214) );
  nor02 U240 ( .Y(n226), .A0(n212), .A1(n214) );
  nor02 U241 ( .Y(n227), .A0(n212), .A1(n213) );
  nor02 U242 ( .Y(n211), .A0(n227), .A1(n228) );
  nor02 U243 ( .Y(n229), .A0(A[16]), .A1(carry_16_) );
  inv01 U244 ( .Y(n216), .A(n229) );
  nor02 U245 ( .Y(n230), .A0(B[16]), .A1(carry_16_) );
  inv01 U246 ( .Y(n218), .A(n230) );
  nor02 U247 ( .Y(n231), .A0(B[16]), .A1(A[16]) );
  inv01 U248 ( .Y(n220), .A(n231) );
  nor02 U249 ( .Y(n232), .A0(n212), .A1(n213) );
  inv01 U250 ( .Y(n222), .A(n232) );
  nor02 U251 ( .Y(n233), .A0(n215), .A1(n217) );
  inv01 U252 ( .Y(n223), .A(n233) );
  nor02 U253 ( .Y(n234), .A0(n219), .A1(n221) );
  inv01 U254 ( .Y(n224), .A(n234) );
  nor02 U255 ( .Y(n235), .A0(n225), .A1(n226) );
  inv01 U256 ( .Y(n228), .A(n235) );
  inv01 U257 ( .Y(SUM[15]), .A(n236) );
  inv02 U258 ( .Y(carry_16_), .A(n237) );
  inv02 U259 ( .Y(n238), .A(B[15]) );
  inv02 U260 ( .Y(n239), .A(A[15]) );
  inv02 U261 ( .Y(n240), .A(carry_15_) );
  nor02 U262 ( .Y(n241), .A0(n238), .A1(n242) );
  nor02 U263 ( .Y(n243), .A0(n239), .A1(n244) );
  nor02 U264 ( .Y(n245), .A0(n240), .A1(n246) );
  nor02 U265 ( .Y(n247), .A0(n240), .A1(n248) );
  nor02 U266 ( .Y(n236), .A0(n249), .A1(n250) );
  nor02 U267 ( .Y(n251), .A0(n239), .A1(n240) );
  nor02 U268 ( .Y(n252), .A0(n238), .A1(n240) );
  nor02 U269 ( .Y(n253), .A0(n238), .A1(n239) );
  nor02 U270 ( .Y(n237), .A0(n253), .A1(n254) );
  nor02 U271 ( .Y(n255), .A0(A[15]), .A1(carry_15_) );
  inv01 U272 ( .Y(n242), .A(n255) );
  nor02 U273 ( .Y(n256), .A0(B[15]), .A1(carry_15_) );
  inv01 U274 ( .Y(n244), .A(n256) );
  nor02 U275 ( .Y(n257), .A0(B[15]), .A1(A[15]) );
  inv01 U276 ( .Y(n246), .A(n257) );
  nor02 U277 ( .Y(n258), .A0(n238), .A1(n239) );
  inv01 U278 ( .Y(n248), .A(n258) );
  nor02 U279 ( .Y(n259), .A0(n241), .A1(n243) );
  inv01 U280 ( .Y(n249), .A(n259) );
  nor02 U281 ( .Y(n260), .A0(n245), .A1(n247) );
  inv01 U282 ( .Y(n250), .A(n260) );
  nor02 U283 ( .Y(n261), .A0(n251), .A1(n252) );
  inv01 U284 ( .Y(n254), .A(n261) );
  inv01 U285 ( .Y(SUM[14]), .A(n262) );
  inv02 U286 ( .Y(carry_15_), .A(n263) );
  inv02 U287 ( .Y(n264), .A(B[14]) );
  inv02 U288 ( .Y(n265), .A(A[14]) );
  inv02 U289 ( .Y(n266), .A(carry_14_) );
  nor02 U290 ( .Y(n267), .A0(n264), .A1(n268) );
  nor02 U291 ( .Y(n269), .A0(n265), .A1(n270) );
  nor02 U292 ( .Y(n271), .A0(n266), .A1(n272) );
  nor02 U293 ( .Y(n273), .A0(n266), .A1(n274) );
  nor02 U294 ( .Y(n262), .A0(n275), .A1(n276) );
  nor02 U295 ( .Y(n277), .A0(n265), .A1(n266) );
  nor02 U296 ( .Y(n278), .A0(n264), .A1(n266) );
  nor02 U297 ( .Y(n279), .A0(n264), .A1(n265) );
  nor02 U298 ( .Y(n263), .A0(n279), .A1(n280) );
  nor02 U299 ( .Y(n281), .A0(A[14]), .A1(carry_14_) );
  inv01 U300 ( .Y(n268), .A(n281) );
  nor02 U301 ( .Y(n282), .A0(B[14]), .A1(carry_14_) );
  inv01 U302 ( .Y(n270), .A(n282) );
  nor02 U303 ( .Y(n283), .A0(B[14]), .A1(A[14]) );
  inv01 U304 ( .Y(n272), .A(n283) );
  nor02 U305 ( .Y(n284), .A0(n264), .A1(n265) );
  inv01 U306 ( .Y(n274), .A(n284) );
  nor02 U307 ( .Y(n285), .A0(n267), .A1(n269) );
  inv01 U308 ( .Y(n275), .A(n285) );
  nor02 U309 ( .Y(n286), .A0(n271), .A1(n273) );
  inv01 U310 ( .Y(n276), .A(n286) );
  nor02 U311 ( .Y(n287), .A0(n277), .A1(n278) );
  inv01 U312 ( .Y(n280), .A(n287) );
  inv01 U313 ( .Y(SUM[13]), .A(n288) );
  inv02 U314 ( .Y(carry_14_), .A(n289) );
  inv02 U315 ( .Y(n290), .A(B[13]) );
  inv02 U316 ( .Y(n291), .A(A[13]) );
  inv02 U317 ( .Y(n292), .A(carry_13_) );
  nor02 U318 ( .Y(n293), .A0(n290), .A1(n294) );
  nor02 U319 ( .Y(n295), .A0(n291), .A1(n296) );
  nor02 U320 ( .Y(n297), .A0(n292), .A1(n298) );
  nor02 U321 ( .Y(n299), .A0(n292), .A1(n300) );
  nor02 U322 ( .Y(n288), .A0(n301), .A1(n302) );
  nor02 U323 ( .Y(n303), .A0(n291), .A1(n292) );
  nor02 U324 ( .Y(n304), .A0(n290), .A1(n292) );
  nor02 U325 ( .Y(n305), .A0(n290), .A1(n291) );
  nor02 U326 ( .Y(n289), .A0(n305), .A1(n306) );
  nor02 U327 ( .Y(n307), .A0(A[13]), .A1(carry_13_) );
  inv01 U328 ( .Y(n294), .A(n307) );
  nor02 U329 ( .Y(n308), .A0(B[13]), .A1(carry_13_) );
  inv01 U330 ( .Y(n296), .A(n308) );
  nor02 U331 ( .Y(n309), .A0(B[13]), .A1(A[13]) );
  inv01 U332 ( .Y(n298), .A(n309) );
  nor02 U333 ( .Y(n310), .A0(n290), .A1(n291) );
  inv01 U334 ( .Y(n300), .A(n310) );
  nor02 U335 ( .Y(n311), .A0(n293), .A1(n295) );
  inv01 U336 ( .Y(n301), .A(n311) );
  nor02 U337 ( .Y(n312), .A0(n297), .A1(n299) );
  inv01 U338 ( .Y(n302), .A(n312) );
  nor02 U339 ( .Y(n313), .A0(n303), .A1(n304) );
  inv01 U340 ( .Y(n306), .A(n313) );
  inv01 U341 ( .Y(SUM[12]), .A(n314) );
  inv02 U342 ( .Y(carry_13_), .A(n315) );
  inv02 U343 ( .Y(n316), .A(B[12]) );
  inv02 U344 ( .Y(n317), .A(A[12]) );
  inv02 U345 ( .Y(n318), .A(carry_12_) );
  nor02 U346 ( .Y(n319), .A0(n316), .A1(n320) );
  nor02 U347 ( .Y(n321), .A0(n317), .A1(n322) );
  nor02 U348 ( .Y(n323), .A0(n318), .A1(n324) );
  nor02 U349 ( .Y(n325), .A0(n318), .A1(n326) );
  nor02 U350 ( .Y(n314), .A0(n327), .A1(n328) );
  nor02 U351 ( .Y(n329), .A0(n317), .A1(n318) );
  nor02 U352 ( .Y(n330), .A0(n316), .A1(n318) );
  nor02 U353 ( .Y(n331), .A0(n316), .A1(n317) );
  nor02 U354 ( .Y(n315), .A0(n331), .A1(n332) );
  nor02 U355 ( .Y(n333), .A0(A[12]), .A1(carry_12_) );
  inv01 U356 ( .Y(n320), .A(n333) );
  nor02 U357 ( .Y(n334), .A0(B[12]), .A1(carry_12_) );
  inv01 U358 ( .Y(n322), .A(n334) );
  nor02 U359 ( .Y(n335), .A0(B[12]), .A1(A[12]) );
  inv01 U360 ( .Y(n324), .A(n335) );
  nor02 U361 ( .Y(n336), .A0(n316), .A1(n317) );
  inv01 U362 ( .Y(n326), .A(n336) );
  nor02 U363 ( .Y(n337), .A0(n319), .A1(n321) );
  inv01 U364 ( .Y(n327), .A(n337) );
  nor02 U365 ( .Y(n338), .A0(n323), .A1(n325) );
  inv01 U366 ( .Y(n328), .A(n338) );
  nor02 U367 ( .Y(n339), .A0(n329), .A1(n330) );
  inv01 U368 ( .Y(n332), .A(n339) );
  inv01 U369 ( .Y(SUM[11]), .A(n340) );
  inv02 U370 ( .Y(carry_12_), .A(n341) );
  inv02 U371 ( .Y(n342), .A(B[11]) );
  inv02 U372 ( .Y(n343), .A(A[11]) );
  inv02 U373 ( .Y(n344), .A(carry_11_) );
  nor02 U374 ( .Y(n345), .A0(n342), .A1(n346) );
  nor02 U375 ( .Y(n347), .A0(n343), .A1(n348) );
  nor02 U376 ( .Y(n349), .A0(n344), .A1(n350) );
  nor02 U377 ( .Y(n351), .A0(n344), .A1(n352) );
  nor02 U378 ( .Y(n340), .A0(n353), .A1(n354) );
  nor02 U379 ( .Y(n355), .A0(n343), .A1(n344) );
  nor02 U380 ( .Y(n356), .A0(n342), .A1(n344) );
  nor02 U381 ( .Y(n357), .A0(n342), .A1(n343) );
  nor02 U382 ( .Y(n341), .A0(n357), .A1(n358) );
  nor02 U383 ( .Y(n359), .A0(A[11]), .A1(carry_11_) );
  inv01 U384 ( .Y(n346), .A(n359) );
  nor02 U385 ( .Y(n360), .A0(B[11]), .A1(carry_11_) );
  inv01 U386 ( .Y(n348), .A(n360) );
  nor02 U387 ( .Y(n361), .A0(B[11]), .A1(A[11]) );
  inv01 U388 ( .Y(n350), .A(n361) );
  nor02 U389 ( .Y(n362), .A0(n342), .A1(n343) );
  inv01 U390 ( .Y(n352), .A(n362) );
  nor02 U391 ( .Y(n363), .A0(n345), .A1(n347) );
  inv01 U392 ( .Y(n353), .A(n363) );
  nor02 U393 ( .Y(n364), .A0(n349), .A1(n351) );
  inv01 U394 ( .Y(n354), .A(n364) );
  nor02 U395 ( .Y(n365), .A0(n355), .A1(n356) );
  inv01 U396 ( .Y(n358), .A(n365) );
  inv01 U397 ( .Y(SUM[10]), .A(n366) );
  inv02 U398 ( .Y(carry_11_), .A(n367) );
  inv02 U399 ( .Y(n368), .A(B[10]) );
  inv02 U400 ( .Y(n369), .A(A[10]) );
  inv02 U401 ( .Y(n370), .A(carry_10_) );
  nor02 U402 ( .Y(n371), .A0(n368), .A1(n372) );
  nor02 U403 ( .Y(n373), .A0(n369), .A1(n374) );
  nor02 U404 ( .Y(n375), .A0(n370), .A1(n376) );
  nor02 U405 ( .Y(n377), .A0(n370), .A1(n378) );
  nor02 U406 ( .Y(n366), .A0(n379), .A1(n380) );
  nor02 U407 ( .Y(n381), .A0(n369), .A1(n370) );
  nor02 U408 ( .Y(n382), .A0(n368), .A1(n370) );
  nor02 U409 ( .Y(n383), .A0(n368), .A1(n369) );
  nor02 U410 ( .Y(n367), .A0(n383), .A1(n384) );
  nor02 U411 ( .Y(n385), .A0(A[10]), .A1(carry_10_) );
  inv01 U412 ( .Y(n372), .A(n385) );
  nor02 U413 ( .Y(n386), .A0(B[10]), .A1(carry_10_) );
  inv01 U414 ( .Y(n374), .A(n386) );
  nor02 U415 ( .Y(n387), .A0(B[10]), .A1(A[10]) );
  inv01 U416 ( .Y(n376), .A(n387) );
  nor02 U417 ( .Y(n388), .A0(n368), .A1(n369) );
  inv01 U418 ( .Y(n378), .A(n388) );
  nor02 U419 ( .Y(n389), .A0(n371), .A1(n373) );
  inv01 U420 ( .Y(n379), .A(n389) );
  nor02 U421 ( .Y(n390), .A0(n375), .A1(n377) );
  inv01 U422 ( .Y(n380), .A(n390) );
  nor02 U423 ( .Y(n391), .A0(n381), .A1(n382) );
  inv01 U424 ( .Y(n384), .A(n391) );
  inv01 U425 ( .Y(SUM[9]), .A(n392) );
  inv02 U426 ( .Y(carry_10_), .A(n393) );
  inv02 U427 ( .Y(n394), .A(B[9]) );
  inv02 U428 ( .Y(n395), .A(A[9]) );
  inv02 U429 ( .Y(n396), .A(carry_9_) );
  nor02 U430 ( .Y(n397), .A0(n394), .A1(n398) );
  nor02 U431 ( .Y(n399), .A0(n395), .A1(n400) );
  nor02 U432 ( .Y(n401), .A0(n396), .A1(n402) );
  nor02 U433 ( .Y(n403), .A0(n396), .A1(n404) );
  nor02 U434 ( .Y(n392), .A0(n405), .A1(n406) );
  nor02 U435 ( .Y(n407), .A0(n395), .A1(n396) );
  nor02 U436 ( .Y(n408), .A0(n394), .A1(n396) );
  nor02 U437 ( .Y(n409), .A0(n394), .A1(n395) );
  nor02 U438 ( .Y(n393), .A0(n409), .A1(n410) );
  nor02 U439 ( .Y(n411), .A0(A[9]), .A1(carry_9_) );
  inv01 U440 ( .Y(n398), .A(n411) );
  nor02 U441 ( .Y(n412), .A0(B[9]), .A1(carry_9_) );
  inv01 U442 ( .Y(n400), .A(n412) );
  nor02 U443 ( .Y(n413), .A0(B[9]), .A1(A[9]) );
  inv01 U444 ( .Y(n402), .A(n413) );
  nor02 U445 ( .Y(n414), .A0(n394), .A1(n395) );
  inv01 U446 ( .Y(n404), .A(n414) );
  nor02 U447 ( .Y(n415), .A0(n397), .A1(n399) );
  inv01 U448 ( .Y(n405), .A(n415) );
  nor02 U449 ( .Y(n416), .A0(n401), .A1(n403) );
  inv01 U450 ( .Y(n406), .A(n416) );
  nor02 U451 ( .Y(n417), .A0(n407), .A1(n408) );
  inv01 U452 ( .Y(n410), .A(n417) );
  inv01 U453 ( .Y(SUM[8]), .A(n418) );
  inv02 U454 ( .Y(carry_9_), .A(n419) );
  inv02 U455 ( .Y(n420), .A(B[8]) );
  inv02 U456 ( .Y(n421), .A(A[8]) );
  inv02 U457 ( .Y(n422), .A(carry_8_) );
  nor02 U458 ( .Y(n423), .A0(n420), .A1(n424) );
  nor02 U459 ( .Y(n425), .A0(n421), .A1(n426) );
  nor02 U460 ( .Y(n427), .A0(n422), .A1(n428) );
  nor02 U461 ( .Y(n429), .A0(n422), .A1(n430) );
  nor02 U462 ( .Y(n418), .A0(n431), .A1(n432) );
  nor02 U463 ( .Y(n433), .A0(n421), .A1(n422) );
  nor02 U464 ( .Y(n434), .A0(n420), .A1(n422) );
  nor02 U465 ( .Y(n435), .A0(n420), .A1(n421) );
  nor02 U466 ( .Y(n419), .A0(n435), .A1(n436) );
  nor02 U467 ( .Y(n437), .A0(A[8]), .A1(carry_8_) );
  inv01 U468 ( .Y(n424), .A(n437) );
  nor02 U469 ( .Y(n438), .A0(B[8]), .A1(carry_8_) );
  inv01 U470 ( .Y(n426), .A(n438) );
  nor02 U471 ( .Y(n439), .A0(B[8]), .A1(A[8]) );
  inv01 U472 ( .Y(n428), .A(n439) );
  nor02 U473 ( .Y(n440), .A0(n420), .A1(n421) );
  inv01 U474 ( .Y(n430), .A(n440) );
  nor02 U475 ( .Y(n441), .A0(n423), .A1(n425) );
  inv01 U476 ( .Y(n431), .A(n441) );
  nor02 U477 ( .Y(n442), .A0(n427), .A1(n429) );
  inv01 U478 ( .Y(n432), .A(n442) );
  nor02 U479 ( .Y(n443), .A0(n433), .A1(n434) );
  inv01 U480 ( .Y(n436), .A(n443) );
  inv01 U481 ( .Y(SUM[7]), .A(n444) );
  inv02 U482 ( .Y(carry_8_), .A(n445) );
  inv02 U483 ( .Y(n446), .A(B[7]) );
  inv02 U484 ( .Y(n447), .A(A[7]) );
  inv02 U485 ( .Y(n448), .A(carry_7_) );
  nor02 U486 ( .Y(n449), .A0(n446), .A1(n450) );
  nor02 U487 ( .Y(n451), .A0(n447), .A1(n452) );
  nor02 U488 ( .Y(n453), .A0(n448), .A1(n454) );
  nor02 U489 ( .Y(n455), .A0(n448), .A1(n456) );
  nor02 U490 ( .Y(n444), .A0(n457), .A1(n458) );
  nor02 U491 ( .Y(n459), .A0(n447), .A1(n448) );
  nor02 U492 ( .Y(n460), .A0(n446), .A1(n448) );
  nor02 U493 ( .Y(n461), .A0(n446), .A1(n447) );
  nor02 U494 ( .Y(n445), .A0(n461), .A1(n462) );
  nor02 U495 ( .Y(n463), .A0(A[7]), .A1(carry_7_) );
  inv01 U496 ( .Y(n450), .A(n463) );
  nor02 U497 ( .Y(n464), .A0(B[7]), .A1(carry_7_) );
  inv01 U498 ( .Y(n452), .A(n464) );
  nor02 U499 ( .Y(n465), .A0(B[7]), .A1(A[7]) );
  inv01 U500 ( .Y(n454), .A(n465) );
  nor02 U501 ( .Y(n466), .A0(n446), .A1(n447) );
  inv01 U502 ( .Y(n456), .A(n466) );
  nor02 U503 ( .Y(n467), .A0(n449), .A1(n451) );
  inv01 U504 ( .Y(n457), .A(n467) );
  nor02 U505 ( .Y(n468), .A0(n453), .A1(n455) );
  inv01 U506 ( .Y(n458), .A(n468) );
  nor02 U507 ( .Y(n469), .A0(n459), .A1(n460) );
  inv01 U508 ( .Y(n462), .A(n469) );
  inv01 U509 ( .Y(SUM[6]), .A(n470) );
  inv02 U510 ( .Y(carry_7_), .A(n471) );
  inv02 U511 ( .Y(n472), .A(B[6]) );
  inv02 U512 ( .Y(n473), .A(A[6]) );
  inv02 U513 ( .Y(n474), .A(carry_6_) );
  nor02 U514 ( .Y(n475), .A0(n472), .A1(n476) );
  nor02 U515 ( .Y(n477), .A0(n473), .A1(n478) );
  nor02 U516 ( .Y(n479), .A0(n474), .A1(n480) );
  nor02 U517 ( .Y(n481), .A0(n474), .A1(n482) );
  nor02 U518 ( .Y(n470), .A0(n483), .A1(n484) );
  nor02 U519 ( .Y(n485), .A0(n473), .A1(n474) );
  nor02 U520 ( .Y(n486), .A0(n472), .A1(n474) );
  nor02 U521 ( .Y(n487), .A0(n472), .A1(n473) );
  nor02 U522 ( .Y(n471), .A0(n487), .A1(n488) );
  nor02 U523 ( .Y(n489), .A0(A[6]), .A1(carry_6_) );
  inv01 U524 ( .Y(n476), .A(n489) );
  nor02 U525 ( .Y(n490), .A0(B[6]), .A1(carry_6_) );
  inv01 U526 ( .Y(n478), .A(n490) );
  nor02 U527 ( .Y(n491), .A0(B[6]), .A1(A[6]) );
  inv01 U528 ( .Y(n480), .A(n491) );
  nor02 U529 ( .Y(n492), .A0(n472), .A1(n473) );
  inv01 U530 ( .Y(n482), .A(n492) );
  nor02 U531 ( .Y(n493), .A0(n475), .A1(n477) );
  inv01 U532 ( .Y(n483), .A(n493) );
  nor02 U533 ( .Y(n494), .A0(n479), .A1(n481) );
  inv01 U534 ( .Y(n484), .A(n494) );
  nor02 U535 ( .Y(n495), .A0(n485), .A1(n486) );
  inv01 U536 ( .Y(n488), .A(n495) );
  inv01 U537 ( .Y(SUM[5]), .A(n496) );
  inv02 U538 ( .Y(carry_6_), .A(n497) );
  inv02 U539 ( .Y(n498), .A(B[5]) );
  inv02 U540 ( .Y(n499), .A(A[5]) );
  inv02 U541 ( .Y(n500), .A(carry_5_) );
  nor02 U542 ( .Y(n501), .A0(n498), .A1(n502) );
  nor02 U543 ( .Y(n503), .A0(n499), .A1(n504) );
  nor02 U544 ( .Y(n505), .A0(n500), .A1(n506) );
  nor02 U545 ( .Y(n507), .A0(n500), .A1(n508) );
  nor02 U546 ( .Y(n496), .A0(n509), .A1(n510) );
  nor02 U547 ( .Y(n511), .A0(n499), .A1(n500) );
  nor02 U548 ( .Y(n512), .A0(n498), .A1(n500) );
  nor02 U549 ( .Y(n513), .A0(n498), .A1(n499) );
  nor02 U550 ( .Y(n497), .A0(n513), .A1(n514) );
  nor02 U551 ( .Y(n515), .A0(A[5]), .A1(carry_5_) );
  inv01 U552 ( .Y(n502), .A(n515) );
  nor02 U553 ( .Y(n516), .A0(B[5]), .A1(carry_5_) );
  inv01 U554 ( .Y(n504), .A(n516) );
  nor02 U555 ( .Y(n517), .A0(B[5]), .A1(A[5]) );
  inv01 U556 ( .Y(n506), .A(n517) );
  nor02 U557 ( .Y(n518), .A0(n498), .A1(n499) );
  inv01 U558 ( .Y(n508), .A(n518) );
  nor02 U559 ( .Y(n519), .A0(n501), .A1(n503) );
  inv01 U560 ( .Y(n509), .A(n519) );
  nor02 U561 ( .Y(n520), .A0(n505), .A1(n507) );
  inv01 U562 ( .Y(n510), .A(n520) );
  nor02 U563 ( .Y(n521), .A0(n511), .A1(n512) );
  inv01 U564 ( .Y(n514), .A(n521) );
  inv01 U565 ( .Y(SUM[4]), .A(n522) );
  inv02 U566 ( .Y(carry_5_), .A(n523) );
  inv02 U567 ( .Y(n524), .A(B[4]) );
  inv02 U568 ( .Y(n525), .A(A[4]) );
  inv02 U569 ( .Y(n526), .A(carry_4_) );
  nor02 U570 ( .Y(n527), .A0(n524), .A1(n528) );
  nor02 U571 ( .Y(n529), .A0(n525), .A1(n530) );
  nor02 U572 ( .Y(n531), .A0(n526), .A1(n532) );
  nor02 U573 ( .Y(n533), .A0(n526), .A1(n534) );
  nor02 U574 ( .Y(n522), .A0(n535), .A1(n536) );
  nor02 U575 ( .Y(n537), .A0(n525), .A1(n526) );
  nor02 U576 ( .Y(n538), .A0(n524), .A1(n526) );
  nor02 U577 ( .Y(n539), .A0(n524), .A1(n525) );
  nor02 U578 ( .Y(n523), .A0(n539), .A1(n540) );
  nor02 U579 ( .Y(n541), .A0(A[4]), .A1(carry_4_) );
  inv01 U580 ( .Y(n528), .A(n541) );
  nor02 U581 ( .Y(n542), .A0(B[4]), .A1(carry_4_) );
  inv01 U582 ( .Y(n530), .A(n542) );
  nor02 U583 ( .Y(n543), .A0(B[4]), .A1(A[4]) );
  inv01 U584 ( .Y(n532), .A(n543) );
  nor02 U585 ( .Y(n544), .A0(n524), .A1(n525) );
  inv01 U586 ( .Y(n534), .A(n544) );
  nor02 U587 ( .Y(n545), .A0(n527), .A1(n529) );
  inv01 U588 ( .Y(n535), .A(n545) );
  nor02 U589 ( .Y(n546), .A0(n531), .A1(n533) );
  inv01 U590 ( .Y(n536), .A(n546) );
  nor02 U591 ( .Y(n547), .A0(n537), .A1(n538) );
  inv01 U592 ( .Y(n540), .A(n547) );
  inv01 U593 ( .Y(SUM[3]), .A(n548) );
  inv02 U594 ( .Y(carry_4_), .A(n549) );
  inv02 U595 ( .Y(n550), .A(B[3]) );
  inv02 U596 ( .Y(n551), .A(A[3]) );
  inv02 U597 ( .Y(n552), .A(carry_3_) );
  nor02 U598 ( .Y(n553), .A0(n550), .A1(n554) );
  nor02 U599 ( .Y(n555), .A0(n551), .A1(n556) );
  nor02 U600 ( .Y(n557), .A0(n552), .A1(n558) );
  nor02 U601 ( .Y(n559), .A0(n552), .A1(n560) );
  nor02 U602 ( .Y(n548), .A0(n561), .A1(n562) );
  nor02 U603 ( .Y(n563), .A0(n551), .A1(n552) );
  nor02 U604 ( .Y(n564), .A0(n550), .A1(n552) );
  nor02 U605 ( .Y(n565), .A0(n550), .A1(n551) );
  nor02 U606 ( .Y(n549), .A0(n565), .A1(n566) );
  nor02 U607 ( .Y(n567), .A0(A[3]), .A1(carry_3_) );
  inv01 U608 ( .Y(n554), .A(n567) );
  nor02 U609 ( .Y(n568), .A0(B[3]), .A1(carry_3_) );
  inv01 U610 ( .Y(n556), .A(n568) );
  nor02 U611 ( .Y(n569), .A0(B[3]), .A1(A[3]) );
  inv01 U612 ( .Y(n558), .A(n569) );
  nor02 U613 ( .Y(n570), .A0(n550), .A1(n551) );
  inv01 U614 ( .Y(n560), .A(n570) );
  nor02 U615 ( .Y(n571), .A0(n553), .A1(n555) );
  inv01 U616 ( .Y(n561), .A(n571) );
  nor02 U617 ( .Y(n572), .A0(n557), .A1(n559) );
  inv01 U618 ( .Y(n562), .A(n572) );
  nor02 U619 ( .Y(n573), .A0(n563), .A1(n564) );
  inv01 U620 ( .Y(n566), .A(n573) );
  inv01 U621 ( .Y(SUM[2]), .A(n574) );
  inv02 U622 ( .Y(carry_3_), .A(n575) );
  inv02 U623 ( .Y(n576), .A(B[2]) );
  inv02 U624 ( .Y(n577), .A(A[2]) );
  inv02 U625 ( .Y(n578), .A(carry_2_) );
  nor02 U626 ( .Y(n579), .A0(n576), .A1(n580) );
  nor02 U627 ( .Y(n581), .A0(n577), .A1(n582) );
  nor02 U628 ( .Y(n583), .A0(n578), .A1(n584) );
  nor02 U629 ( .Y(n585), .A0(n578), .A1(n586) );
  nor02 U630 ( .Y(n574), .A0(n587), .A1(n588) );
  nor02 U631 ( .Y(n589), .A0(n577), .A1(n578) );
  nor02 U632 ( .Y(n590), .A0(n576), .A1(n578) );
  nor02 U633 ( .Y(n591), .A0(n576), .A1(n577) );
  nor02 U634 ( .Y(n575), .A0(n591), .A1(n592) );
  nor02 U635 ( .Y(n593), .A0(A[2]), .A1(carry_2_) );
  inv01 U636 ( .Y(n580), .A(n593) );
  nor02 U637 ( .Y(n594), .A0(B[2]), .A1(carry_2_) );
  inv01 U638 ( .Y(n582), .A(n594) );
  nor02 U639 ( .Y(n595), .A0(B[2]), .A1(A[2]) );
  inv01 U640 ( .Y(n584), .A(n595) );
  nor02 U641 ( .Y(n596), .A0(n576), .A1(n577) );
  inv01 U642 ( .Y(n586), .A(n596) );
  nor02 U643 ( .Y(n597), .A0(n579), .A1(n581) );
  inv01 U644 ( .Y(n587), .A(n597) );
  nor02 U645 ( .Y(n598), .A0(n583), .A1(n585) );
  inv01 U646 ( .Y(n588), .A(n598) );
  nor02 U647 ( .Y(n599), .A0(n589), .A1(n590) );
  inv01 U648 ( .Y(n592), .A(n599) );
  inv01 U649 ( .Y(SUM[1]), .A(n600) );
  inv02 U650 ( .Y(carry_2_), .A(n601) );
  inv02 U651 ( .Y(n602), .A(B[1]) );
  inv02 U652 ( .Y(n603), .A(A[1]) );
  inv02 U653 ( .Y(n604), .A(carry_1_) );
  nor02 U654 ( .Y(n605), .A0(n602), .A1(n606) );
  nor02 U655 ( .Y(n607), .A0(n603), .A1(n608) );
  nor02 U656 ( .Y(n609), .A0(n604), .A1(n610) );
  nor02 U657 ( .Y(n611), .A0(n604), .A1(n612) );
  nor02 U658 ( .Y(n600), .A0(n613), .A1(n614) );
  nor02 U659 ( .Y(n615), .A0(n603), .A1(n604) );
  nor02 U660 ( .Y(n616), .A0(n602), .A1(n604) );
  nor02 U661 ( .Y(n617), .A0(n602), .A1(n603) );
  nor02 U662 ( .Y(n601), .A0(n617), .A1(n618) );
  nor02 U663 ( .Y(n619), .A0(A[1]), .A1(n1) );
  inv01 U664 ( .Y(n606), .A(n619) );
  nor02 U665 ( .Y(n620), .A0(B[1]), .A1(n1) );
  inv01 U666 ( .Y(n608), .A(n620) );
  nor02 U667 ( .Y(n621), .A0(B[1]), .A1(A[1]) );
  inv01 U668 ( .Y(n610), .A(n621) );
  nor02 U669 ( .Y(n622), .A0(n602), .A1(n603) );
  inv01 U670 ( .Y(n612), .A(n622) );
  nor02 U671 ( .Y(n623), .A0(n605), .A1(n607) );
  inv01 U672 ( .Y(n613), .A(n623) );
  nor02 U673 ( .Y(n624), .A0(n609), .A1(n611) );
  inv01 U674 ( .Y(n614), .A(n624) );
  nor02 U675 ( .Y(n625), .A0(n615), .A1(n616) );
  inv01 U676 ( .Y(n618), .A(n625) );
  and02 U677 ( .Y(carry_1_), .A0(A[0]), .A1(B[0]) );
  xor2 U678 ( .Y(SUM[0]), .A0(B[0]), .A1(A[0]) );
  fadd1 U1_25 ( .S(SUM[25]), .A(A[25]), .B(B[25]), .CI(carry_25_) );
endmodule


module sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_sub_26_0 ( A, B, CI, DIFF, CO );
  input [25:0] A;
  input [25:0] B;
  output [25:0] DIFF;
  input CI;
  output CO;
  wire   carry_25_, carry_24_, carry_23_, carry_22_, carry_21_, carry_20_,
         carry_19_, carry_18_, carry_17_, carry_16_, carry_15_, carry_14_,
         carry_13_, carry_12_, carry_11_, carry_10_, carry_9_, carry_8_,
         carry_7_, carry_6_, carry_5_, carry_4_, carry_3_, carry_2_, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580;
  wire   [25:0] B_not;

  inv02 U6 ( .Y(B_not[25]), .A(B[25]) );
  nor02 U7 ( .Y(n5), .A0(B_not[0]), .A1(A[0]) );
  inv02 U8 ( .Y(n6), .A(n5) );
  buf02 U9 ( .Y(n7), .A(carry_25_) );
  inv01 U10 ( .Y(DIFF[23]), .A(n8) );
  inv02 U11 ( .Y(carry_24_), .A(n9) );
  inv02 U12 ( .Y(n10), .A(B_not[23]) );
  inv02 U13 ( .Y(n11), .A(A[23]) );
  inv02 U14 ( .Y(n12), .A(carry_23_) );
  nor02 U15 ( .Y(n13), .A0(n10), .A1(n14) );
  nor02 U16 ( .Y(n15), .A0(n11), .A1(n16) );
  nor02 U17 ( .Y(n17), .A0(n12), .A1(n18) );
  nor02 U18 ( .Y(n19), .A0(n12), .A1(n20) );
  nor02 U19 ( .Y(n8), .A0(n21), .A1(n22) );
  nor02 U20 ( .Y(n23), .A0(n11), .A1(n12) );
  nor02 U21 ( .Y(n24), .A0(n10), .A1(n12) );
  nor02 U22 ( .Y(n25), .A0(n10), .A1(n11) );
  nor02 U23 ( .Y(n9), .A0(n25), .A1(n26) );
  nor02 U24 ( .Y(n27), .A0(A[23]), .A1(carry_23_) );
  inv01 U25 ( .Y(n14), .A(n27) );
  nor02 U26 ( .Y(n28), .A0(B_not[23]), .A1(carry_23_) );
  inv01 U27 ( .Y(n16), .A(n28) );
  nor02 U28 ( .Y(n29), .A0(B_not[23]), .A1(A[23]) );
  inv01 U29 ( .Y(n18), .A(n29) );
  nor02 U30 ( .Y(n30), .A0(n10), .A1(n11) );
  inv01 U31 ( .Y(n20), .A(n30) );
  nor02 U32 ( .Y(n31), .A0(n13), .A1(n15) );
  inv01 U33 ( .Y(n21), .A(n31) );
  nor02 U34 ( .Y(n32), .A0(n17), .A1(n19) );
  inv01 U35 ( .Y(n22), .A(n32) );
  nor02 U36 ( .Y(n33), .A0(n23), .A1(n24) );
  inv01 U37 ( .Y(n26), .A(n33) );
  inv02 U38 ( .Y(B_not[23]), .A(B[23]) );
  inv01 U39 ( .Y(DIFF[22]), .A(n34) );
  inv02 U40 ( .Y(carry_23_), .A(n35) );
  inv02 U41 ( .Y(n36), .A(B_not[22]) );
  inv02 U42 ( .Y(n37), .A(A[22]) );
  inv02 U43 ( .Y(n38), .A(carry_22_) );
  nor02 U44 ( .Y(n39), .A0(n36), .A1(n40) );
  nor02 U45 ( .Y(n41), .A0(n37), .A1(n42) );
  nor02 U46 ( .Y(n43), .A0(n38), .A1(n44) );
  nor02 U47 ( .Y(n45), .A0(n38), .A1(n46) );
  nor02 U48 ( .Y(n34), .A0(n47), .A1(n48) );
  nor02 U49 ( .Y(n49), .A0(n37), .A1(n38) );
  nor02 U50 ( .Y(n50), .A0(n36), .A1(n38) );
  nor02 U51 ( .Y(n51), .A0(n36), .A1(n37) );
  nor02 U52 ( .Y(n35), .A0(n51), .A1(n52) );
  nor02 U53 ( .Y(n53), .A0(A[22]), .A1(carry_22_) );
  inv01 U54 ( .Y(n40), .A(n53) );
  nor02 U55 ( .Y(n54), .A0(B_not[22]), .A1(carry_22_) );
  inv01 U56 ( .Y(n42), .A(n54) );
  nor02 U57 ( .Y(n55), .A0(B_not[22]), .A1(A[22]) );
  inv01 U58 ( .Y(n44), .A(n55) );
  nor02 U59 ( .Y(n56), .A0(n36), .A1(n37) );
  inv01 U60 ( .Y(n46), .A(n56) );
  nor02 U61 ( .Y(n57), .A0(n39), .A1(n41) );
  inv01 U62 ( .Y(n47), .A(n57) );
  nor02 U63 ( .Y(n58), .A0(n43), .A1(n45) );
  inv01 U64 ( .Y(n48), .A(n58) );
  nor02 U65 ( .Y(n59), .A0(n49), .A1(n50) );
  inv01 U66 ( .Y(n52), .A(n59) );
  inv02 U67 ( .Y(B_not[22]), .A(B[22]) );
  inv01 U68 ( .Y(DIFF[21]), .A(n60) );
  inv02 U69 ( .Y(carry_22_), .A(n61) );
  inv02 U70 ( .Y(n62), .A(B_not[21]) );
  inv02 U71 ( .Y(n63), .A(A[21]) );
  inv02 U72 ( .Y(n64), .A(carry_21_) );
  nor02 U73 ( .Y(n65), .A0(n62), .A1(n66) );
  nor02 U74 ( .Y(n67), .A0(n63), .A1(n68) );
  nor02 U75 ( .Y(n69), .A0(n64), .A1(n70) );
  nor02 U76 ( .Y(n71), .A0(n64), .A1(n72) );
  nor02 U77 ( .Y(n60), .A0(n73), .A1(n74) );
  nor02 U78 ( .Y(n75), .A0(n63), .A1(n64) );
  nor02 U79 ( .Y(n76), .A0(n62), .A1(n64) );
  nor02 U80 ( .Y(n77), .A0(n62), .A1(n63) );
  nor02 U81 ( .Y(n61), .A0(n77), .A1(n78) );
  nor02 U82 ( .Y(n79), .A0(A[21]), .A1(carry_21_) );
  inv01 U83 ( .Y(n66), .A(n79) );
  nor02 U84 ( .Y(n80), .A0(B_not[21]), .A1(carry_21_) );
  inv01 U85 ( .Y(n68), .A(n80) );
  nor02 U86 ( .Y(n81), .A0(B_not[21]), .A1(A[21]) );
  inv01 U87 ( .Y(n70), .A(n81) );
  nor02 U88 ( .Y(n82), .A0(n62), .A1(n63) );
  inv01 U89 ( .Y(n72), .A(n82) );
  nor02 U90 ( .Y(n83), .A0(n65), .A1(n67) );
  inv01 U91 ( .Y(n73), .A(n83) );
  nor02 U92 ( .Y(n84), .A0(n69), .A1(n71) );
  inv01 U93 ( .Y(n74), .A(n84) );
  nor02 U94 ( .Y(n85), .A0(n75), .A1(n76) );
  inv01 U95 ( .Y(n78), .A(n85) );
  inv02 U96 ( .Y(B_not[21]), .A(B[21]) );
  inv01 U97 ( .Y(DIFF[20]), .A(n86) );
  inv02 U98 ( .Y(carry_21_), .A(n87) );
  inv02 U99 ( .Y(n88), .A(B_not[20]) );
  inv02 U100 ( .Y(n89), .A(A[20]) );
  inv02 U101 ( .Y(n90), .A(carry_20_) );
  nor02 U102 ( .Y(n91), .A0(n88), .A1(n92) );
  nor02 U103 ( .Y(n93), .A0(n89), .A1(n94) );
  nor02 U104 ( .Y(n95), .A0(n90), .A1(n96) );
  nor02 U105 ( .Y(n97), .A0(n90), .A1(n98) );
  nor02 U106 ( .Y(n86), .A0(n99), .A1(n100) );
  nor02 U107 ( .Y(n101), .A0(n89), .A1(n90) );
  nor02 U108 ( .Y(n102), .A0(n88), .A1(n90) );
  nor02 U109 ( .Y(n103), .A0(n88), .A1(n89) );
  nor02 U110 ( .Y(n87), .A0(n103), .A1(n104) );
  nor02 U111 ( .Y(n105), .A0(A[20]), .A1(carry_20_) );
  inv01 U112 ( .Y(n92), .A(n105) );
  nor02 U113 ( .Y(n106), .A0(B_not[20]), .A1(carry_20_) );
  inv01 U114 ( .Y(n94), .A(n106) );
  nor02 U115 ( .Y(n107), .A0(B_not[20]), .A1(A[20]) );
  inv01 U116 ( .Y(n96), .A(n107) );
  nor02 U117 ( .Y(n108), .A0(n88), .A1(n89) );
  inv01 U118 ( .Y(n98), .A(n108) );
  nor02 U119 ( .Y(n109), .A0(n91), .A1(n93) );
  inv01 U120 ( .Y(n99), .A(n109) );
  nor02 U121 ( .Y(n110), .A0(n95), .A1(n97) );
  inv01 U122 ( .Y(n100), .A(n110) );
  nor02 U123 ( .Y(n111), .A0(n101), .A1(n102) );
  inv01 U124 ( .Y(n104), .A(n111) );
  inv02 U125 ( .Y(B_not[20]), .A(B[20]) );
  inv01 U126 ( .Y(DIFF[19]), .A(n112) );
  inv02 U127 ( .Y(carry_20_), .A(n113) );
  inv02 U128 ( .Y(n114), .A(B_not[19]) );
  inv02 U129 ( .Y(n115), .A(A[19]) );
  inv02 U130 ( .Y(n116), .A(carry_19_) );
  nor02 U131 ( .Y(n117), .A0(n114), .A1(n118) );
  nor02 U132 ( .Y(n119), .A0(n115), .A1(n120) );
  nor02 U133 ( .Y(n121), .A0(n116), .A1(n122) );
  nor02 U134 ( .Y(n123), .A0(n116), .A1(n124) );
  nor02 U135 ( .Y(n112), .A0(n125), .A1(n126) );
  nor02 U136 ( .Y(n127), .A0(n115), .A1(n116) );
  nor02 U137 ( .Y(n128), .A0(n114), .A1(n116) );
  nor02 U138 ( .Y(n129), .A0(n114), .A1(n115) );
  nor02 U139 ( .Y(n113), .A0(n129), .A1(n130) );
  nor02 U140 ( .Y(n131), .A0(A[19]), .A1(carry_19_) );
  inv01 U141 ( .Y(n118), .A(n131) );
  nor02 U142 ( .Y(n132), .A0(B_not[19]), .A1(carry_19_) );
  inv01 U143 ( .Y(n120), .A(n132) );
  nor02 U144 ( .Y(n133), .A0(B_not[19]), .A1(A[19]) );
  inv01 U145 ( .Y(n122), .A(n133) );
  nor02 U146 ( .Y(n134), .A0(n114), .A1(n115) );
  inv01 U147 ( .Y(n124), .A(n134) );
  nor02 U148 ( .Y(n135), .A0(n117), .A1(n119) );
  inv01 U149 ( .Y(n125), .A(n135) );
  nor02 U150 ( .Y(n136), .A0(n121), .A1(n123) );
  inv01 U151 ( .Y(n126), .A(n136) );
  nor02 U152 ( .Y(n137), .A0(n127), .A1(n128) );
  inv01 U153 ( .Y(n130), .A(n137) );
  inv02 U154 ( .Y(B_not[19]), .A(B[19]) );
  inv01 U155 ( .Y(DIFF[18]), .A(n138) );
  inv02 U156 ( .Y(carry_19_), .A(n139) );
  inv02 U157 ( .Y(n140), .A(B_not[18]) );
  inv02 U158 ( .Y(n141), .A(A[18]) );
  inv02 U159 ( .Y(n142), .A(carry_18_) );
  nor02 U160 ( .Y(n143), .A0(n140), .A1(n144) );
  nor02 U161 ( .Y(n145), .A0(n141), .A1(n146) );
  nor02 U162 ( .Y(n147), .A0(n142), .A1(n148) );
  nor02 U163 ( .Y(n149), .A0(n142), .A1(n150) );
  nor02 U164 ( .Y(n138), .A0(n151), .A1(n152) );
  nor02 U165 ( .Y(n153), .A0(n141), .A1(n142) );
  nor02 U166 ( .Y(n154), .A0(n140), .A1(n142) );
  nor02 U167 ( .Y(n155), .A0(n140), .A1(n141) );
  nor02 U168 ( .Y(n139), .A0(n155), .A1(n156) );
  nor02 U169 ( .Y(n157), .A0(A[18]), .A1(carry_18_) );
  inv01 U170 ( .Y(n144), .A(n157) );
  nor02 U171 ( .Y(n158), .A0(B_not[18]), .A1(carry_18_) );
  inv01 U172 ( .Y(n146), .A(n158) );
  nor02 U173 ( .Y(n159), .A0(B_not[18]), .A1(A[18]) );
  inv01 U174 ( .Y(n148), .A(n159) );
  nor02 U175 ( .Y(n160), .A0(n140), .A1(n141) );
  inv01 U176 ( .Y(n150), .A(n160) );
  nor02 U177 ( .Y(n161), .A0(n143), .A1(n145) );
  inv01 U178 ( .Y(n151), .A(n161) );
  nor02 U179 ( .Y(n162), .A0(n147), .A1(n149) );
  inv01 U180 ( .Y(n152), .A(n162) );
  nor02 U181 ( .Y(n163), .A0(n153), .A1(n154) );
  inv01 U182 ( .Y(n156), .A(n163) );
  inv02 U183 ( .Y(B_not[18]), .A(B[18]) );
  inv01 U184 ( .Y(DIFF[17]), .A(n164) );
  inv02 U185 ( .Y(carry_18_), .A(n165) );
  inv02 U186 ( .Y(n166), .A(B_not[17]) );
  inv02 U187 ( .Y(n167), .A(A[17]) );
  inv02 U188 ( .Y(n168), .A(carry_17_) );
  nor02 U189 ( .Y(n169), .A0(n166), .A1(n170) );
  nor02 U190 ( .Y(n171), .A0(n167), .A1(n172) );
  nor02 U191 ( .Y(n173), .A0(n168), .A1(n174) );
  nor02 U192 ( .Y(n175), .A0(n168), .A1(n176) );
  nor02 U193 ( .Y(n164), .A0(n177), .A1(n178) );
  nor02 U194 ( .Y(n179), .A0(n167), .A1(n168) );
  nor02 U195 ( .Y(n180), .A0(n166), .A1(n168) );
  nor02 U196 ( .Y(n181), .A0(n166), .A1(n167) );
  nor02 U197 ( .Y(n165), .A0(n181), .A1(n182) );
  nor02 U198 ( .Y(n183), .A0(A[17]), .A1(carry_17_) );
  inv01 U199 ( .Y(n170), .A(n183) );
  nor02 U200 ( .Y(n184), .A0(B_not[17]), .A1(carry_17_) );
  inv01 U201 ( .Y(n172), .A(n184) );
  nor02 U202 ( .Y(n185), .A0(B_not[17]), .A1(A[17]) );
  inv01 U203 ( .Y(n174), .A(n185) );
  nor02 U204 ( .Y(n186), .A0(n166), .A1(n167) );
  inv01 U205 ( .Y(n176), .A(n186) );
  nor02 U206 ( .Y(n187), .A0(n169), .A1(n171) );
  inv01 U207 ( .Y(n177), .A(n187) );
  nor02 U208 ( .Y(n188), .A0(n173), .A1(n175) );
  inv01 U209 ( .Y(n178), .A(n188) );
  nor02 U210 ( .Y(n189), .A0(n179), .A1(n180) );
  inv01 U211 ( .Y(n182), .A(n189) );
  inv02 U212 ( .Y(B_not[17]), .A(B[17]) );
  inv01 U213 ( .Y(DIFF[16]), .A(n190) );
  inv02 U214 ( .Y(carry_17_), .A(n191) );
  inv02 U215 ( .Y(n192), .A(B_not[16]) );
  inv02 U216 ( .Y(n193), .A(A[16]) );
  inv02 U217 ( .Y(n194), .A(carry_16_) );
  nor02 U218 ( .Y(n195), .A0(n192), .A1(n196) );
  nor02 U219 ( .Y(n197), .A0(n193), .A1(n198) );
  nor02 U220 ( .Y(n199), .A0(n194), .A1(n200) );
  nor02 U221 ( .Y(n201), .A0(n194), .A1(n202) );
  nor02 U222 ( .Y(n190), .A0(n203), .A1(n204) );
  nor02 U223 ( .Y(n205), .A0(n193), .A1(n194) );
  nor02 U224 ( .Y(n206), .A0(n192), .A1(n194) );
  nor02 U225 ( .Y(n207), .A0(n192), .A1(n193) );
  nor02 U226 ( .Y(n191), .A0(n207), .A1(n208) );
  nor02 U227 ( .Y(n209), .A0(A[16]), .A1(carry_16_) );
  inv01 U228 ( .Y(n196), .A(n209) );
  nor02 U229 ( .Y(n210), .A0(B_not[16]), .A1(carry_16_) );
  inv01 U230 ( .Y(n198), .A(n210) );
  nor02 U231 ( .Y(n211), .A0(B_not[16]), .A1(A[16]) );
  inv01 U232 ( .Y(n200), .A(n211) );
  nor02 U233 ( .Y(n212), .A0(n192), .A1(n193) );
  inv01 U234 ( .Y(n202), .A(n212) );
  nor02 U235 ( .Y(n213), .A0(n195), .A1(n197) );
  inv01 U236 ( .Y(n203), .A(n213) );
  nor02 U237 ( .Y(n214), .A0(n199), .A1(n201) );
  inv01 U238 ( .Y(n204), .A(n214) );
  nor02 U239 ( .Y(n215), .A0(n205), .A1(n206) );
  inv01 U240 ( .Y(n208), .A(n215) );
  inv02 U241 ( .Y(B_not[16]), .A(B[16]) );
  inv01 U242 ( .Y(DIFF[15]), .A(n216) );
  inv02 U243 ( .Y(carry_16_), .A(n217) );
  inv02 U244 ( .Y(n218), .A(B_not[15]) );
  inv02 U245 ( .Y(n219), .A(A[15]) );
  inv02 U246 ( .Y(n220), .A(carry_15_) );
  nor02 U247 ( .Y(n221), .A0(n218), .A1(n222) );
  nor02 U248 ( .Y(n223), .A0(n219), .A1(n224) );
  nor02 U249 ( .Y(n225), .A0(n220), .A1(n226) );
  nor02 U250 ( .Y(n227), .A0(n220), .A1(n228) );
  nor02 U251 ( .Y(n216), .A0(n229), .A1(n230) );
  nor02 U252 ( .Y(n231), .A0(n219), .A1(n220) );
  nor02 U253 ( .Y(n232), .A0(n218), .A1(n220) );
  nor02 U254 ( .Y(n233), .A0(n218), .A1(n219) );
  nor02 U255 ( .Y(n217), .A0(n233), .A1(n234) );
  nor02 U256 ( .Y(n235), .A0(A[15]), .A1(carry_15_) );
  inv01 U257 ( .Y(n222), .A(n235) );
  nor02 U258 ( .Y(n236), .A0(B_not[15]), .A1(carry_15_) );
  inv01 U259 ( .Y(n224), .A(n236) );
  nor02 U260 ( .Y(n237), .A0(B_not[15]), .A1(A[15]) );
  inv01 U261 ( .Y(n226), .A(n237) );
  nor02 U262 ( .Y(n238), .A0(n218), .A1(n219) );
  inv01 U263 ( .Y(n228), .A(n238) );
  nor02 U264 ( .Y(n239), .A0(n221), .A1(n223) );
  inv01 U265 ( .Y(n229), .A(n239) );
  nor02 U266 ( .Y(n240), .A0(n225), .A1(n227) );
  inv01 U267 ( .Y(n230), .A(n240) );
  nor02 U268 ( .Y(n241), .A0(n231), .A1(n232) );
  inv01 U269 ( .Y(n234), .A(n241) );
  inv02 U270 ( .Y(B_not[15]), .A(B[15]) );
  inv01 U271 ( .Y(DIFF[14]), .A(n242) );
  inv02 U272 ( .Y(carry_15_), .A(n243) );
  inv02 U273 ( .Y(n244), .A(B_not[14]) );
  inv02 U274 ( .Y(n245), .A(A[14]) );
  inv02 U275 ( .Y(n246), .A(carry_14_) );
  nor02 U276 ( .Y(n247), .A0(n244), .A1(n248) );
  nor02 U277 ( .Y(n249), .A0(n245), .A1(n250) );
  nor02 U278 ( .Y(n251), .A0(n246), .A1(n252) );
  nor02 U279 ( .Y(n253), .A0(n246), .A1(n254) );
  nor02 U280 ( .Y(n242), .A0(n255), .A1(n256) );
  nor02 U281 ( .Y(n257), .A0(n245), .A1(n246) );
  nor02 U282 ( .Y(n258), .A0(n244), .A1(n246) );
  nor02 U283 ( .Y(n259), .A0(n244), .A1(n245) );
  nor02 U284 ( .Y(n243), .A0(n259), .A1(n260) );
  nor02 U285 ( .Y(n261), .A0(A[14]), .A1(carry_14_) );
  inv01 U286 ( .Y(n248), .A(n261) );
  nor02 U287 ( .Y(n262), .A0(B_not[14]), .A1(carry_14_) );
  inv01 U288 ( .Y(n250), .A(n262) );
  nor02 U289 ( .Y(n263), .A0(B_not[14]), .A1(A[14]) );
  inv01 U290 ( .Y(n252), .A(n263) );
  nor02 U291 ( .Y(n264), .A0(n244), .A1(n245) );
  inv01 U292 ( .Y(n254), .A(n264) );
  nor02 U293 ( .Y(n265), .A0(n247), .A1(n249) );
  inv01 U294 ( .Y(n255), .A(n265) );
  nor02 U295 ( .Y(n266), .A0(n251), .A1(n253) );
  inv01 U296 ( .Y(n256), .A(n266) );
  nor02 U297 ( .Y(n267), .A0(n257), .A1(n258) );
  inv01 U298 ( .Y(n260), .A(n267) );
  inv02 U299 ( .Y(B_not[14]), .A(B[14]) );
  inv01 U300 ( .Y(DIFF[13]), .A(n268) );
  inv02 U301 ( .Y(carry_14_), .A(n269) );
  inv02 U302 ( .Y(n270), .A(B_not[13]) );
  inv02 U303 ( .Y(n271), .A(A[13]) );
  inv02 U304 ( .Y(n272), .A(carry_13_) );
  nor02 U305 ( .Y(n273), .A0(n270), .A1(n274) );
  nor02 U306 ( .Y(n275), .A0(n271), .A1(n276) );
  nor02 U307 ( .Y(n277), .A0(n272), .A1(n278) );
  nor02 U308 ( .Y(n279), .A0(n272), .A1(n280) );
  nor02 U309 ( .Y(n268), .A0(n281), .A1(n282) );
  nor02 U310 ( .Y(n283), .A0(n271), .A1(n272) );
  nor02 U311 ( .Y(n284), .A0(n270), .A1(n272) );
  nor02 U312 ( .Y(n285), .A0(n270), .A1(n271) );
  nor02 U313 ( .Y(n269), .A0(n285), .A1(n286) );
  nor02 U314 ( .Y(n287), .A0(A[13]), .A1(carry_13_) );
  inv01 U315 ( .Y(n274), .A(n287) );
  nor02 U316 ( .Y(n288), .A0(B_not[13]), .A1(carry_13_) );
  inv01 U317 ( .Y(n276), .A(n288) );
  nor02 U318 ( .Y(n289), .A0(B_not[13]), .A1(A[13]) );
  inv01 U319 ( .Y(n278), .A(n289) );
  nor02 U320 ( .Y(n290), .A0(n270), .A1(n271) );
  inv01 U321 ( .Y(n280), .A(n290) );
  nor02 U322 ( .Y(n291), .A0(n273), .A1(n275) );
  inv01 U323 ( .Y(n281), .A(n291) );
  nor02 U324 ( .Y(n292), .A0(n277), .A1(n279) );
  inv01 U325 ( .Y(n282), .A(n292) );
  nor02 U326 ( .Y(n293), .A0(n283), .A1(n284) );
  inv01 U327 ( .Y(n286), .A(n293) );
  inv02 U328 ( .Y(B_not[13]), .A(B[13]) );
  inv01 U329 ( .Y(DIFF[12]), .A(n294) );
  inv02 U330 ( .Y(carry_13_), .A(n295) );
  inv02 U331 ( .Y(n296), .A(B_not[12]) );
  inv02 U332 ( .Y(n297), .A(A[12]) );
  inv02 U333 ( .Y(n298), .A(carry_12_) );
  nor02 U334 ( .Y(n299), .A0(n296), .A1(n300) );
  nor02 U335 ( .Y(n301), .A0(n297), .A1(n302) );
  nor02 U336 ( .Y(n303), .A0(n298), .A1(n304) );
  nor02 U337 ( .Y(n305), .A0(n298), .A1(n306) );
  nor02 U338 ( .Y(n294), .A0(n307), .A1(n308) );
  nor02 U339 ( .Y(n309), .A0(n297), .A1(n298) );
  nor02 U340 ( .Y(n310), .A0(n296), .A1(n298) );
  nor02 U341 ( .Y(n311), .A0(n296), .A1(n297) );
  nor02 U342 ( .Y(n295), .A0(n311), .A1(n312) );
  nor02 U343 ( .Y(n313), .A0(A[12]), .A1(carry_12_) );
  inv01 U344 ( .Y(n300), .A(n313) );
  nor02 U345 ( .Y(n314), .A0(B_not[12]), .A1(carry_12_) );
  inv01 U346 ( .Y(n302), .A(n314) );
  nor02 U347 ( .Y(n315), .A0(B_not[12]), .A1(A[12]) );
  inv01 U348 ( .Y(n304), .A(n315) );
  nor02 U349 ( .Y(n316), .A0(n296), .A1(n297) );
  inv01 U350 ( .Y(n306), .A(n316) );
  nor02 U351 ( .Y(n317), .A0(n299), .A1(n301) );
  inv01 U352 ( .Y(n307), .A(n317) );
  nor02 U353 ( .Y(n318), .A0(n303), .A1(n305) );
  inv01 U354 ( .Y(n308), .A(n318) );
  nor02 U355 ( .Y(n319), .A0(n309), .A1(n310) );
  inv01 U356 ( .Y(n312), .A(n319) );
  inv02 U357 ( .Y(B_not[12]), .A(B[12]) );
  inv01 U358 ( .Y(DIFF[11]), .A(n320) );
  inv02 U359 ( .Y(carry_12_), .A(n321) );
  inv02 U360 ( .Y(n322), .A(B_not[11]) );
  inv02 U361 ( .Y(n323), .A(A[11]) );
  inv02 U362 ( .Y(n324), .A(carry_11_) );
  nor02 U363 ( .Y(n325), .A0(n322), .A1(n326) );
  nor02 U364 ( .Y(n327), .A0(n323), .A1(n328) );
  nor02 U365 ( .Y(n329), .A0(n324), .A1(n330) );
  nor02 U366 ( .Y(n331), .A0(n324), .A1(n332) );
  nor02 U367 ( .Y(n320), .A0(n333), .A1(n334) );
  nor02 U368 ( .Y(n335), .A0(n323), .A1(n324) );
  nor02 U369 ( .Y(n336), .A0(n322), .A1(n324) );
  nor02 U370 ( .Y(n337), .A0(n322), .A1(n323) );
  nor02 U371 ( .Y(n321), .A0(n337), .A1(n338) );
  nor02 U372 ( .Y(n339), .A0(A[11]), .A1(carry_11_) );
  inv01 U373 ( .Y(n326), .A(n339) );
  nor02 U374 ( .Y(n340), .A0(B_not[11]), .A1(carry_11_) );
  inv01 U375 ( .Y(n328), .A(n340) );
  nor02 U376 ( .Y(n341), .A0(B_not[11]), .A1(A[11]) );
  inv01 U377 ( .Y(n330), .A(n341) );
  nor02 U378 ( .Y(n342), .A0(n322), .A1(n323) );
  inv01 U379 ( .Y(n332), .A(n342) );
  nor02 U380 ( .Y(n343), .A0(n325), .A1(n327) );
  inv01 U381 ( .Y(n333), .A(n343) );
  nor02 U382 ( .Y(n344), .A0(n329), .A1(n331) );
  inv01 U383 ( .Y(n334), .A(n344) );
  nor02 U384 ( .Y(n345), .A0(n335), .A1(n336) );
  inv01 U385 ( .Y(n338), .A(n345) );
  inv02 U386 ( .Y(B_not[11]), .A(B[11]) );
  inv01 U387 ( .Y(DIFF[10]), .A(n346) );
  inv02 U388 ( .Y(carry_11_), .A(n347) );
  inv02 U389 ( .Y(n348), .A(B_not[10]) );
  inv02 U390 ( .Y(n349), .A(A[10]) );
  inv02 U391 ( .Y(n350), .A(carry_10_) );
  nor02 U392 ( .Y(n351), .A0(n348), .A1(n352) );
  nor02 U393 ( .Y(n353), .A0(n349), .A1(n354) );
  nor02 U394 ( .Y(n355), .A0(n350), .A1(n356) );
  nor02 U395 ( .Y(n357), .A0(n350), .A1(n358) );
  nor02 U396 ( .Y(n346), .A0(n359), .A1(n360) );
  nor02 U397 ( .Y(n361), .A0(n349), .A1(n350) );
  nor02 U398 ( .Y(n362), .A0(n348), .A1(n350) );
  nor02 U399 ( .Y(n363), .A0(n348), .A1(n349) );
  nor02 U400 ( .Y(n347), .A0(n363), .A1(n364) );
  nor02 U401 ( .Y(n365), .A0(A[10]), .A1(carry_10_) );
  inv01 U402 ( .Y(n352), .A(n365) );
  nor02 U403 ( .Y(n366), .A0(B_not[10]), .A1(carry_10_) );
  inv01 U404 ( .Y(n354), .A(n366) );
  nor02 U405 ( .Y(n367), .A0(B_not[10]), .A1(A[10]) );
  inv01 U406 ( .Y(n356), .A(n367) );
  nor02 U407 ( .Y(n368), .A0(n348), .A1(n349) );
  inv01 U408 ( .Y(n358), .A(n368) );
  nor02 U409 ( .Y(n369), .A0(n351), .A1(n353) );
  inv01 U410 ( .Y(n359), .A(n369) );
  nor02 U411 ( .Y(n370), .A0(n355), .A1(n357) );
  inv01 U412 ( .Y(n360), .A(n370) );
  nor02 U413 ( .Y(n371), .A0(n361), .A1(n362) );
  inv01 U414 ( .Y(n364), .A(n371) );
  inv02 U415 ( .Y(B_not[10]), .A(B[10]) );
  inv01 U416 ( .Y(DIFF[9]), .A(n372) );
  inv02 U417 ( .Y(carry_10_), .A(n373) );
  inv02 U418 ( .Y(n374), .A(B_not[9]) );
  inv02 U419 ( .Y(n375), .A(A[9]) );
  inv02 U420 ( .Y(n376), .A(carry_9_) );
  nor02 U421 ( .Y(n377), .A0(n374), .A1(n378) );
  nor02 U422 ( .Y(n379), .A0(n375), .A1(n380) );
  nor02 U423 ( .Y(n381), .A0(n376), .A1(n382) );
  nor02 U424 ( .Y(n383), .A0(n376), .A1(n384) );
  nor02 U425 ( .Y(n372), .A0(n385), .A1(n386) );
  nor02 U426 ( .Y(n387), .A0(n375), .A1(n376) );
  nor02 U427 ( .Y(n388), .A0(n374), .A1(n376) );
  nor02 U428 ( .Y(n389), .A0(n374), .A1(n375) );
  nor02 U429 ( .Y(n373), .A0(n389), .A1(n390) );
  nor02 U430 ( .Y(n391), .A0(A[9]), .A1(carry_9_) );
  inv01 U431 ( .Y(n378), .A(n391) );
  nor02 U432 ( .Y(n392), .A0(B_not[9]), .A1(carry_9_) );
  inv01 U433 ( .Y(n380), .A(n392) );
  nor02 U434 ( .Y(n393), .A0(B_not[9]), .A1(A[9]) );
  inv01 U435 ( .Y(n382), .A(n393) );
  nor02 U436 ( .Y(n394), .A0(n374), .A1(n375) );
  inv01 U437 ( .Y(n384), .A(n394) );
  nor02 U438 ( .Y(n395), .A0(n377), .A1(n379) );
  inv01 U439 ( .Y(n385), .A(n395) );
  nor02 U440 ( .Y(n396), .A0(n381), .A1(n383) );
  inv01 U441 ( .Y(n386), .A(n396) );
  nor02 U442 ( .Y(n397), .A0(n387), .A1(n388) );
  inv01 U443 ( .Y(n390), .A(n397) );
  inv02 U444 ( .Y(B_not[9]), .A(B[9]) );
  inv01 U445 ( .Y(DIFF[8]), .A(n398) );
  inv02 U446 ( .Y(carry_9_), .A(n399) );
  inv02 U447 ( .Y(n400), .A(B_not[8]) );
  inv02 U448 ( .Y(n401), .A(A[8]) );
  inv02 U449 ( .Y(n402), .A(carry_8_) );
  nor02 U450 ( .Y(n403), .A0(n400), .A1(n404) );
  nor02 U451 ( .Y(n405), .A0(n401), .A1(n406) );
  nor02 U452 ( .Y(n407), .A0(n402), .A1(n408) );
  nor02 U453 ( .Y(n409), .A0(n402), .A1(n410) );
  nor02 U454 ( .Y(n398), .A0(n411), .A1(n412) );
  nor02 U455 ( .Y(n413), .A0(n401), .A1(n402) );
  nor02 U456 ( .Y(n414), .A0(n400), .A1(n402) );
  nor02 U457 ( .Y(n415), .A0(n400), .A1(n401) );
  nor02 U458 ( .Y(n399), .A0(n415), .A1(n416) );
  nor02 U459 ( .Y(n417), .A0(A[8]), .A1(carry_8_) );
  inv01 U460 ( .Y(n404), .A(n417) );
  nor02 U461 ( .Y(n418), .A0(B_not[8]), .A1(carry_8_) );
  inv01 U462 ( .Y(n406), .A(n418) );
  nor02 U463 ( .Y(n419), .A0(B_not[8]), .A1(A[8]) );
  inv01 U464 ( .Y(n408), .A(n419) );
  nor02 U465 ( .Y(n420), .A0(n400), .A1(n401) );
  inv01 U466 ( .Y(n410), .A(n420) );
  nor02 U467 ( .Y(n421), .A0(n403), .A1(n405) );
  inv01 U468 ( .Y(n411), .A(n421) );
  nor02 U469 ( .Y(n422), .A0(n407), .A1(n409) );
  inv01 U470 ( .Y(n412), .A(n422) );
  nor02 U471 ( .Y(n423), .A0(n413), .A1(n414) );
  inv01 U472 ( .Y(n416), .A(n423) );
  inv02 U473 ( .Y(B_not[8]), .A(B[8]) );
  inv01 U474 ( .Y(DIFF[7]), .A(n424) );
  inv02 U475 ( .Y(carry_8_), .A(n425) );
  inv02 U476 ( .Y(n426), .A(B_not[7]) );
  inv02 U477 ( .Y(n427), .A(A[7]) );
  inv02 U478 ( .Y(n428), .A(carry_7_) );
  nor02 U479 ( .Y(n429), .A0(n426), .A1(n430) );
  nor02 U480 ( .Y(n431), .A0(n427), .A1(n432) );
  nor02 U481 ( .Y(n433), .A0(n428), .A1(n434) );
  nor02 U482 ( .Y(n435), .A0(n428), .A1(n436) );
  nor02 U483 ( .Y(n424), .A0(n437), .A1(n438) );
  nor02 U484 ( .Y(n439), .A0(n427), .A1(n428) );
  nor02 U485 ( .Y(n440), .A0(n426), .A1(n428) );
  nor02 U486 ( .Y(n441), .A0(n426), .A1(n427) );
  nor02 U487 ( .Y(n425), .A0(n441), .A1(n442) );
  nor02 U488 ( .Y(n443), .A0(A[7]), .A1(carry_7_) );
  inv01 U489 ( .Y(n430), .A(n443) );
  nor02 U490 ( .Y(n444), .A0(B_not[7]), .A1(carry_7_) );
  inv01 U491 ( .Y(n432), .A(n444) );
  nor02 U492 ( .Y(n445), .A0(B_not[7]), .A1(A[7]) );
  inv01 U493 ( .Y(n434), .A(n445) );
  nor02 U494 ( .Y(n446), .A0(n426), .A1(n427) );
  inv01 U495 ( .Y(n436), .A(n446) );
  nor02 U496 ( .Y(n447), .A0(n429), .A1(n431) );
  inv01 U497 ( .Y(n437), .A(n447) );
  nor02 U498 ( .Y(n448), .A0(n433), .A1(n435) );
  inv01 U499 ( .Y(n438), .A(n448) );
  nor02 U500 ( .Y(n449), .A0(n439), .A1(n440) );
  inv01 U501 ( .Y(n442), .A(n449) );
  inv02 U502 ( .Y(B_not[7]), .A(B[7]) );
  inv01 U503 ( .Y(DIFF[6]), .A(n450) );
  inv02 U504 ( .Y(carry_7_), .A(n451) );
  inv02 U505 ( .Y(n452), .A(B_not[6]) );
  inv02 U506 ( .Y(n453), .A(A[6]) );
  inv02 U507 ( .Y(n454), .A(carry_6_) );
  nor02 U508 ( .Y(n455), .A0(n452), .A1(n456) );
  nor02 U509 ( .Y(n457), .A0(n453), .A1(n458) );
  nor02 U510 ( .Y(n459), .A0(n454), .A1(n460) );
  nor02 U511 ( .Y(n461), .A0(n454), .A1(n462) );
  nor02 U512 ( .Y(n450), .A0(n463), .A1(n464) );
  nor02 U513 ( .Y(n465), .A0(n453), .A1(n454) );
  nor02 U514 ( .Y(n466), .A0(n452), .A1(n454) );
  nor02 U515 ( .Y(n467), .A0(n452), .A1(n453) );
  nor02 U516 ( .Y(n451), .A0(n467), .A1(n468) );
  nor02 U517 ( .Y(n469), .A0(A[6]), .A1(carry_6_) );
  inv01 U518 ( .Y(n456), .A(n469) );
  nor02 U519 ( .Y(n470), .A0(B_not[6]), .A1(carry_6_) );
  inv01 U520 ( .Y(n458), .A(n470) );
  nor02 U521 ( .Y(n471), .A0(B_not[6]), .A1(A[6]) );
  inv01 U522 ( .Y(n460), .A(n471) );
  nor02 U523 ( .Y(n472), .A0(n452), .A1(n453) );
  inv01 U524 ( .Y(n462), .A(n472) );
  nor02 U525 ( .Y(n473), .A0(n455), .A1(n457) );
  inv01 U526 ( .Y(n463), .A(n473) );
  nor02 U527 ( .Y(n474), .A0(n459), .A1(n461) );
  inv01 U528 ( .Y(n464), .A(n474) );
  nor02 U529 ( .Y(n475), .A0(n465), .A1(n466) );
  inv01 U530 ( .Y(n468), .A(n475) );
  inv02 U531 ( .Y(B_not[6]), .A(B[6]) );
  inv01 U532 ( .Y(DIFF[5]), .A(n476) );
  inv02 U533 ( .Y(carry_6_), .A(n477) );
  inv02 U534 ( .Y(n478), .A(B_not[5]) );
  inv02 U535 ( .Y(n479), .A(A[5]) );
  inv02 U536 ( .Y(n480), .A(carry_5_) );
  nor02 U537 ( .Y(n481), .A0(n478), .A1(n482) );
  nor02 U538 ( .Y(n483), .A0(n479), .A1(n484) );
  nor02 U539 ( .Y(n485), .A0(n480), .A1(n486) );
  nor02 U540 ( .Y(n487), .A0(n480), .A1(n488) );
  nor02 U541 ( .Y(n476), .A0(n489), .A1(n490) );
  nor02 U542 ( .Y(n491), .A0(n479), .A1(n480) );
  nor02 U543 ( .Y(n492), .A0(n478), .A1(n480) );
  nor02 U544 ( .Y(n493), .A0(n478), .A1(n479) );
  nor02 U545 ( .Y(n477), .A0(n493), .A1(n494) );
  nor02 U546 ( .Y(n495), .A0(A[5]), .A1(carry_5_) );
  inv01 U547 ( .Y(n482), .A(n495) );
  nor02 U548 ( .Y(n496), .A0(B_not[5]), .A1(carry_5_) );
  inv01 U549 ( .Y(n484), .A(n496) );
  nor02 U550 ( .Y(n497), .A0(B_not[5]), .A1(A[5]) );
  inv01 U551 ( .Y(n486), .A(n497) );
  nor02 U552 ( .Y(n498), .A0(n478), .A1(n479) );
  inv01 U553 ( .Y(n488), .A(n498) );
  nor02 U554 ( .Y(n499), .A0(n481), .A1(n483) );
  inv01 U555 ( .Y(n489), .A(n499) );
  nor02 U556 ( .Y(n500), .A0(n485), .A1(n487) );
  inv01 U557 ( .Y(n490), .A(n500) );
  nor02 U558 ( .Y(n501), .A0(n491), .A1(n492) );
  inv01 U559 ( .Y(n494), .A(n501) );
  inv02 U560 ( .Y(B_not[5]), .A(B[5]) );
  inv01 U561 ( .Y(DIFF[4]), .A(n502) );
  inv02 U562 ( .Y(carry_5_), .A(n503) );
  inv02 U563 ( .Y(n504), .A(B_not[4]) );
  inv02 U564 ( .Y(n505), .A(A[4]) );
  inv02 U565 ( .Y(n506), .A(carry_4_) );
  nor02 U566 ( .Y(n507), .A0(n504), .A1(n508) );
  nor02 U567 ( .Y(n509), .A0(n505), .A1(n510) );
  nor02 U568 ( .Y(n511), .A0(n506), .A1(n512) );
  nor02 U569 ( .Y(n513), .A0(n506), .A1(n514) );
  nor02 U570 ( .Y(n502), .A0(n515), .A1(n516) );
  nor02 U571 ( .Y(n517), .A0(n505), .A1(n506) );
  nor02 U572 ( .Y(n518), .A0(n504), .A1(n506) );
  nor02 U573 ( .Y(n519), .A0(n504), .A1(n505) );
  nor02 U574 ( .Y(n503), .A0(n519), .A1(n520) );
  nor02 U575 ( .Y(n521), .A0(A[4]), .A1(carry_4_) );
  inv01 U576 ( .Y(n508), .A(n521) );
  nor02 U577 ( .Y(n522), .A0(B_not[4]), .A1(carry_4_) );
  inv01 U578 ( .Y(n510), .A(n522) );
  nor02 U579 ( .Y(n523), .A0(B_not[4]), .A1(A[4]) );
  inv01 U580 ( .Y(n512), .A(n523) );
  nor02 U581 ( .Y(n524), .A0(n504), .A1(n505) );
  inv01 U582 ( .Y(n514), .A(n524) );
  nor02 U583 ( .Y(n525), .A0(n507), .A1(n509) );
  inv01 U584 ( .Y(n515), .A(n525) );
  nor02 U585 ( .Y(n526), .A0(n511), .A1(n513) );
  inv01 U586 ( .Y(n516), .A(n526) );
  nor02 U587 ( .Y(n527), .A0(n517), .A1(n518) );
  inv01 U588 ( .Y(n520), .A(n527) );
  inv02 U589 ( .Y(B_not[4]), .A(B[4]) );
  inv01 U590 ( .Y(DIFF[3]), .A(n528) );
  inv02 U591 ( .Y(carry_4_), .A(n529) );
  inv02 U592 ( .Y(n530), .A(B_not[3]) );
  inv02 U593 ( .Y(n531), .A(A[3]) );
  inv02 U594 ( .Y(n532), .A(carry_3_) );
  nor02 U595 ( .Y(n533), .A0(n530), .A1(n534) );
  nor02 U596 ( .Y(n535), .A0(n531), .A1(n536) );
  nor02 U597 ( .Y(n537), .A0(n532), .A1(n538) );
  nor02 U598 ( .Y(n539), .A0(n532), .A1(n540) );
  nor02 U599 ( .Y(n528), .A0(n541), .A1(n542) );
  nor02 U600 ( .Y(n543), .A0(n531), .A1(n532) );
  nor02 U601 ( .Y(n544), .A0(n530), .A1(n532) );
  nor02 U602 ( .Y(n545), .A0(n530), .A1(n531) );
  nor02 U603 ( .Y(n529), .A0(n545), .A1(n546) );
  nor02 U604 ( .Y(n547), .A0(A[3]), .A1(carry_3_) );
  inv01 U605 ( .Y(n534), .A(n547) );
  nor02 U606 ( .Y(n548), .A0(B_not[3]), .A1(carry_3_) );
  inv01 U607 ( .Y(n536), .A(n548) );
  nor02 U608 ( .Y(n549), .A0(B_not[3]), .A1(A[3]) );
  inv01 U609 ( .Y(n538), .A(n549) );
  nor02 U610 ( .Y(n550), .A0(n530), .A1(n531) );
  inv01 U611 ( .Y(n540), .A(n550) );
  nor02 U612 ( .Y(n551), .A0(n533), .A1(n535) );
  inv01 U613 ( .Y(n541), .A(n551) );
  nor02 U614 ( .Y(n552), .A0(n537), .A1(n539) );
  inv01 U615 ( .Y(n542), .A(n552) );
  nor02 U616 ( .Y(n553), .A0(n543), .A1(n544) );
  inv01 U617 ( .Y(n546), .A(n553) );
  inv02 U618 ( .Y(B_not[3]), .A(B[3]) );
  inv01 U619 ( .Y(DIFF[2]), .A(n554) );
  inv02 U620 ( .Y(carry_3_), .A(n555) );
  inv02 U621 ( .Y(n556), .A(B_not[2]) );
  inv02 U622 ( .Y(n557), .A(A[2]) );
  inv02 U623 ( .Y(n558), .A(n580) );
  nor02 U624 ( .Y(n559), .A0(n556), .A1(n560) );
  nor02 U625 ( .Y(n561), .A0(n557), .A1(n562) );
  nor02 U626 ( .Y(n563), .A0(n558), .A1(n564) );
  nor02 U627 ( .Y(n565), .A0(n558), .A1(n566) );
  nor02 U628 ( .Y(n554), .A0(n567), .A1(n568) );
  nor02 U629 ( .Y(n569), .A0(n557), .A1(n558) );
  nor02 U630 ( .Y(n570), .A0(n556), .A1(n558) );
  nor02 U631 ( .Y(n571), .A0(n556), .A1(n557) );
  nor02 U632 ( .Y(n555), .A0(n571), .A1(n572) );
  nor02 U633 ( .Y(n573), .A0(A[2]), .A1(n580) );
  inv01 U634 ( .Y(n560), .A(n573) );
  nor02 U635 ( .Y(n574), .A0(B_not[2]), .A1(n580) );
  inv01 U636 ( .Y(n562), .A(n574) );
  nor02 U637 ( .Y(n575), .A0(B_not[2]), .A1(A[2]) );
  inv01 U638 ( .Y(n564), .A(n575) );
  nor02 U639 ( .Y(n576), .A0(n556), .A1(n557) );
  inv01 U640 ( .Y(n566), .A(n576) );
  nor02 U641 ( .Y(n577), .A0(n559), .A1(n561) );
  inv01 U642 ( .Y(n567), .A(n577) );
  nor02 U643 ( .Y(n578), .A0(n563), .A1(n565) );
  inv01 U644 ( .Y(n568), .A(n578) );
  nor02 U645 ( .Y(n579), .A0(n569), .A1(n570) );
  inv01 U646 ( .Y(n572), .A(n579) );
  inv02 U647 ( .Y(B_not[2]), .A(B[2]) );
  buf02 U648 ( .Y(n580), .A(carry_2_) );
  xnor2 U649 ( .Y(DIFF[0]), .A0(B_not[0]), .A1(A[0]) );
  inv04 U650 ( .Y(B_not[24]), .A(B[24]) );
  inv04 U651 ( .Y(B_not[1]), .A(B[1]) );
  inv04 U652 ( .Y(B_not[0]), .A(B[0]) );
  fadd1 U2_1 ( .S(DIFF[1]), .CO(carry_2_), .A(A[1]), .B(B_not[1]), .CI(n6) );
  fadd1 U2_24 ( .S(DIFF[24]), .CO(carry_25_), .A(A[24]), .B(B_not[24]), .CI(
        carry_24_) );
  fadd1 U2_25 ( .S(DIFF[25]), .A(A[25]), .B(B_not[25]), .CI(n7) );
endmodule


module sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_add_52_0 ( A, B, CI, SUM, CO );
  input [51:0] A;
  input [51:0] B;
  output [51:0] SUM;
  input CI;
  output CO;
  wire   carry_51_, carry_50_, carry_49_, carry_48_, carry_47_, carry_46_,
         carry_45_, carry_44_, carry_43_, carry_42_, carry_41_, carry_40_,
         carry_39_, carry_38_, carry_37_, carry_36_, carry_35_, carry_34_,
         carry_33_, carry_32_, carry_31_, carry_30_, carry_29_, carry_28_,
         carry_27_, carry_26_, carry_25_, carry_24_, carry_23_, carry_22_,
         carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, carry_6_, carry_5_, carry_4_, carry_3_,
         carry_2_, n1325, n1, n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324;

  or02 U4 ( .Y(n1), .A0(n329), .A1(n330) );
  inv02 U5 ( .Y(n2), .A(n1) );
  nand02 U6 ( .Y(n3), .A0(A[0]), .A1(B[0]) );
  inv02 U7 ( .Y(n4), .A(n3) );
  inv02 U8 ( .Y(SUM[50]), .A(n292) );
  inv02 U9 ( .Y(SUM[49]), .A(n441) );
  inv02 U10 ( .Y(SUM[48]), .A(n363) );
  inv02 U11 ( .Y(SUM[47]), .A(n545) );
  inv02 U12 ( .Y(SUM[46]), .A(n467) );
  inv02 U13 ( .Y(SUM[45]), .A(n623) );
  inv02 U14 ( .Y(SUM[44]), .A(n58) );
  inv02 U15 ( .Y(SUM[43]), .A(n240) );
  inv02 U16 ( .Y(SUM[22]), .A(n805) );
  inv02 U17 ( .Y(SUM[42]), .A(n214) );
  inv02 U18 ( .Y(SUM[23]), .A(n831) );
  inv02 U19 ( .Y(SUM[41]), .A(n6) );
  inv02 U20 ( .Y(SUM[21]), .A(n961) );
  inv02 U21 ( .Y(SUM[24]), .A(n701) );
  inv02 U22 ( .Y(SUM[40]), .A(n136) );
  inv02 U23 ( .Y(SUM[20]), .A(n909) );
  inv02 U24 ( .Y(SUM[25]), .A(n727) );
  inv02 U25 ( .Y(SUM[19]), .A(n987) );
  inv02 U26 ( .Y(SUM[39]), .A(n32) );
  inv02 U27 ( .Y(SUM[26]), .A(n571) );
  inv02 U28 ( .Y(SUM[18]), .A(n1143) );
  inv02 U29 ( .Y(SUM[38]), .A(n110) );
  inv02 U30 ( .Y(SUM[27]), .A(n597) );
  inv02 U31 ( .Y(SUM[37]), .A(n84) );
  inv02 U32 ( .Y(SUM[17]), .A(n1273) );
  inv02 U33 ( .Y(SUM[28]), .A(n493) );
  inv02 U34 ( .Y(SUM[36]), .A(n188) );
  inv02 U35 ( .Y(SUM[16]), .A(n1065) );
  inv02 U36 ( .Y(SUM[29]), .A(n649) );
  inv02 U37 ( .Y(SUM[35]), .A(n162) );
  inv02 U38 ( .Y(SUM[15]), .A(n1039) );
  inv02 U39 ( .Y(SUM[30]), .A(n519) );
  inv02 U40 ( .Y(SUM[14]), .A(n1169) );
  inv02 U41 ( .Y(SUM[34]), .A(n337) );
  inv02 U42 ( .Y(SUM[31]), .A(n389) );
  inv02 U43 ( .Y(SUM[33]), .A(n266) );
  inv02 U44 ( .Y(SUM[13]), .A(n1117) );
  inv02 U45 ( .Y(SUM[32]), .A(n415) );
  inv02 U46 ( .Y(SUM[12]), .A(n1247) );
  inv02 U47 ( .Y(SUM[11]), .A(n753) );
  inv02 U48 ( .Y(SUM[10]), .A(n675) );
  inv02 U49 ( .Y(SUM[9]), .A(n857) );
  inv02 U50 ( .Y(SUM[8]), .A(n779) );
  inv02 U51 ( .Y(SUM[7]), .A(n935) );
  inv02 U52 ( .Y(SUM[6]), .A(n883) );
  inv02 U53 ( .Y(SUM[5]), .A(n1013) );
  inv02 U54 ( .Y(SUM[4]), .A(n1091) );
  inv02 U55 ( .Y(SUM[3]), .A(n1221) );
  inv02 U56 ( .Y(SUM[2]), .A(n1195) );
  inv02 U57 ( .Y(SUM[1]), .A(n1299) );
  buf02 U58 ( .Y(SUM[0]), .A(n1325) );
  inv02 U59 ( .Y(carry_42_), .A(n7) );
  inv02 U60 ( .Y(n8), .A(B[41]) );
  inv02 U61 ( .Y(n9), .A(A[41]) );
  inv04 U62 ( .Y(n10), .A(carry_41_) );
  nor02 U63 ( .Y(n11), .A0(n8), .A1(n12) );
  nor02 U64 ( .Y(n13), .A0(n9), .A1(n14) );
  nor02 U65 ( .Y(n15), .A0(n10), .A1(n16) );
  nor02 U66 ( .Y(n17), .A0(n10), .A1(n18) );
  nor02 U67 ( .Y(n6), .A0(n19), .A1(n20) );
  nor02 U68 ( .Y(n21), .A0(n9), .A1(n10) );
  nor02 U69 ( .Y(n22), .A0(n8), .A1(n10) );
  nor02 U70 ( .Y(n23), .A0(n8), .A1(n9) );
  nor02 U71 ( .Y(n7), .A0(n23), .A1(n24) );
  nor02 U72 ( .Y(n25), .A0(A[41]), .A1(carry_41_) );
  inv01 U73 ( .Y(n12), .A(n25) );
  nor02 U74 ( .Y(n26), .A0(B[41]), .A1(carry_41_) );
  inv01 U75 ( .Y(n14), .A(n26) );
  nor02 U76 ( .Y(n27), .A0(B[41]), .A1(A[41]) );
  inv01 U77 ( .Y(n16), .A(n27) );
  nor02 U78 ( .Y(n28), .A0(n8), .A1(n9) );
  inv01 U79 ( .Y(n18), .A(n28) );
  nor02 U80 ( .Y(n29), .A0(n11), .A1(n13) );
  inv02 U81 ( .Y(n19), .A(n29) );
  nor02 U82 ( .Y(n30), .A0(n15), .A1(n17) );
  inv02 U83 ( .Y(n20), .A(n30) );
  nor02 U84 ( .Y(n31), .A0(n21), .A1(n22) );
  inv01 U85 ( .Y(n24), .A(n31) );
  inv02 U86 ( .Y(carry_40_), .A(n33) );
  inv02 U87 ( .Y(n34), .A(B[39]) );
  inv02 U88 ( .Y(n35), .A(A[39]) );
  inv04 U89 ( .Y(n36), .A(carry_39_) );
  nor02 U90 ( .Y(n37), .A0(n34), .A1(n38) );
  nor02 U91 ( .Y(n39), .A0(n35), .A1(n40) );
  nor02 U92 ( .Y(n41), .A0(n36), .A1(n42) );
  nor02 U93 ( .Y(n43), .A0(n36), .A1(n44) );
  nor02 U94 ( .Y(n32), .A0(n45), .A1(n46) );
  nor02 U95 ( .Y(n47), .A0(n35), .A1(n36) );
  nor02 U96 ( .Y(n48), .A0(n34), .A1(n36) );
  nor02 U97 ( .Y(n49), .A0(n34), .A1(n35) );
  nor02 U98 ( .Y(n33), .A0(n49), .A1(n50) );
  nor02 U99 ( .Y(n51), .A0(A[39]), .A1(carry_39_) );
  inv01 U100 ( .Y(n38), .A(n51) );
  nor02 U101 ( .Y(n52), .A0(B[39]), .A1(carry_39_) );
  inv01 U102 ( .Y(n40), .A(n52) );
  nor02 U103 ( .Y(n53), .A0(B[39]), .A1(A[39]) );
  inv01 U104 ( .Y(n42), .A(n53) );
  nor02 U105 ( .Y(n54), .A0(n34), .A1(n35) );
  inv01 U106 ( .Y(n44), .A(n54) );
  nor02 U107 ( .Y(n55), .A0(n37), .A1(n39) );
  inv02 U108 ( .Y(n45), .A(n55) );
  nor02 U109 ( .Y(n56), .A0(n41), .A1(n43) );
  inv02 U110 ( .Y(n46), .A(n56) );
  nor02 U111 ( .Y(n57), .A0(n47), .A1(n48) );
  inv01 U112 ( .Y(n50), .A(n57) );
  inv02 U113 ( .Y(carry_45_), .A(n59) );
  inv02 U114 ( .Y(n60), .A(B[44]) );
  inv02 U115 ( .Y(n61), .A(A[44]) );
  inv04 U116 ( .Y(n62), .A(carry_44_) );
  nor02 U117 ( .Y(n63), .A0(n60), .A1(n64) );
  nor02 U118 ( .Y(n65), .A0(n61), .A1(n66) );
  nor02 U119 ( .Y(n67), .A0(n62), .A1(n68) );
  nor02 U120 ( .Y(n69), .A0(n62), .A1(n70) );
  nor02 U121 ( .Y(n58), .A0(n71), .A1(n72) );
  nor02 U122 ( .Y(n73), .A0(n61), .A1(n62) );
  nor02 U123 ( .Y(n74), .A0(n60), .A1(n62) );
  nor02 U124 ( .Y(n75), .A0(n60), .A1(n61) );
  nor02 U125 ( .Y(n59), .A0(n75), .A1(n76) );
  nor02 U126 ( .Y(n77), .A0(A[44]), .A1(carry_44_) );
  inv01 U127 ( .Y(n64), .A(n77) );
  nor02 U128 ( .Y(n78), .A0(B[44]), .A1(carry_44_) );
  inv01 U129 ( .Y(n66), .A(n78) );
  nor02 U130 ( .Y(n79), .A0(B[44]), .A1(A[44]) );
  inv01 U131 ( .Y(n68), .A(n79) );
  nor02 U132 ( .Y(n80), .A0(n60), .A1(n61) );
  inv01 U133 ( .Y(n70), .A(n80) );
  nor02 U134 ( .Y(n81), .A0(n63), .A1(n65) );
  inv02 U135 ( .Y(n71), .A(n81) );
  nor02 U136 ( .Y(n82), .A0(n67), .A1(n69) );
  inv02 U137 ( .Y(n72), .A(n82) );
  nor02 U138 ( .Y(n83), .A0(n73), .A1(n74) );
  inv01 U139 ( .Y(n76), .A(n83) );
  inv02 U140 ( .Y(carry_38_), .A(n85) );
  inv02 U141 ( .Y(n86), .A(B[37]) );
  inv02 U142 ( .Y(n87), .A(A[37]) );
  inv04 U143 ( .Y(n88), .A(carry_37_) );
  nor02 U144 ( .Y(n89), .A0(n86), .A1(n90) );
  nor02 U145 ( .Y(n91), .A0(n87), .A1(n92) );
  nor02 U146 ( .Y(n93), .A0(n88), .A1(n94) );
  nor02 U147 ( .Y(n95), .A0(n88), .A1(n96) );
  nor02 U148 ( .Y(n84), .A0(n97), .A1(n98) );
  nor02 U149 ( .Y(n99), .A0(n87), .A1(n88) );
  nor02 U150 ( .Y(n100), .A0(n86), .A1(n88) );
  nor02 U151 ( .Y(n101), .A0(n86), .A1(n87) );
  nor02 U152 ( .Y(n85), .A0(n101), .A1(n102) );
  nor02 U153 ( .Y(n103), .A0(A[37]), .A1(carry_37_) );
  inv01 U154 ( .Y(n90), .A(n103) );
  nor02 U155 ( .Y(n104), .A0(B[37]), .A1(carry_37_) );
  inv01 U156 ( .Y(n92), .A(n104) );
  nor02 U157 ( .Y(n105), .A0(B[37]), .A1(A[37]) );
  inv01 U158 ( .Y(n94), .A(n105) );
  nor02 U159 ( .Y(n106), .A0(n86), .A1(n87) );
  inv01 U160 ( .Y(n96), .A(n106) );
  nor02 U161 ( .Y(n107), .A0(n89), .A1(n91) );
  inv02 U162 ( .Y(n97), .A(n107) );
  nor02 U163 ( .Y(n108), .A0(n93), .A1(n95) );
  inv02 U164 ( .Y(n98), .A(n108) );
  nor02 U165 ( .Y(n109), .A0(n99), .A1(n100) );
  inv01 U166 ( .Y(n102), .A(n109) );
  inv02 U167 ( .Y(carry_39_), .A(n111) );
  inv02 U168 ( .Y(n112), .A(B[38]) );
  inv02 U169 ( .Y(n113), .A(A[38]) );
  inv04 U170 ( .Y(n114), .A(carry_38_) );
  nor02 U171 ( .Y(n115), .A0(n112), .A1(n116) );
  nor02 U172 ( .Y(n117), .A0(n113), .A1(n118) );
  nor02 U173 ( .Y(n119), .A0(n114), .A1(n120) );
  nor02 U174 ( .Y(n121), .A0(n114), .A1(n122) );
  nor02 U175 ( .Y(n110), .A0(n123), .A1(n124) );
  nor02 U176 ( .Y(n125), .A0(n113), .A1(n114) );
  nor02 U177 ( .Y(n126), .A0(n112), .A1(n114) );
  nor02 U178 ( .Y(n127), .A0(n112), .A1(n113) );
  nor02 U179 ( .Y(n111), .A0(n127), .A1(n128) );
  nor02 U180 ( .Y(n129), .A0(A[38]), .A1(carry_38_) );
  inv01 U181 ( .Y(n116), .A(n129) );
  nor02 U182 ( .Y(n130), .A0(B[38]), .A1(carry_38_) );
  inv01 U183 ( .Y(n118), .A(n130) );
  nor02 U184 ( .Y(n131), .A0(B[38]), .A1(A[38]) );
  inv01 U185 ( .Y(n120), .A(n131) );
  nor02 U186 ( .Y(n132), .A0(n112), .A1(n113) );
  inv01 U187 ( .Y(n122), .A(n132) );
  nor02 U188 ( .Y(n133), .A0(n115), .A1(n117) );
  inv02 U189 ( .Y(n123), .A(n133) );
  nor02 U190 ( .Y(n134), .A0(n119), .A1(n121) );
  inv02 U191 ( .Y(n124), .A(n134) );
  nor02 U192 ( .Y(n135), .A0(n125), .A1(n126) );
  inv01 U193 ( .Y(n128), .A(n135) );
  inv02 U194 ( .Y(carry_41_), .A(n137) );
  inv02 U195 ( .Y(n138), .A(B[40]) );
  inv02 U196 ( .Y(n139), .A(A[40]) );
  inv02 U197 ( .Y(n140), .A(carry_40_) );
  nor02 U198 ( .Y(n141), .A0(n138), .A1(n142) );
  nor02 U199 ( .Y(n143), .A0(n139), .A1(n144) );
  nor02 U200 ( .Y(n145), .A0(n140), .A1(n146) );
  nor02 U201 ( .Y(n147), .A0(n140), .A1(n148) );
  nor02 U202 ( .Y(n136), .A0(n149), .A1(n150) );
  nor02 U203 ( .Y(n151), .A0(n139), .A1(n140) );
  nor02 U204 ( .Y(n152), .A0(n138), .A1(n140) );
  nor02 U205 ( .Y(n153), .A0(n138), .A1(n139) );
  nor02 U206 ( .Y(n137), .A0(n153), .A1(n154) );
  nor02 U207 ( .Y(n155), .A0(A[40]), .A1(carry_40_) );
  inv01 U208 ( .Y(n142), .A(n155) );
  nor02 U209 ( .Y(n156), .A0(B[40]), .A1(carry_40_) );
  inv01 U210 ( .Y(n144), .A(n156) );
  nor02 U211 ( .Y(n157), .A0(B[40]), .A1(A[40]) );
  inv01 U212 ( .Y(n146), .A(n157) );
  nor02 U213 ( .Y(n158), .A0(n138), .A1(n139) );
  inv01 U214 ( .Y(n148), .A(n158) );
  nor02 U215 ( .Y(n159), .A0(n141), .A1(n143) );
  inv02 U216 ( .Y(n149), .A(n159) );
  nor02 U217 ( .Y(n160), .A0(n145), .A1(n147) );
  inv02 U218 ( .Y(n150), .A(n160) );
  nor02 U219 ( .Y(n161), .A0(n151), .A1(n152) );
  inv01 U220 ( .Y(n154), .A(n161) );
  inv02 U221 ( .Y(carry_36_), .A(n163) );
  inv02 U222 ( .Y(n164), .A(B[35]) );
  inv02 U223 ( .Y(n165), .A(A[35]) );
  inv04 U224 ( .Y(n166), .A(carry_35_) );
  nor02 U225 ( .Y(n167), .A0(n164), .A1(n168) );
  nor02 U226 ( .Y(n169), .A0(n165), .A1(n170) );
  nor02 U227 ( .Y(n171), .A0(n166), .A1(n172) );
  nor02 U228 ( .Y(n173), .A0(n166), .A1(n174) );
  nor02 U229 ( .Y(n162), .A0(n175), .A1(n176) );
  nor02 U230 ( .Y(n177), .A0(n165), .A1(n166) );
  nor02 U231 ( .Y(n178), .A0(n164), .A1(n166) );
  nor02 U232 ( .Y(n179), .A0(n164), .A1(n165) );
  nor02 U233 ( .Y(n163), .A0(n179), .A1(n180) );
  nor02 U234 ( .Y(n181), .A0(A[35]), .A1(carry_35_) );
  inv01 U235 ( .Y(n168), .A(n181) );
  nor02 U236 ( .Y(n182), .A0(B[35]), .A1(carry_35_) );
  inv01 U237 ( .Y(n170), .A(n182) );
  nor02 U238 ( .Y(n183), .A0(B[35]), .A1(A[35]) );
  inv01 U239 ( .Y(n172), .A(n183) );
  nor02 U240 ( .Y(n184), .A0(n164), .A1(n165) );
  inv01 U241 ( .Y(n174), .A(n184) );
  nor02 U242 ( .Y(n185), .A0(n167), .A1(n169) );
  inv02 U243 ( .Y(n175), .A(n185) );
  nor02 U244 ( .Y(n186), .A0(n171), .A1(n173) );
  inv02 U245 ( .Y(n176), .A(n186) );
  nor02 U246 ( .Y(n187), .A0(n177), .A1(n178) );
  inv01 U247 ( .Y(n180), .A(n187) );
  inv02 U248 ( .Y(carry_37_), .A(n189) );
  inv02 U249 ( .Y(n190), .A(B[36]) );
  inv02 U250 ( .Y(n191), .A(A[36]) );
  inv04 U251 ( .Y(n192), .A(carry_36_) );
  nor02 U252 ( .Y(n193), .A0(n190), .A1(n194) );
  nor02 U253 ( .Y(n195), .A0(n191), .A1(n196) );
  nor02 U254 ( .Y(n197), .A0(n192), .A1(n198) );
  nor02 U255 ( .Y(n199), .A0(n192), .A1(n200) );
  nor02 U256 ( .Y(n188), .A0(n201), .A1(n202) );
  nor02 U257 ( .Y(n203), .A0(n191), .A1(n192) );
  nor02 U258 ( .Y(n204), .A0(n190), .A1(n192) );
  nor02 U259 ( .Y(n205), .A0(n190), .A1(n191) );
  nor02 U260 ( .Y(n189), .A0(n205), .A1(n206) );
  nor02 U261 ( .Y(n207), .A0(A[36]), .A1(carry_36_) );
  inv01 U262 ( .Y(n194), .A(n207) );
  nor02 U263 ( .Y(n208), .A0(B[36]), .A1(carry_36_) );
  inv01 U264 ( .Y(n196), .A(n208) );
  nor02 U265 ( .Y(n209), .A0(B[36]), .A1(A[36]) );
  inv01 U266 ( .Y(n198), .A(n209) );
  nor02 U267 ( .Y(n210), .A0(n190), .A1(n191) );
  inv01 U268 ( .Y(n200), .A(n210) );
  nor02 U269 ( .Y(n211), .A0(n193), .A1(n195) );
  inv02 U270 ( .Y(n201), .A(n211) );
  nor02 U271 ( .Y(n212), .A0(n197), .A1(n199) );
  inv02 U272 ( .Y(n202), .A(n212) );
  nor02 U273 ( .Y(n213), .A0(n203), .A1(n204) );
  inv01 U274 ( .Y(n206), .A(n213) );
  inv02 U275 ( .Y(carry_43_), .A(n215) );
  inv02 U276 ( .Y(n216), .A(B[42]) );
  inv02 U277 ( .Y(n217), .A(A[42]) );
  inv02 U278 ( .Y(n218), .A(carry_42_) );
  nor02 U279 ( .Y(n219), .A0(n216), .A1(n220) );
  nor02 U280 ( .Y(n221), .A0(n217), .A1(n222) );
  nor02 U281 ( .Y(n223), .A0(n218), .A1(n224) );
  nor02 U282 ( .Y(n225), .A0(n218), .A1(n226) );
  nor02 U283 ( .Y(n214), .A0(n227), .A1(n228) );
  nor02 U284 ( .Y(n229), .A0(n217), .A1(n218) );
  nor02 U285 ( .Y(n230), .A0(n216), .A1(n218) );
  nor02 U286 ( .Y(n231), .A0(n216), .A1(n217) );
  nor02 U287 ( .Y(n215), .A0(n231), .A1(n232) );
  nor02 U288 ( .Y(n233), .A0(A[42]), .A1(carry_42_) );
  inv01 U289 ( .Y(n220), .A(n233) );
  nor02 U290 ( .Y(n234), .A0(B[42]), .A1(carry_42_) );
  inv01 U291 ( .Y(n222), .A(n234) );
  nor02 U292 ( .Y(n235), .A0(B[42]), .A1(A[42]) );
  inv01 U293 ( .Y(n224), .A(n235) );
  nor02 U294 ( .Y(n236), .A0(n216), .A1(n217) );
  inv01 U295 ( .Y(n226), .A(n236) );
  nor02 U296 ( .Y(n237), .A0(n219), .A1(n221) );
  inv02 U297 ( .Y(n227), .A(n237) );
  nor02 U298 ( .Y(n238), .A0(n223), .A1(n225) );
  inv02 U299 ( .Y(n228), .A(n238) );
  nor02 U300 ( .Y(n239), .A0(n229), .A1(n230) );
  inv01 U301 ( .Y(n232), .A(n239) );
  inv02 U302 ( .Y(carry_44_), .A(n241) );
  inv02 U303 ( .Y(n242), .A(B[43]) );
  inv02 U304 ( .Y(n243), .A(A[43]) );
  inv04 U305 ( .Y(n244), .A(carry_43_) );
  nor02 U306 ( .Y(n245), .A0(n242), .A1(n246) );
  nor02 U307 ( .Y(n247), .A0(n243), .A1(n248) );
  nor02 U308 ( .Y(n249), .A0(n244), .A1(n250) );
  nor02 U309 ( .Y(n251), .A0(n244), .A1(n252) );
  nor02 U310 ( .Y(n240), .A0(n253), .A1(n254) );
  nor02 U311 ( .Y(n255), .A0(n243), .A1(n244) );
  nor02 U312 ( .Y(n256), .A0(n242), .A1(n244) );
  nor02 U313 ( .Y(n257), .A0(n242), .A1(n243) );
  nor02 U314 ( .Y(n241), .A0(n257), .A1(n258) );
  nor02 U315 ( .Y(n259), .A0(A[43]), .A1(carry_43_) );
  inv01 U316 ( .Y(n246), .A(n259) );
  nor02 U317 ( .Y(n260), .A0(B[43]), .A1(carry_43_) );
  inv01 U318 ( .Y(n248), .A(n260) );
  nor02 U319 ( .Y(n261), .A0(B[43]), .A1(A[43]) );
  inv01 U320 ( .Y(n250), .A(n261) );
  nor02 U321 ( .Y(n262), .A0(n242), .A1(n243) );
  inv01 U322 ( .Y(n252), .A(n262) );
  nor02 U323 ( .Y(n263), .A0(n245), .A1(n247) );
  inv02 U324 ( .Y(n253), .A(n263) );
  nor02 U325 ( .Y(n264), .A0(n249), .A1(n251) );
  inv02 U326 ( .Y(n254), .A(n264) );
  nor02 U327 ( .Y(n265), .A0(n255), .A1(n256) );
  inv01 U328 ( .Y(n258), .A(n265) );
  inv02 U329 ( .Y(carry_34_), .A(n267) );
  inv02 U330 ( .Y(n268), .A(B[33]) );
  inv02 U331 ( .Y(n269), .A(A[33]) );
  inv04 U332 ( .Y(n270), .A(carry_33_) );
  nor02 U333 ( .Y(n271), .A0(n268), .A1(n272) );
  nor02 U334 ( .Y(n273), .A0(n269), .A1(n274) );
  nor02 U335 ( .Y(n275), .A0(n270), .A1(n276) );
  nor02 U336 ( .Y(n277), .A0(n270), .A1(n278) );
  nor02 U337 ( .Y(n266), .A0(n279), .A1(n280) );
  nor02 U338 ( .Y(n281), .A0(n269), .A1(n270) );
  nor02 U339 ( .Y(n282), .A0(n268), .A1(n270) );
  nor02 U340 ( .Y(n283), .A0(n268), .A1(n269) );
  nor02 U341 ( .Y(n267), .A0(n283), .A1(n284) );
  nor02 U342 ( .Y(n285), .A0(A[33]), .A1(carry_33_) );
  inv01 U343 ( .Y(n272), .A(n285) );
  nor02 U344 ( .Y(n286), .A0(B[33]), .A1(carry_33_) );
  inv01 U345 ( .Y(n274), .A(n286) );
  nor02 U346 ( .Y(n287), .A0(B[33]), .A1(A[33]) );
  inv01 U347 ( .Y(n276), .A(n287) );
  nor02 U348 ( .Y(n288), .A0(n268), .A1(n269) );
  inv01 U349 ( .Y(n278), .A(n288) );
  nor02 U350 ( .Y(n289), .A0(n271), .A1(n273) );
  inv02 U351 ( .Y(n279), .A(n289) );
  nor02 U352 ( .Y(n290), .A0(n275), .A1(n277) );
  inv02 U353 ( .Y(n280), .A(n290) );
  nor02 U354 ( .Y(n291), .A0(n281), .A1(n282) );
  inv01 U355 ( .Y(n284), .A(n291) );
  inv02 U356 ( .Y(carry_51_), .A(n293) );
  inv02 U357 ( .Y(n294), .A(B[50]) );
  inv02 U358 ( .Y(n295), .A(A[50]) );
  inv04 U359 ( .Y(n296), .A(carry_50_) );
  nor02 U360 ( .Y(n297), .A0(n294), .A1(n298) );
  nor02 U361 ( .Y(n299), .A0(n295), .A1(n300) );
  nor02 U362 ( .Y(n301), .A0(n296), .A1(n302) );
  nor02 U363 ( .Y(n303), .A0(n296), .A1(n304) );
  nor02 U364 ( .Y(n292), .A0(n305), .A1(n306) );
  nor02 U365 ( .Y(n307), .A0(n295), .A1(n296) );
  nor02 U366 ( .Y(n308), .A0(n294), .A1(n296) );
  nor02 U367 ( .Y(n309), .A0(n294), .A1(n295) );
  nor02 U368 ( .Y(n293), .A0(n309), .A1(n310) );
  nor02 U369 ( .Y(n311), .A0(A[50]), .A1(carry_50_) );
  inv01 U370 ( .Y(n298), .A(n311) );
  nor02 U371 ( .Y(n312), .A0(B[50]), .A1(carry_50_) );
  inv01 U372 ( .Y(n300), .A(n312) );
  nor02 U373 ( .Y(n313), .A0(B[50]), .A1(A[50]) );
  inv01 U374 ( .Y(n302), .A(n313) );
  nor02 U375 ( .Y(n314), .A0(n294), .A1(n295) );
  inv01 U376 ( .Y(n304), .A(n314) );
  nor02 U377 ( .Y(n315), .A0(n297), .A1(n299) );
  inv02 U378 ( .Y(n305), .A(n315) );
  nor02 U379 ( .Y(n316), .A0(n301), .A1(n303) );
  inv02 U380 ( .Y(n306), .A(n316) );
  nor02 U381 ( .Y(n317), .A0(n307), .A1(n308) );
  inv01 U382 ( .Y(n310), .A(n317) );
  inv04 U383 ( .Y(SUM[51]), .A(n2) );
  inv01 U384 ( .Y(n318), .A(B[51]) );
  inv01 U385 ( .Y(n319), .A(A[51]) );
  inv02 U386 ( .Y(n320), .A(carry_51_) );
  nor02 U387 ( .Y(n321), .A0(n318), .A1(n322) );
  nor02 U388 ( .Y(n323), .A0(n319), .A1(n324) );
  nor02 U389 ( .Y(n325), .A0(n320), .A1(n326) );
  nor02 U390 ( .Y(n327), .A0(n320), .A1(n328) );
  nor02 U391 ( .Y(n331), .A0(A[51]), .A1(carry_51_) );
  inv01 U392 ( .Y(n322), .A(n331) );
  nor02 U393 ( .Y(n332), .A0(B[51]), .A1(carry_51_) );
  inv01 U394 ( .Y(n324), .A(n332) );
  nor02 U395 ( .Y(n333), .A0(B[51]), .A1(A[51]) );
  inv01 U396 ( .Y(n326), .A(n333) );
  nor02 U397 ( .Y(n334), .A0(n318), .A1(n319) );
  inv01 U398 ( .Y(n328), .A(n334) );
  nor02 U399 ( .Y(n335), .A0(n321), .A1(n323) );
  inv02 U400 ( .Y(n329), .A(n335) );
  nor02 U401 ( .Y(n336), .A0(n325), .A1(n327) );
  inv02 U402 ( .Y(n330), .A(n336) );
  inv02 U403 ( .Y(carry_35_), .A(n338) );
  inv02 U404 ( .Y(n339), .A(B[34]) );
  inv02 U405 ( .Y(n340), .A(A[34]) );
  inv04 U406 ( .Y(n341), .A(carry_34_) );
  nor02 U407 ( .Y(n342), .A0(n339), .A1(n343) );
  nor02 U408 ( .Y(n344), .A0(n340), .A1(n345) );
  nor02 U409 ( .Y(n346), .A0(n341), .A1(n347) );
  nor02 U410 ( .Y(n348), .A0(n341), .A1(n349) );
  nor02 U411 ( .Y(n337), .A0(n350), .A1(n351) );
  nor02 U412 ( .Y(n352), .A0(n340), .A1(n341) );
  nor02 U413 ( .Y(n353), .A0(n339), .A1(n341) );
  nor02 U414 ( .Y(n354), .A0(n339), .A1(n340) );
  nor02 U415 ( .Y(n338), .A0(n354), .A1(n355) );
  nor02 U416 ( .Y(n356), .A0(A[34]), .A1(carry_34_) );
  inv01 U417 ( .Y(n343), .A(n356) );
  nor02 U418 ( .Y(n357), .A0(B[34]), .A1(carry_34_) );
  inv01 U419 ( .Y(n345), .A(n357) );
  nor02 U420 ( .Y(n358), .A0(B[34]), .A1(A[34]) );
  inv01 U421 ( .Y(n347), .A(n358) );
  nor02 U422 ( .Y(n359), .A0(n339), .A1(n340) );
  inv01 U423 ( .Y(n349), .A(n359) );
  nor02 U424 ( .Y(n360), .A0(n342), .A1(n344) );
  inv02 U425 ( .Y(n350), .A(n360) );
  nor02 U426 ( .Y(n361), .A0(n346), .A1(n348) );
  inv02 U427 ( .Y(n351), .A(n361) );
  nor02 U428 ( .Y(n362), .A0(n352), .A1(n353) );
  inv01 U429 ( .Y(n355), .A(n362) );
  inv02 U430 ( .Y(carry_49_), .A(n364) );
  inv02 U431 ( .Y(n365), .A(B[48]) );
  inv02 U432 ( .Y(n366), .A(A[48]) );
  inv04 U433 ( .Y(n367), .A(carry_48_) );
  nor02 U434 ( .Y(n368), .A0(n365), .A1(n369) );
  nor02 U435 ( .Y(n370), .A0(n366), .A1(n371) );
  nor02 U436 ( .Y(n372), .A0(n367), .A1(n373) );
  nor02 U437 ( .Y(n374), .A0(n367), .A1(n375) );
  nor02 U438 ( .Y(n363), .A0(n376), .A1(n377) );
  nor02 U439 ( .Y(n378), .A0(n366), .A1(n367) );
  nor02 U440 ( .Y(n379), .A0(n365), .A1(n367) );
  nor02 U441 ( .Y(n380), .A0(n365), .A1(n366) );
  nor02 U442 ( .Y(n364), .A0(n380), .A1(n381) );
  nor02 U443 ( .Y(n382), .A0(A[48]), .A1(carry_48_) );
  inv01 U444 ( .Y(n369), .A(n382) );
  nor02 U445 ( .Y(n383), .A0(B[48]), .A1(carry_48_) );
  inv01 U446 ( .Y(n371), .A(n383) );
  nor02 U447 ( .Y(n384), .A0(B[48]), .A1(A[48]) );
  inv01 U448 ( .Y(n373), .A(n384) );
  nor02 U449 ( .Y(n385), .A0(n365), .A1(n366) );
  inv01 U450 ( .Y(n375), .A(n385) );
  nor02 U451 ( .Y(n386), .A0(n368), .A1(n370) );
  inv02 U452 ( .Y(n376), .A(n386) );
  nor02 U453 ( .Y(n387), .A0(n372), .A1(n374) );
  inv02 U454 ( .Y(n377), .A(n387) );
  nor02 U455 ( .Y(n388), .A0(n378), .A1(n379) );
  inv01 U456 ( .Y(n381), .A(n388) );
  inv02 U457 ( .Y(carry_32_), .A(n390) );
  inv02 U458 ( .Y(n391), .A(B[31]) );
  inv02 U459 ( .Y(n392), .A(A[31]) );
  inv04 U460 ( .Y(n393), .A(carry_31_) );
  nor02 U461 ( .Y(n394), .A0(n391), .A1(n395) );
  nor02 U462 ( .Y(n396), .A0(n392), .A1(n397) );
  nor02 U463 ( .Y(n398), .A0(n393), .A1(n399) );
  nor02 U464 ( .Y(n400), .A0(n393), .A1(n401) );
  nor02 U465 ( .Y(n389), .A0(n402), .A1(n403) );
  nor02 U466 ( .Y(n404), .A0(n392), .A1(n393) );
  nor02 U467 ( .Y(n405), .A0(n391), .A1(n393) );
  nor02 U468 ( .Y(n406), .A0(n391), .A1(n392) );
  nor02 U469 ( .Y(n390), .A0(n406), .A1(n407) );
  nor02 U470 ( .Y(n408), .A0(A[31]), .A1(carry_31_) );
  inv01 U471 ( .Y(n395), .A(n408) );
  nor02 U472 ( .Y(n409), .A0(B[31]), .A1(carry_31_) );
  inv01 U473 ( .Y(n397), .A(n409) );
  nor02 U474 ( .Y(n410), .A0(B[31]), .A1(A[31]) );
  inv01 U475 ( .Y(n399), .A(n410) );
  nor02 U476 ( .Y(n411), .A0(n391), .A1(n392) );
  inv01 U477 ( .Y(n401), .A(n411) );
  nor02 U478 ( .Y(n412), .A0(n394), .A1(n396) );
  inv02 U479 ( .Y(n402), .A(n412) );
  nor02 U480 ( .Y(n413), .A0(n398), .A1(n400) );
  inv02 U481 ( .Y(n403), .A(n413) );
  nor02 U482 ( .Y(n414), .A0(n404), .A1(n405) );
  inv01 U483 ( .Y(n407), .A(n414) );
  inv02 U484 ( .Y(carry_33_), .A(n416) );
  inv02 U485 ( .Y(n417), .A(B[32]) );
  inv02 U486 ( .Y(n418), .A(A[32]) );
  inv04 U487 ( .Y(n419), .A(carry_32_) );
  nor02 U488 ( .Y(n420), .A0(n417), .A1(n421) );
  nor02 U489 ( .Y(n422), .A0(n418), .A1(n423) );
  nor02 U490 ( .Y(n424), .A0(n419), .A1(n425) );
  nor02 U491 ( .Y(n426), .A0(n419), .A1(n427) );
  nor02 U492 ( .Y(n415), .A0(n428), .A1(n429) );
  nor02 U493 ( .Y(n430), .A0(n418), .A1(n419) );
  nor02 U494 ( .Y(n431), .A0(n417), .A1(n419) );
  nor02 U495 ( .Y(n432), .A0(n417), .A1(n418) );
  nor02 U496 ( .Y(n416), .A0(n432), .A1(n433) );
  nor02 U497 ( .Y(n434), .A0(A[32]), .A1(carry_32_) );
  inv01 U498 ( .Y(n421), .A(n434) );
  nor02 U499 ( .Y(n435), .A0(B[32]), .A1(carry_32_) );
  inv01 U500 ( .Y(n423), .A(n435) );
  nor02 U501 ( .Y(n436), .A0(B[32]), .A1(A[32]) );
  inv01 U502 ( .Y(n425), .A(n436) );
  nor02 U503 ( .Y(n437), .A0(n417), .A1(n418) );
  inv01 U504 ( .Y(n427), .A(n437) );
  nor02 U505 ( .Y(n438), .A0(n420), .A1(n422) );
  inv02 U506 ( .Y(n428), .A(n438) );
  nor02 U507 ( .Y(n439), .A0(n424), .A1(n426) );
  inv02 U508 ( .Y(n429), .A(n439) );
  nor02 U509 ( .Y(n440), .A0(n430), .A1(n431) );
  inv01 U510 ( .Y(n433), .A(n440) );
  inv02 U511 ( .Y(carry_50_), .A(n442) );
  inv02 U512 ( .Y(n443), .A(B[49]) );
  inv02 U513 ( .Y(n444), .A(A[49]) );
  inv04 U514 ( .Y(n445), .A(carry_49_) );
  nor02 U515 ( .Y(n446), .A0(n443), .A1(n447) );
  nor02 U516 ( .Y(n448), .A0(n444), .A1(n449) );
  nor02 U517 ( .Y(n450), .A0(n445), .A1(n451) );
  nor02 U518 ( .Y(n452), .A0(n445), .A1(n453) );
  nor02 U519 ( .Y(n441), .A0(n454), .A1(n455) );
  nor02 U520 ( .Y(n456), .A0(n444), .A1(n445) );
  nor02 U521 ( .Y(n457), .A0(n443), .A1(n445) );
  nor02 U522 ( .Y(n458), .A0(n443), .A1(n444) );
  nor02 U523 ( .Y(n442), .A0(n458), .A1(n459) );
  nor02 U524 ( .Y(n460), .A0(A[49]), .A1(carry_49_) );
  inv01 U525 ( .Y(n447), .A(n460) );
  nor02 U526 ( .Y(n461), .A0(B[49]), .A1(carry_49_) );
  inv01 U527 ( .Y(n449), .A(n461) );
  nor02 U528 ( .Y(n462), .A0(B[49]), .A1(A[49]) );
  inv01 U529 ( .Y(n451), .A(n462) );
  nor02 U530 ( .Y(n463), .A0(n443), .A1(n444) );
  inv01 U531 ( .Y(n453), .A(n463) );
  nor02 U532 ( .Y(n464), .A0(n446), .A1(n448) );
  inv02 U533 ( .Y(n454), .A(n464) );
  nor02 U534 ( .Y(n465), .A0(n450), .A1(n452) );
  inv02 U535 ( .Y(n455), .A(n465) );
  nor02 U536 ( .Y(n466), .A0(n456), .A1(n457) );
  inv01 U537 ( .Y(n459), .A(n466) );
  inv02 U538 ( .Y(carry_47_), .A(n468) );
  inv02 U539 ( .Y(n469), .A(B[46]) );
  inv02 U540 ( .Y(n470), .A(A[46]) );
  inv04 U541 ( .Y(n471), .A(carry_46_) );
  nor02 U542 ( .Y(n472), .A0(n469), .A1(n473) );
  nor02 U543 ( .Y(n474), .A0(n470), .A1(n475) );
  nor02 U544 ( .Y(n476), .A0(n471), .A1(n477) );
  nor02 U545 ( .Y(n478), .A0(n471), .A1(n479) );
  nor02 U546 ( .Y(n467), .A0(n480), .A1(n481) );
  nor02 U547 ( .Y(n482), .A0(n470), .A1(n471) );
  nor02 U548 ( .Y(n483), .A0(n469), .A1(n471) );
  nor02 U549 ( .Y(n484), .A0(n469), .A1(n470) );
  nor02 U550 ( .Y(n468), .A0(n484), .A1(n485) );
  nor02 U551 ( .Y(n486), .A0(A[46]), .A1(carry_46_) );
  inv01 U552 ( .Y(n473), .A(n486) );
  nor02 U553 ( .Y(n487), .A0(B[46]), .A1(carry_46_) );
  inv01 U554 ( .Y(n475), .A(n487) );
  nor02 U555 ( .Y(n488), .A0(B[46]), .A1(A[46]) );
  inv01 U556 ( .Y(n477), .A(n488) );
  nor02 U557 ( .Y(n489), .A0(n469), .A1(n470) );
  inv01 U558 ( .Y(n479), .A(n489) );
  nor02 U559 ( .Y(n490), .A0(n472), .A1(n474) );
  inv02 U560 ( .Y(n480), .A(n490) );
  nor02 U561 ( .Y(n491), .A0(n476), .A1(n478) );
  inv02 U562 ( .Y(n481), .A(n491) );
  nor02 U563 ( .Y(n492), .A0(n482), .A1(n483) );
  inv01 U564 ( .Y(n485), .A(n492) );
  inv02 U565 ( .Y(carry_29_), .A(n494) );
  inv02 U566 ( .Y(n495), .A(B[28]) );
  inv02 U567 ( .Y(n496), .A(A[28]) );
  inv04 U568 ( .Y(n497), .A(carry_28_) );
  nor02 U569 ( .Y(n498), .A0(n495), .A1(n499) );
  nor02 U570 ( .Y(n500), .A0(n496), .A1(n501) );
  nor02 U571 ( .Y(n502), .A0(n497), .A1(n503) );
  nor02 U572 ( .Y(n504), .A0(n497), .A1(n505) );
  nor02 U573 ( .Y(n493), .A0(n506), .A1(n507) );
  nor02 U574 ( .Y(n508), .A0(n496), .A1(n497) );
  nor02 U575 ( .Y(n509), .A0(n495), .A1(n497) );
  nor02 U576 ( .Y(n510), .A0(n495), .A1(n496) );
  nor02 U577 ( .Y(n494), .A0(n510), .A1(n511) );
  nor02 U578 ( .Y(n512), .A0(A[28]), .A1(carry_28_) );
  inv01 U579 ( .Y(n499), .A(n512) );
  nor02 U580 ( .Y(n513), .A0(B[28]), .A1(carry_28_) );
  inv01 U581 ( .Y(n501), .A(n513) );
  nor02 U582 ( .Y(n514), .A0(B[28]), .A1(A[28]) );
  inv01 U583 ( .Y(n503), .A(n514) );
  nor02 U584 ( .Y(n515), .A0(n495), .A1(n496) );
  inv01 U585 ( .Y(n505), .A(n515) );
  nor02 U586 ( .Y(n516), .A0(n498), .A1(n500) );
  inv02 U587 ( .Y(n506), .A(n516) );
  nor02 U588 ( .Y(n517), .A0(n502), .A1(n504) );
  inv02 U589 ( .Y(n507), .A(n517) );
  nor02 U590 ( .Y(n518), .A0(n508), .A1(n509) );
  inv01 U591 ( .Y(n511), .A(n518) );
  inv02 U592 ( .Y(carry_31_), .A(n520) );
  inv02 U593 ( .Y(n521), .A(B[30]) );
  inv02 U594 ( .Y(n522), .A(A[30]) );
  inv04 U595 ( .Y(n523), .A(carry_30_) );
  nor02 U596 ( .Y(n524), .A0(n521), .A1(n525) );
  nor02 U597 ( .Y(n526), .A0(n522), .A1(n527) );
  nor02 U598 ( .Y(n528), .A0(n523), .A1(n529) );
  nor02 U599 ( .Y(n530), .A0(n523), .A1(n531) );
  nor02 U600 ( .Y(n519), .A0(n532), .A1(n533) );
  nor02 U601 ( .Y(n534), .A0(n522), .A1(n523) );
  nor02 U602 ( .Y(n535), .A0(n521), .A1(n523) );
  nor02 U603 ( .Y(n536), .A0(n521), .A1(n522) );
  nor02 U604 ( .Y(n520), .A0(n536), .A1(n537) );
  nor02 U605 ( .Y(n538), .A0(A[30]), .A1(carry_30_) );
  inv01 U606 ( .Y(n525), .A(n538) );
  nor02 U607 ( .Y(n539), .A0(B[30]), .A1(carry_30_) );
  inv01 U608 ( .Y(n527), .A(n539) );
  nor02 U609 ( .Y(n540), .A0(B[30]), .A1(A[30]) );
  inv01 U610 ( .Y(n529), .A(n540) );
  nor02 U611 ( .Y(n541), .A0(n521), .A1(n522) );
  inv01 U612 ( .Y(n531), .A(n541) );
  nor02 U613 ( .Y(n542), .A0(n524), .A1(n526) );
  inv02 U614 ( .Y(n532), .A(n542) );
  nor02 U615 ( .Y(n543), .A0(n528), .A1(n530) );
  inv02 U616 ( .Y(n533), .A(n543) );
  nor02 U617 ( .Y(n544), .A0(n534), .A1(n535) );
  inv01 U618 ( .Y(n537), .A(n544) );
  inv02 U619 ( .Y(carry_48_), .A(n546) );
  inv02 U620 ( .Y(n547), .A(B[47]) );
  inv02 U621 ( .Y(n548), .A(A[47]) );
  inv04 U622 ( .Y(n549), .A(carry_47_) );
  nor02 U623 ( .Y(n550), .A0(n547), .A1(n551) );
  nor02 U624 ( .Y(n552), .A0(n548), .A1(n553) );
  nor02 U625 ( .Y(n554), .A0(n549), .A1(n555) );
  nor02 U626 ( .Y(n556), .A0(n549), .A1(n557) );
  nor02 U627 ( .Y(n545), .A0(n558), .A1(n559) );
  nor02 U628 ( .Y(n560), .A0(n548), .A1(n549) );
  nor02 U629 ( .Y(n561), .A0(n547), .A1(n549) );
  nor02 U630 ( .Y(n562), .A0(n547), .A1(n548) );
  nor02 U631 ( .Y(n546), .A0(n562), .A1(n563) );
  nor02 U632 ( .Y(n564), .A0(A[47]), .A1(carry_47_) );
  inv01 U633 ( .Y(n551), .A(n564) );
  nor02 U634 ( .Y(n565), .A0(B[47]), .A1(carry_47_) );
  inv01 U635 ( .Y(n553), .A(n565) );
  nor02 U636 ( .Y(n566), .A0(B[47]), .A1(A[47]) );
  inv01 U637 ( .Y(n555), .A(n566) );
  nor02 U638 ( .Y(n567), .A0(n547), .A1(n548) );
  inv01 U639 ( .Y(n557), .A(n567) );
  nor02 U640 ( .Y(n568), .A0(n550), .A1(n552) );
  inv02 U641 ( .Y(n558), .A(n568) );
  nor02 U642 ( .Y(n569), .A0(n554), .A1(n556) );
  inv02 U643 ( .Y(n559), .A(n569) );
  nor02 U644 ( .Y(n570), .A0(n560), .A1(n561) );
  inv01 U645 ( .Y(n563), .A(n570) );
  inv02 U646 ( .Y(carry_27_), .A(n572) );
  inv02 U647 ( .Y(n573), .A(B[26]) );
  inv02 U648 ( .Y(n574), .A(A[26]) );
  inv04 U649 ( .Y(n575), .A(carry_26_) );
  nor02 U650 ( .Y(n576), .A0(n573), .A1(n577) );
  nor02 U651 ( .Y(n578), .A0(n574), .A1(n579) );
  nor02 U652 ( .Y(n580), .A0(n575), .A1(n581) );
  nor02 U653 ( .Y(n582), .A0(n575), .A1(n583) );
  nor02 U654 ( .Y(n571), .A0(n584), .A1(n585) );
  nor02 U655 ( .Y(n586), .A0(n574), .A1(n575) );
  nor02 U656 ( .Y(n587), .A0(n573), .A1(n575) );
  nor02 U657 ( .Y(n588), .A0(n573), .A1(n574) );
  nor02 U658 ( .Y(n572), .A0(n588), .A1(n589) );
  nor02 U659 ( .Y(n590), .A0(A[26]), .A1(carry_26_) );
  inv01 U660 ( .Y(n577), .A(n590) );
  nor02 U661 ( .Y(n591), .A0(B[26]), .A1(carry_26_) );
  inv01 U662 ( .Y(n579), .A(n591) );
  nor02 U663 ( .Y(n592), .A0(B[26]), .A1(A[26]) );
  inv01 U664 ( .Y(n581), .A(n592) );
  nor02 U665 ( .Y(n593), .A0(n573), .A1(n574) );
  inv01 U666 ( .Y(n583), .A(n593) );
  nor02 U667 ( .Y(n594), .A0(n576), .A1(n578) );
  inv02 U668 ( .Y(n584), .A(n594) );
  nor02 U669 ( .Y(n595), .A0(n580), .A1(n582) );
  inv02 U670 ( .Y(n585), .A(n595) );
  nor02 U671 ( .Y(n596), .A0(n586), .A1(n587) );
  inv01 U672 ( .Y(n589), .A(n596) );
  inv02 U673 ( .Y(carry_28_), .A(n598) );
  inv02 U674 ( .Y(n599), .A(B[27]) );
  inv02 U675 ( .Y(n600), .A(A[27]) );
  inv04 U676 ( .Y(n601), .A(carry_27_) );
  nor02 U677 ( .Y(n602), .A0(n599), .A1(n603) );
  nor02 U678 ( .Y(n604), .A0(n600), .A1(n605) );
  nor02 U679 ( .Y(n606), .A0(n601), .A1(n607) );
  nor02 U680 ( .Y(n608), .A0(n601), .A1(n609) );
  nor02 U681 ( .Y(n597), .A0(n610), .A1(n611) );
  nor02 U682 ( .Y(n612), .A0(n600), .A1(n601) );
  nor02 U683 ( .Y(n613), .A0(n599), .A1(n601) );
  nor02 U684 ( .Y(n614), .A0(n599), .A1(n600) );
  nor02 U685 ( .Y(n598), .A0(n614), .A1(n615) );
  nor02 U686 ( .Y(n616), .A0(A[27]), .A1(carry_27_) );
  inv01 U687 ( .Y(n603), .A(n616) );
  nor02 U688 ( .Y(n617), .A0(B[27]), .A1(carry_27_) );
  inv01 U689 ( .Y(n605), .A(n617) );
  nor02 U690 ( .Y(n618), .A0(B[27]), .A1(A[27]) );
  inv01 U691 ( .Y(n607), .A(n618) );
  nor02 U692 ( .Y(n619), .A0(n599), .A1(n600) );
  inv01 U693 ( .Y(n609), .A(n619) );
  nor02 U694 ( .Y(n620), .A0(n602), .A1(n604) );
  inv02 U695 ( .Y(n610), .A(n620) );
  nor02 U696 ( .Y(n621), .A0(n606), .A1(n608) );
  inv02 U697 ( .Y(n611), .A(n621) );
  nor02 U698 ( .Y(n622), .A0(n612), .A1(n613) );
  inv01 U699 ( .Y(n615), .A(n622) );
  inv02 U700 ( .Y(carry_46_), .A(n624) );
  inv02 U701 ( .Y(n625), .A(B[45]) );
  inv02 U702 ( .Y(n626), .A(A[45]) );
  inv02 U703 ( .Y(n627), .A(carry_45_) );
  nor02 U704 ( .Y(n628), .A0(n625), .A1(n629) );
  nor02 U705 ( .Y(n630), .A0(n626), .A1(n631) );
  nor02 U706 ( .Y(n632), .A0(n627), .A1(n633) );
  nor02 U707 ( .Y(n634), .A0(n627), .A1(n635) );
  nor02 U708 ( .Y(n623), .A0(n636), .A1(n637) );
  nor02 U709 ( .Y(n638), .A0(n626), .A1(n627) );
  nor02 U710 ( .Y(n639), .A0(n625), .A1(n627) );
  nor02 U711 ( .Y(n640), .A0(n625), .A1(n626) );
  nor02 U712 ( .Y(n624), .A0(n640), .A1(n641) );
  nor02 U713 ( .Y(n642), .A0(A[45]), .A1(carry_45_) );
  inv01 U714 ( .Y(n629), .A(n642) );
  nor02 U715 ( .Y(n643), .A0(B[45]), .A1(carry_45_) );
  inv01 U716 ( .Y(n631), .A(n643) );
  nor02 U717 ( .Y(n644), .A0(B[45]), .A1(A[45]) );
  inv01 U718 ( .Y(n633), .A(n644) );
  nor02 U719 ( .Y(n645), .A0(n625), .A1(n626) );
  inv01 U720 ( .Y(n635), .A(n645) );
  nor02 U721 ( .Y(n646), .A0(n628), .A1(n630) );
  inv02 U722 ( .Y(n636), .A(n646) );
  nor02 U723 ( .Y(n647), .A0(n632), .A1(n634) );
  inv02 U724 ( .Y(n637), .A(n647) );
  nor02 U725 ( .Y(n648), .A0(n638), .A1(n639) );
  inv01 U726 ( .Y(n641), .A(n648) );
  inv02 U727 ( .Y(carry_30_), .A(n650) );
  inv02 U728 ( .Y(n651), .A(B[29]) );
  inv02 U729 ( .Y(n652), .A(A[29]) );
  inv02 U730 ( .Y(n653), .A(carry_29_) );
  nor02 U731 ( .Y(n654), .A0(n651), .A1(n655) );
  nor02 U732 ( .Y(n656), .A0(n652), .A1(n657) );
  nor02 U733 ( .Y(n658), .A0(n653), .A1(n659) );
  nor02 U734 ( .Y(n660), .A0(n653), .A1(n661) );
  nor02 U735 ( .Y(n649), .A0(n662), .A1(n663) );
  nor02 U736 ( .Y(n664), .A0(n652), .A1(n653) );
  nor02 U737 ( .Y(n665), .A0(n651), .A1(n653) );
  nor02 U738 ( .Y(n666), .A0(n651), .A1(n652) );
  nor02 U739 ( .Y(n650), .A0(n666), .A1(n667) );
  nor02 U740 ( .Y(n668), .A0(A[29]), .A1(carry_29_) );
  inv01 U741 ( .Y(n655), .A(n668) );
  nor02 U742 ( .Y(n669), .A0(B[29]), .A1(carry_29_) );
  inv01 U743 ( .Y(n657), .A(n669) );
  nor02 U744 ( .Y(n670), .A0(B[29]), .A1(A[29]) );
  inv01 U745 ( .Y(n659), .A(n670) );
  nor02 U746 ( .Y(n671), .A0(n651), .A1(n652) );
  inv01 U747 ( .Y(n661), .A(n671) );
  nor02 U748 ( .Y(n672), .A0(n654), .A1(n656) );
  inv02 U749 ( .Y(n662), .A(n672) );
  nor02 U750 ( .Y(n673), .A0(n658), .A1(n660) );
  inv02 U751 ( .Y(n663), .A(n673) );
  nor02 U752 ( .Y(n674), .A0(n664), .A1(n665) );
  inv01 U753 ( .Y(n667), .A(n674) );
  inv02 U754 ( .Y(carry_11_), .A(n676) );
  inv02 U755 ( .Y(n677), .A(B[10]) );
  inv02 U756 ( .Y(n678), .A(A[10]) );
  inv04 U757 ( .Y(n679), .A(carry_10_) );
  nor02 U758 ( .Y(n680), .A0(n677), .A1(n681) );
  nor02 U759 ( .Y(n682), .A0(n678), .A1(n683) );
  nor02 U760 ( .Y(n684), .A0(n679), .A1(n685) );
  nor02 U761 ( .Y(n686), .A0(n679), .A1(n687) );
  nor02 U762 ( .Y(n675), .A0(n688), .A1(n689) );
  nor02 U763 ( .Y(n690), .A0(n678), .A1(n679) );
  nor02 U764 ( .Y(n691), .A0(n677), .A1(n679) );
  nor02 U765 ( .Y(n692), .A0(n677), .A1(n678) );
  nor02 U766 ( .Y(n676), .A0(n692), .A1(n693) );
  nor02 U767 ( .Y(n694), .A0(A[10]), .A1(carry_10_) );
  inv01 U768 ( .Y(n681), .A(n694) );
  nor02 U769 ( .Y(n695), .A0(B[10]), .A1(carry_10_) );
  inv01 U770 ( .Y(n683), .A(n695) );
  nor02 U771 ( .Y(n696), .A0(B[10]), .A1(A[10]) );
  inv01 U772 ( .Y(n685), .A(n696) );
  nor02 U773 ( .Y(n697), .A0(n677), .A1(n678) );
  inv01 U774 ( .Y(n687), .A(n697) );
  nor02 U775 ( .Y(n698), .A0(n680), .A1(n682) );
  inv02 U776 ( .Y(n688), .A(n698) );
  nor02 U777 ( .Y(n699), .A0(n684), .A1(n686) );
  inv02 U778 ( .Y(n689), .A(n699) );
  nor02 U779 ( .Y(n700), .A0(n690), .A1(n691) );
  inv01 U780 ( .Y(n693), .A(n700) );
  inv02 U781 ( .Y(carry_25_), .A(n702) );
  inv02 U782 ( .Y(n703), .A(B[24]) );
  inv02 U783 ( .Y(n704), .A(A[24]) );
  inv04 U784 ( .Y(n705), .A(carry_24_) );
  nor02 U785 ( .Y(n706), .A0(n703), .A1(n707) );
  nor02 U786 ( .Y(n708), .A0(n704), .A1(n709) );
  nor02 U787 ( .Y(n710), .A0(n705), .A1(n711) );
  nor02 U788 ( .Y(n712), .A0(n705), .A1(n713) );
  nor02 U789 ( .Y(n701), .A0(n714), .A1(n715) );
  nor02 U790 ( .Y(n716), .A0(n704), .A1(n705) );
  nor02 U791 ( .Y(n717), .A0(n703), .A1(n705) );
  nor02 U792 ( .Y(n718), .A0(n703), .A1(n704) );
  nor02 U793 ( .Y(n702), .A0(n718), .A1(n719) );
  nor02 U794 ( .Y(n720), .A0(A[24]), .A1(carry_24_) );
  inv01 U795 ( .Y(n707), .A(n720) );
  nor02 U796 ( .Y(n721), .A0(B[24]), .A1(carry_24_) );
  inv01 U797 ( .Y(n709), .A(n721) );
  nor02 U798 ( .Y(n722), .A0(B[24]), .A1(A[24]) );
  inv01 U799 ( .Y(n711), .A(n722) );
  nor02 U800 ( .Y(n723), .A0(n703), .A1(n704) );
  inv01 U801 ( .Y(n713), .A(n723) );
  nor02 U802 ( .Y(n724), .A0(n706), .A1(n708) );
  inv02 U803 ( .Y(n714), .A(n724) );
  nor02 U804 ( .Y(n725), .A0(n710), .A1(n712) );
  inv02 U805 ( .Y(n715), .A(n725) );
  nor02 U806 ( .Y(n726), .A0(n716), .A1(n717) );
  inv01 U807 ( .Y(n719), .A(n726) );
  inv02 U808 ( .Y(carry_26_), .A(n728) );
  inv02 U809 ( .Y(n729), .A(B[25]) );
  inv02 U810 ( .Y(n730), .A(A[25]) );
  inv04 U811 ( .Y(n731), .A(carry_25_) );
  nor02 U812 ( .Y(n732), .A0(n729), .A1(n733) );
  nor02 U813 ( .Y(n734), .A0(n730), .A1(n735) );
  nor02 U814 ( .Y(n736), .A0(n731), .A1(n737) );
  nor02 U815 ( .Y(n738), .A0(n731), .A1(n739) );
  nor02 U816 ( .Y(n727), .A0(n740), .A1(n741) );
  nor02 U817 ( .Y(n742), .A0(n730), .A1(n731) );
  nor02 U818 ( .Y(n743), .A0(n729), .A1(n731) );
  nor02 U819 ( .Y(n744), .A0(n729), .A1(n730) );
  nor02 U820 ( .Y(n728), .A0(n744), .A1(n745) );
  nor02 U821 ( .Y(n746), .A0(A[25]), .A1(carry_25_) );
  inv01 U822 ( .Y(n733), .A(n746) );
  nor02 U823 ( .Y(n747), .A0(B[25]), .A1(carry_25_) );
  inv01 U824 ( .Y(n735), .A(n747) );
  nor02 U825 ( .Y(n748), .A0(B[25]), .A1(A[25]) );
  inv01 U826 ( .Y(n737), .A(n748) );
  nor02 U827 ( .Y(n749), .A0(n729), .A1(n730) );
  inv01 U828 ( .Y(n739), .A(n749) );
  nor02 U829 ( .Y(n750), .A0(n732), .A1(n734) );
  inv02 U830 ( .Y(n740), .A(n750) );
  nor02 U831 ( .Y(n751), .A0(n736), .A1(n738) );
  inv02 U832 ( .Y(n741), .A(n751) );
  nor02 U833 ( .Y(n752), .A0(n742), .A1(n743) );
  inv01 U834 ( .Y(n745), .A(n752) );
  inv02 U835 ( .Y(carry_12_), .A(n754) );
  inv02 U836 ( .Y(n755), .A(B[11]) );
  inv02 U837 ( .Y(n756), .A(A[11]) );
  inv04 U838 ( .Y(n757), .A(carry_11_) );
  nor02 U839 ( .Y(n758), .A0(n755), .A1(n759) );
  nor02 U840 ( .Y(n760), .A0(n756), .A1(n761) );
  nor02 U841 ( .Y(n762), .A0(n757), .A1(n763) );
  nor02 U842 ( .Y(n764), .A0(n757), .A1(n765) );
  nor02 U843 ( .Y(n753), .A0(n766), .A1(n767) );
  nor02 U844 ( .Y(n768), .A0(n756), .A1(n757) );
  nor02 U845 ( .Y(n769), .A0(n755), .A1(n757) );
  nor02 U846 ( .Y(n770), .A0(n755), .A1(n756) );
  nor02 U847 ( .Y(n754), .A0(n770), .A1(n771) );
  nor02 U848 ( .Y(n772), .A0(A[11]), .A1(carry_11_) );
  inv01 U849 ( .Y(n759), .A(n772) );
  nor02 U850 ( .Y(n773), .A0(B[11]), .A1(carry_11_) );
  inv01 U851 ( .Y(n761), .A(n773) );
  nor02 U852 ( .Y(n774), .A0(B[11]), .A1(A[11]) );
  inv01 U853 ( .Y(n763), .A(n774) );
  nor02 U854 ( .Y(n775), .A0(n755), .A1(n756) );
  inv01 U855 ( .Y(n765), .A(n775) );
  nor02 U856 ( .Y(n776), .A0(n758), .A1(n760) );
  inv02 U857 ( .Y(n766), .A(n776) );
  nor02 U858 ( .Y(n777), .A0(n762), .A1(n764) );
  inv02 U859 ( .Y(n767), .A(n777) );
  nor02 U860 ( .Y(n778), .A0(n768), .A1(n769) );
  inv01 U861 ( .Y(n771), .A(n778) );
  inv02 U862 ( .Y(carry_9_), .A(n780) );
  inv02 U863 ( .Y(n781), .A(B[8]) );
  inv02 U864 ( .Y(n782), .A(A[8]) );
  inv04 U865 ( .Y(n783), .A(carry_8_) );
  nor02 U866 ( .Y(n784), .A0(n781), .A1(n785) );
  nor02 U867 ( .Y(n786), .A0(n782), .A1(n787) );
  nor02 U868 ( .Y(n788), .A0(n783), .A1(n789) );
  nor02 U869 ( .Y(n790), .A0(n783), .A1(n791) );
  nor02 U870 ( .Y(n779), .A0(n792), .A1(n793) );
  nor02 U871 ( .Y(n794), .A0(n782), .A1(n783) );
  nor02 U872 ( .Y(n795), .A0(n781), .A1(n783) );
  nor02 U873 ( .Y(n796), .A0(n781), .A1(n782) );
  nor02 U874 ( .Y(n780), .A0(n796), .A1(n797) );
  nor02 U875 ( .Y(n798), .A0(A[8]), .A1(carry_8_) );
  inv01 U876 ( .Y(n785), .A(n798) );
  nor02 U877 ( .Y(n799), .A0(B[8]), .A1(carry_8_) );
  inv01 U878 ( .Y(n787), .A(n799) );
  nor02 U879 ( .Y(n800), .A0(B[8]), .A1(A[8]) );
  inv01 U880 ( .Y(n789), .A(n800) );
  nor02 U881 ( .Y(n801), .A0(n781), .A1(n782) );
  inv01 U882 ( .Y(n791), .A(n801) );
  nor02 U883 ( .Y(n802), .A0(n784), .A1(n786) );
  inv02 U884 ( .Y(n792), .A(n802) );
  nor02 U885 ( .Y(n803), .A0(n788), .A1(n790) );
  inv02 U886 ( .Y(n793), .A(n803) );
  nor02 U887 ( .Y(n804), .A0(n794), .A1(n795) );
  inv01 U888 ( .Y(n797), .A(n804) );
  inv02 U889 ( .Y(carry_23_), .A(n806) );
  inv02 U890 ( .Y(n807), .A(B[22]) );
  inv02 U891 ( .Y(n808), .A(A[22]) );
  inv04 U892 ( .Y(n809), .A(carry_22_) );
  nor02 U893 ( .Y(n810), .A0(n807), .A1(n811) );
  nor02 U894 ( .Y(n812), .A0(n808), .A1(n813) );
  nor02 U895 ( .Y(n814), .A0(n809), .A1(n815) );
  nor02 U896 ( .Y(n816), .A0(n809), .A1(n817) );
  nor02 U897 ( .Y(n805), .A0(n818), .A1(n819) );
  nor02 U898 ( .Y(n820), .A0(n808), .A1(n809) );
  nor02 U899 ( .Y(n821), .A0(n807), .A1(n809) );
  nor02 U900 ( .Y(n822), .A0(n807), .A1(n808) );
  nor02 U901 ( .Y(n806), .A0(n822), .A1(n823) );
  nor02 U902 ( .Y(n824), .A0(A[22]), .A1(carry_22_) );
  inv01 U903 ( .Y(n811), .A(n824) );
  nor02 U904 ( .Y(n825), .A0(B[22]), .A1(carry_22_) );
  inv01 U905 ( .Y(n813), .A(n825) );
  nor02 U906 ( .Y(n826), .A0(B[22]), .A1(A[22]) );
  inv01 U907 ( .Y(n815), .A(n826) );
  nor02 U908 ( .Y(n827), .A0(n807), .A1(n808) );
  inv01 U909 ( .Y(n817), .A(n827) );
  nor02 U910 ( .Y(n828), .A0(n810), .A1(n812) );
  inv02 U911 ( .Y(n818), .A(n828) );
  nor02 U912 ( .Y(n829), .A0(n814), .A1(n816) );
  inv02 U913 ( .Y(n819), .A(n829) );
  nor02 U914 ( .Y(n830), .A0(n820), .A1(n821) );
  inv01 U915 ( .Y(n823), .A(n830) );
  inv02 U916 ( .Y(carry_24_), .A(n832) );
  inv02 U917 ( .Y(n833), .A(B[23]) );
  inv02 U918 ( .Y(n834), .A(A[23]) );
  inv04 U919 ( .Y(n835), .A(carry_23_) );
  nor02 U920 ( .Y(n836), .A0(n833), .A1(n837) );
  nor02 U921 ( .Y(n838), .A0(n834), .A1(n839) );
  nor02 U922 ( .Y(n840), .A0(n835), .A1(n841) );
  nor02 U923 ( .Y(n842), .A0(n835), .A1(n843) );
  nor02 U924 ( .Y(n831), .A0(n844), .A1(n845) );
  nor02 U925 ( .Y(n846), .A0(n834), .A1(n835) );
  nor02 U926 ( .Y(n847), .A0(n833), .A1(n835) );
  nor02 U927 ( .Y(n848), .A0(n833), .A1(n834) );
  nor02 U928 ( .Y(n832), .A0(n848), .A1(n849) );
  nor02 U929 ( .Y(n850), .A0(A[23]), .A1(carry_23_) );
  inv01 U930 ( .Y(n837), .A(n850) );
  nor02 U931 ( .Y(n851), .A0(B[23]), .A1(carry_23_) );
  inv01 U932 ( .Y(n839), .A(n851) );
  nor02 U933 ( .Y(n852), .A0(B[23]), .A1(A[23]) );
  inv01 U934 ( .Y(n841), .A(n852) );
  nor02 U935 ( .Y(n853), .A0(n833), .A1(n834) );
  inv01 U936 ( .Y(n843), .A(n853) );
  nor02 U937 ( .Y(n854), .A0(n836), .A1(n838) );
  inv02 U938 ( .Y(n844), .A(n854) );
  nor02 U939 ( .Y(n855), .A0(n840), .A1(n842) );
  inv02 U940 ( .Y(n845), .A(n855) );
  nor02 U941 ( .Y(n856), .A0(n846), .A1(n847) );
  inv01 U942 ( .Y(n849), .A(n856) );
  inv02 U943 ( .Y(carry_10_), .A(n858) );
  inv02 U944 ( .Y(n859), .A(B[9]) );
  inv02 U945 ( .Y(n860), .A(A[9]) );
  inv04 U946 ( .Y(n861), .A(carry_9_) );
  nor02 U947 ( .Y(n862), .A0(n859), .A1(n863) );
  nor02 U948 ( .Y(n864), .A0(n860), .A1(n865) );
  nor02 U949 ( .Y(n866), .A0(n861), .A1(n867) );
  nor02 U950 ( .Y(n868), .A0(n861), .A1(n869) );
  nor02 U951 ( .Y(n857), .A0(n870), .A1(n871) );
  nor02 U952 ( .Y(n872), .A0(n860), .A1(n861) );
  nor02 U953 ( .Y(n873), .A0(n859), .A1(n861) );
  nor02 U954 ( .Y(n874), .A0(n859), .A1(n860) );
  nor02 U955 ( .Y(n858), .A0(n874), .A1(n875) );
  nor02 U956 ( .Y(n876), .A0(A[9]), .A1(carry_9_) );
  inv01 U957 ( .Y(n863), .A(n876) );
  nor02 U958 ( .Y(n877), .A0(B[9]), .A1(carry_9_) );
  inv01 U959 ( .Y(n865), .A(n877) );
  nor02 U960 ( .Y(n878), .A0(B[9]), .A1(A[9]) );
  inv01 U961 ( .Y(n867), .A(n878) );
  nor02 U962 ( .Y(n879), .A0(n859), .A1(n860) );
  inv01 U963 ( .Y(n869), .A(n879) );
  nor02 U964 ( .Y(n880), .A0(n862), .A1(n864) );
  inv02 U965 ( .Y(n870), .A(n880) );
  nor02 U966 ( .Y(n881), .A0(n866), .A1(n868) );
  inv02 U967 ( .Y(n871), .A(n881) );
  nor02 U968 ( .Y(n882), .A0(n872), .A1(n873) );
  inv01 U969 ( .Y(n875), .A(n882) );
  inv02 U970 ( .Y(carry_7_), .A(n884) );
  inv02 U971 ( .Y(n885), .A(B[6]) );
  inv02 U972 ( .Y(n886), .A(A[6]) );
  inv04 U973 ( .Y(n887), .A(carry_6_) );
  nor02 U974 ( .Y(n888), .A0(n885), .A1(n889) );
  nor02 U975 ( .Y(n890), .A0(n886), .A1(n891) );
  nor02 U976 ( .Y(n892), .A0(n887), .A1(n893) );
  nor02 U977 ( .Y(n894), .A0(n887), .A1(n895) );
  nor02 U978 ( .Y(n883), .A0(n896), .A1(n897) );
  nor02 U979 ( .Y(n898), .A0(n886), .A1(n887) );
  nor02 U980 ( .Y(n899), .A0(n885), .A1(n887) );
  nor02 U981 ( .Y(n900), .A0(n885), .A1(n886) );
  nor02 U982 ( .Y(n884), .A0(n900), .A1(n901) );
  nor02 U983 ( .Y(n902), .A0(A[6]), .A1(carry_6_) );
  inv01 U984 ( .Y(n889), .A(n902) );
  nor02 U985 ( .Y(n903), .A0(B[6]), .A1(carry_6_) );
  inv01 U986 ( .Y(n891), .A(n903) );
  nor02 U987 ( .Y(n904), .A0(B[6]), .A1(A[6]) );
  inv01 U988 ( .Y(n893), .A(n904) );
  nor02 U989 ( .Y(n905), .A0(n885), .A1(n886) );
  inv01 U990 ( .Y(n895), .A(n905) );
  nor02 U991 ( .Y(n906), .A0(n888), .A1(n890) );
  inv02 U992 ( .Y(n896), .A(n906) );
  nor02 U993 ( .Y(n907), .A0(n892), .A1(n894) );
  inv02 U994 ( .Y(n897), .A(n907) );
  nor02 U995 ( .Y(n908), .A0(n898), .A1(n899) );
  inv01 U996 ( .Y(n901), .A(n908) );
  inv02 U997 ( .Y(carry_21_), .A(n910) );
  inv02 U998 ( .Y(n911), .A(B[20]) );
  inv02 U999 ( .Y(n912), .A(A[20]) );
  inv04 U1000 ( .Y(n913), .A(carry_20_) );
  nor02 U1001 ( .Y(n914), .A0(n911), .A1(n915) );
  nor02 U1002 ( .Y(n916), .A0(n912), .A1(n917) );
  nor02 U1003 ( .Y(n918), .A0(n913), .A1(n919) );
  nor02 U1004 ( .Y(n920), .A0(n913), .A1(n921) );
  nor02 U1005 ( .Y(n909), .A0(n922), .A1(n923) );
  nor02 U1006 ( .Y(n924), .A0(n912), .A1(n913) );
  nor02 U1007 ( .Y(n925), .A0(n911), .A1(n913) );
  nor02 U1008 ( .Y(n926), .A0(n911), .A1(n912) );
  nor02 U1009 ( .Y(n910), .A0(n926), .A1(n927) );
  nor02 U1010 ( .Y(n928), .A0(A[20]), .A1(carry_20_) );
  inv01 U1011 ( .Y(n915), .A(n928) );
  nor02 U1012 ( .Y(n929), .A0(B[20]), .A1(carry_20_) );
  inv01 U1013 ( .Y(n917), .A(n929) );
  nor02 U1014 ( .Y(n930), .A0(B[20]), .A1(A[20]) );
  inv01 U1015 ( .Y(n919), .A(n930) );
  nor02 U1016 ( .Y(n931), .A0(n911), .A1(n912) );
  inv01 U1017 ( .Y(n921), .A(n931) );
  nor02 U1018 ( .Y(n932), .A0(n914), .A1(n916) );
  inv02 U1019 ( .Y(n922), .A(n932) );
  nor02 U1020 ( .Y(n933), .A0(n918), .A1(n920) );
  inv02 U1021 ( .Y(n923), .A(n933) );
  nor02 U1022 ( .Y(n934), .A0(n924), .A1(n925) );
  inv01 U1023 ( .Y(n927), .A(n934) );
  inv02 U1024 ( .Y(carry_8_), .A(n936) );
  inv02 U1025 ( .Y(n937), .A(B[7]) );
  inv02 U1026 ( .Y(n938), .A(A[7]) );
  inv04 U1027 ( .Y(n939), .A(carry_7_) );
  nor02 U1028 ( .Y(n940), .A0(n937), .A1(n941) );
  nor02 U1029 ( .Y(n942), .A0(n938), .A1(n943) );
  nor02 U1030 ( .Y(n944), .A0(n939), .A1(n945) );
  nor02 U1031 ( .Y(n946), .A0(n939), .A1(n947) );
  nor02 U1032 ( .Y(n935), .A0(n948), .A1(n949) );
  nor02 U1033 ( .Y(n950), .A0(n938), .A1(n939) );
  nor02 U1034 ( .Y(n951), .A0(n937), .A1(n939) );
  nor02 U1035 ( .Y(n952), .A0(n937), .A1(n938) );
  nor02 U1036 ( .Y(n936), .A0(n952), .A1(n953) );
  nor02 U1037 ( .Y(n954), .A0(A[7]), .A1(carry_7_) );
  inv01 U1038 ( .Y(n941), .A(n954) );
  nor02 U1039 ( .Y(n955), .A0(B[7]), .A1(carry_7_) );
  inv01 U1040 ( .Y(n943), .A(n955) );
  nor02 U1041 ( .Y(n956), .A0(B[7]), .A1(A[7]) );
  inv01 U1042 ( .Y(n945), .A(n956) );
  nor02 U1043 ( .Y(n957), .A0(n937), .A1(n938) );
  inv01 U1044 ( .Y(n947), .A(n957) );
  nor02 U1045 ( .Y(n958), .A0(n940), .A1(n942) );
  inv02 U1046 ( .Y(n948), .A(n958) );
  nor02 U1047 ( .Y(n959), .A0(n944), .A1(n946) );
  inv02 U1048 ( .Y(n949), .A(n959) );
  nor02 U1049 ( .Y(n960), .A0(n950), .A1(n951) );
  inv01 U1050 ( .Y(n953), .A(n960) );
  inv02 U1051 ( .Y(carry_22_), .A(n962) );
  inv02 U1052 ( .Y(n963), .A(B[21]) );
  inv02 U1053 ( .Y(n964), .A(A[21]) );
  inv04 U1054 ( .Y(n965), .A(carry_21_) );
  nor02 U1055 ( .Y(n966), .A0(n963), .A1(n967) );
  nor02 U1056 ( .Y(n968), .A0(n964), .A1(n969) );
  nor02 U1057 ( .Y(n970), .A0(n965), .A1(n971) );
  nor02 U1058 ( .Y(n972), .A0(n965), .A1(n973) );
  nor02 U1059 ( .Y(n961), .A0(n974), .A1(n975) );
  nor02 U1060 ( .Y(n976), .A0(n964), .A1(n965) );
  nor02 U1061 ( .Y(n977), .A0(n963), .A1(n965) );
  nor02 U1062 ( .Y(n978), .A0(n963), .A1(n964) );
  nor02 U1063 ( .Y(n962), .A0(n978), .A1(n979) );
  nor02 U1064 ( .Y(n980), .A0(A[21]), .A1(carry_21_) );
  inv01 U1065 ( .Y(n967), .A(n980) );
  nor02 U1066 ( .Y(n981), .A0(B[21]), .A1(carry_21_) );
  inv01 U1067 ( .Y(n969), .A(n981) );
  nor02 U1068 ( .Y(n982), .A0(B[21]), .A1(A[21]) );
  inv01 U1069 ( .Y(n971), .A(n982) );
  nor02 U1070 ( .Y(n983), .A0(n963), .A1(n964) );
  inv01 U1071 ( .Y(n973), .A(n983) );
  nor02 U1072 ( .Y(n984), .A0(n966), .A1(n968) );
  inv02 U1073 ( .Y(n974), .A(n984) );
  nor02 U1074 ( .Y(n985), .A0(n970), .A1(n972) );
  inv02 U1075 ( .Y(n975), .A(n985) );
  nor02 U1076 ( .Y(n986), .A0(n976), .A1(n977) );
  inv01 U1077 ( .Y(n979), .A(n986) );
  inv02 U1078 ( .Y(carry_20_), .A(n988) );
  inv02 U1079 ( .Y(n989), .A(B[19]) );
  inv02 U1080 ( .Y(n990), .A(A[19]) );
  inv04 U1081 ( .Y(n991), .A(carry_19_) );
  nor02 U1082 ( .Y(n992), .A0(n989), .A1(n993) );
  nor02 U1083 ( .Y(n994), .A0(n990), .A1(n995) );
  nor02 U1084 ( .Y(n996), .A0(n991), .A1(n997) );
  nor02 U1085 ( .Y(n998), .A0(n991), .A1(n999) );
  nor02 U1086 ( .Y(n987), .A0(n1000), .A1(n1001) );
  nor02 U1087 ( .Y(n1002), .A0(n990), .A1(n991) );
  nor02 U1088 ( .Y(n1003), .A0(n989), .A1(n991) );
  nor02 U1089 ( .Y(n1004), .A0(n989), .A1(n990) );
  nor02 U1090 ( .Y(n988), .A0(n1004), .A1(n1005) );
  nor02 U1091 ( .Y(n1006), .A0(A[19]), .A1(carry_19_) );
  inv01 U1092 ( .Y(n993), .A(n1006) );
  nor02 U1093 ( .Y(n1007), .A0(B[19]), .A1(carry_19_) );
  inv01 U1094 ( .Y(n995), .A(n1007) );
  nor02 U1095 ( .Y(n1008), .A0(B[19]), .A1(A[19]) );
  inv01 U1096 ( .Y(n997), .A(n1008) );
  nor02 U1097 ( .Y(n1009), .A0(n989), .A1(n990) );
  inv01 U1098 ( .Y(n999), .A(n1009) );
  nor02 U1099 ( .Y(n1010), .A0(n992), .A1(n994) );
  inv02 U1100 ( .Y(n1000), .A(n1010) );
  nor02 U1101 ( .Y(n1011), .A0(n996), .A1(n998) );
  inv02 U1102 ( .Y(n1001), .A(n1011) );
  nor02 U1103 ( .Y(n1012), .A0(n1002), .A1(n1003) );
  inv01 U1104 ( .Y(n1005), .A(n1012) );
  inv02 U1105 ( .Y(carry_6_), .A(n1014) );
  inv02 U1106 ( .Y(n1015), .A(B[5]) );
  inv02 U1107 ( .Y(n1016), .A(A[5]) );
  inv04 U1108 ( .Y(n1017), .A(carry_5_) );
  nor02 U1109 ( .Y(n1018), .A0(n1015), .A1(n1019) );
  nor02 U1110 ( .Y(n1020), .A0(n1016), .A1(n1021) );
  nor02 U1111 ( .Y(n1022), .A0(n1017), .A1(n1023) );
  nor02 U1112 ( .Y(n1024), .A0(n1017), .A1(n1025) );
  nor02 U1113 ( .Y(n1013), .A0(n1026), .A1(n1027) );
  nor02 U1114 ( .Y(n1028), .A0(n1016), .A1(n1017) );
  nor02 U1115 ( .Y(n1029), .A0(n1015), .A1(n1017) );
  nor02 U1116 ( .Y(n1030), .A0(n1015), .A1(n1016) );
  nor02 U1117 ( .Y(n1014), .A0(n1030), .A1(n1031) );
  nor02 U1118 ( .Y(n1032), .A0(A[5]), .A1(carry_5_) );
  inv01 U1119 ( .Y(n1019), .A(n1032) );
  nor02 U1120 ( .Y(n1033), .A0(B[5]), .A1(carry_5_) );
  inv01 U1121 ( .Y(n1021), .A(n1033) );
  nor02 U1122 ( .Y(n1034), .A0(B[5]), .A1(A[5]) );
  inv01 U1123 ( .Y(n1023), .A(n1034) );
  nor02 U1124 ( .Y(n1035), .A0(n1015), .A1(n1016) );
  inv01 U1125 ( .Y(n1025), .A(n1035) );
  nor02 U1126 ( .Y(n1036), .A0(n1018), .A1(n1020) );
  inv02 U1127 ( .Y(n1026), .A(n1036) );
  nor02 U1128 ( .Y(n1037), .A0(n1022), .A1(n1024) );
  inv02 U1129 ( .Y(n1027), .A(n1037) );
  nor02 U1130 ( .Y(n1038), .A0(n1028), .A1(n1029) );
  inv01 U1131 ( .Y(n1031), .A(n1038) );
  inv02 U1132 ( .Y(carry_16_), .A(n1040) );
  inv02 U1133 ( .Y(n1041), .A(B[15]) );
  inv02 U1134 ( .Y(n1042), .A(A[15]) );
  inv04 U1135 ( .Y(n1043), .A(carry_15_) );
  nor02 U1136 ( .Y(n1044), .A0(n1041), .A1(n1045) );
  nor02 U1137 ( .Y(n1046), .A0(n1042), .A1(n1047) );
  nor02 U1138 ( .Y(n1048), .A0(n1043), .A1(n1049) );
  nor02 U1139 ( .Y(n1050), .A0(n1043), .A1(n1051) );
  nor02 U1140 ( .Y(n1039), .A0(n1052), .A1(n1053) );
  nor02 U1141 ( .Y(n1054), .A0(n1042), .A1(n1043) );
  nor02 U1142 ( .Y(n1055), .A0(n1041), .A1(n1043) );
  nor02 U1143 ( .Y(n1056), .A0(n1041), .A1(n1042) );
  nor02 U1144 ( .Y(n1040), .A0(n1056), .A1(n1057) );
  nor02 U1145 ( .Y(n1058), .A0(A[15]), .A1(carry_15_) );
  inv01 U1146 ( .Y(n1045), .A(n1058) );
  nor02 U1147 ( .Y(n1059), .A0(B[15]), .A1(carry_15_) );
  inv01 U1148 ( .Y(n1047), .A(n1059) );
  nor02 U1149 ( .Y(n1060), .A0(B[15]), .A1(A[15]) );
  inv01 U1150 ( .Y(n1049), .A(n1060) );
  nor02 U1151 ( .Y(n1061), .A0(n1041), .A1(n1042) );
  inv01 U1152 ( .Y(n1051), .A(n1061) );
  nor02 U1153 ( .Y(n1062), .A0(n1044), .A1(n1046) );
  inv02 U1154 ( .Y(n1052), .A(n1062) );
  nor02 U1155 ( .Y(n1063), .A0(n1048), .A1(n1050) );
  inv02 U1156 ( .Y(n1053), .A(n1063) );
  nor02 U1157 ( .Y(n1064), .A0(n1054), .A1(n1055) );
  inv01 U1158 ( .Y(n1057), .A(n1064) );
  inv02 U1159 ( .Y(carry_17_), .A(n1066) );
  inv02 U1160 ( .Y(n1067), .A(B[16]) );
  inv02 U1161 ( .Y(n1068), .A(A[16]) );
  inv04 U1162 ( .Y(n1069), .A(carry_16_) );
  nor02 U1163 ( .Y(n1070), .A0(n1067), .A1(n1071) );
  nor02 U1164 ( .Y(n1072), .A0(n1068), .A1(n1073) );
  nor02 U1165 ( .Y(n1074), .A0(n1069), .A1(n1075) );
  nor02 U1166 ( .Y(n1076), .A0(n1069), .A1(n1077) );
  nor02 U1167 ( .Y(n1065), .A0(n1078), .A1(n1079) );
  nor02 U1168 ( .Y(n1080), .A0(n1068), .A1(n1069) );
  nor02 U1169 ( .Y(n1081), .A0(n1067), .A1(n1069) );
  nor02 U1170 ( .Y(n1082), .A0(n1067), .A1(n1068) );
  nor02 U1171 ( .Y(n1066), .A0(n1082), .A1(n1083) );
  nor02 U1172 ( .Y(n1084), .A0(A[16]), .A1(carry_16_) );
  inv01 U1173 ( .Y(n1071), .A(n1084) );
  nor02 U1174 ( .Y(n1085), .A0(B[16]), .A1(carry_16_) );
  inv01 U1175 ( .Y(n1073), .A(n1085) );
  nor02 U1176 ( .Y(n1086), .A0(B[16]), .A1(A[16]) );
  inv01 U1177 ( .Y(n1075), .A(n1086) );
  nor02 U1178 ( .Y(n1087), .A0(n1067), .A1(n1068) );
  inv01 U1179 ( .Y(n1077), .A(n1087) );
  nor02 U1180 ( .Y(n1088), .A0(n1070), .A1(n1072) );
  inv02 U1181 ( .Y(n1078), .A(n1088) );
  nor02 U1182 ( .Y(n1089), .A0(n1074), .A1(n1076) );
  inv02 U1183 ( .Y(n1079), .A(n1089) );
  nor02 U1184 ( .Y(n1090), .A0(n1080), .A1(n1081) );
  inv01 U1185 ( .Y(n1083), .A(n1090) );
  inv02 U1186 ( .Y(carry_5_), .A(n1092) );
  inv02 U1187 ( .Y(n1093), .A(B[4]) );
  inv02 U1188 ( .Y(n1094), .A(A[4]) );
  inv04 U1189 ( .Y(n1095), .A(carry_4_) );
  nor02 U1190 ( .Y(n1096), .A0(n1093), .A1(n1097) );
  nor02 U1191 ( .Y(n1098), .A0(n1094), .A1(n1099) );
  nor02 U1192 ( .Y(n1100), .A0(n1095), .A1(n1101) );
  nor02 U1193 ( .Y(n1102), .A0(n1095), .A1(n1103) );
  nor02 U1194 ( .Y(n1091), .A0(n1104), .A1(n1105) );
  nor02 U1195 ( .Y(n1106), .A0(n1094), .A1(n1095) );
  nor02 U1196 ( .Y(n1107), .A0(n1093), .A1(n1095) );
  nor02 U1197 ( .Y(n1108), .A0(n1093), .A1(n1094) );
  nor02 U1198 ( .Y(n1092), .A0(n1108), .A1(n1109) );
  nor02 U1199 ( .Y(n1110), .A0(A[4]), .A1(carry_4_) );
  inv01 U1200 ( .Y(n1097), .A(n1110) );
  nor02 U1201 ( .Y(n1111), .A0(B[4]), .A1(carry_4_) );
  inv01 U1202 ( .Y(n1099), .A(n1111) );
  nor02 U1203 ( .Y(n1112), .A0(B[4]), .A1(A[4]) );
  inv01 U1204 ( .Y(n1101), .A(n1112) );
  nor02 U1205 ( .Y(n1113), .A0(n1093), .A1(n1094) );
  inv01 U1206 ( .Y(n1103), .A(n1113) );
  nor02 U1207 ( .Y(n1114), .A0(n1096), .A1(n1098) );
  inv02 U1208 ( .Y(n1104), .A(n1114) );
  nor02 U1209 ( .Y(n1115), .A0(n1100), .A1(n1102) );
  inv02 U1210 ( .Y(n1105), .A(n1115) );
  nor02 U1211 ( .Y(n1116), .A0(n1106), .A1(n1107) );
  inv01 U1212 ( .Y(n1109), .A(n1116) );
  inv02 U1213 ( .Y(carry_14_), .A(n1118) );
  inv02 U1214 ( .Y(n1119), .A(B[13]) );
  inv02 U1215 ( .Y(n1120), .A(A[13]) );
  inv04 U1216 ( .Y(n1121), .A(carry_13_) );
  nor02 U1217 ( .Y(n1122), .A0(n1119), .A1(n1123) );
  nor02 U1218 ( .Y(n1124), .A0(n1120), .A1(n1125) );
  nor02 U1219 ( .Y(n1126), .A0(n1121), .A1(n1127) );
  nor02 U1220 ( .Y(n1128), .A0(n1121), .A1(n1129) );
  nor02 U1221 ( .Y(n1117), .A0(n1130), .A1(n1131) );
  nor02 U1222 ( .Y(n1132), .A0(n1120), .A1(n1121) );
  nor02 U1223 ( .Y(n1133), .A0(n1119), .A1(n1121) );
  nor02 U1224 ( .Y(n1134), .A0(n1119), .A1(n1120) );
  nor02 U1225 ( .Y(n1118), .A0(n1134), .A1(n1135) );
  nor02 U1226 ( .Y(n1136), .A0(A[13]), .A1(carry_13_) );
  inv01 U1227 ( .Y(n1123), .A(n1136) );
  nor02 U1228 ( .Y(n1137), .A0(B[13]), .A1(carry_13_) );
  inv01 U1229 ( .Y(n1125), .A(n1137) );
  nor02 U1230 ( .Y(n1138), .A0(B[13]), .A1(A[13]) );
  inv01 U1231 ( .Y(n1127), .A(n1138) );
  nor02 U1232 ( .Y(n1139), .A0(n1119), .A1(n1120) );
  inv01 U1233 ( .Y(n1129), .A(n1139) );
  nor02 U1234 ( .Y(n1140), .A0(n1122), .A1(n1124) );
  inv02 U1235 ( .Y(n1130), .A(n1140) );
  nor02 U1236 ( .Y(n1141), .A0(n1126), .A1(n1128) );
  inv02 U1237 ( .Y(n1131), .A(n1141) );
  nor02 U1238 ( .Y(n1142), .A0(n1132), .A1(n1133) );
  inv01 U1239 ( .Y(n1135), .A(n1142) );
  inv02 U1240 ( .Y(carry_19_), .A(n1144) );
  inv02 U1241 ( .Y(n1145), .A(B[18]) );
  inv02 U1242 ( .Y(n1146), .A(A[18]) );
  inv04 U1243 ( .Y(n1147), .A(carry_18_) );
  nor02 U1244 ( .Y(n1148), .A0(n1145), .A1(n1149) );
  nor02 U1245 ( .Y(n1150), .A0(n1146), .A1(n1151) );
  nor02 U1246 ( .Y(n1152), .A0(n1147), .A1(n1153) );
  nor02 U1247 ( .Y(n1154), .A0(n1147), .A1(n1155) );
  nor02 U1248 ( .Y(n1143), .A0(n1156), .A1(n1157) );
  nor02 U1249 ( .Y(n1158), .A0(n1146), .A1(n1147) );
  nor02 U1250 ( .Y(n1159), .A0(n1145), .A1(n1147) );
  nor02 U1251 ( .Y(n1160), .A0(n1145), .A1(n1146) );
  nor02 U1252 ( .Y(n1144), .A0(n1160), .A1(n1161) );
  nor02 U1253 ( .Y(n1162), .A0(A[18]), .A1(carry_18_) );
  inv01 U1254 ( .Y(n1149), .A(n1162) );
  nor02 U1255 ( .Y(n1163), .A0(B[18]), .A1(carry_18_) );
  inv01 U1256 ( .Y(n1151), .A(n1163) );
  nor02 U1257 ( .Y(n1164), .A0(B[18]), .A1(A[18]) );
  inv01 U1258 ( .Y(n1153), .A(n1164) );
  nor02 U1259 ( .Y(n1165), .A0(n1145), .A1(n1146) );
  inv01 U1260 ( .Y(n1155), .A(n1165) );
  nor02 U1261 ( .Y(n1166), .A0(n1148), .A1(n1150) );
  inv02 U1262 ( .Y(n1156), .A(n1166) );
  nor02 U1263 ( .Y(n1167), .A0(n1152), .A1(n1154) );
  inv02 U1264 ( .Y(n1157), .A(n1167) );
  nor02 U1265 ( .Y(n1168), .A0(n1158), .A1(n1159) );
  inv01 U1266 ( .Y(n1161), .A(n1168) );
  inv02 U1267 ( .Y(carry_15_), .A(n1170) );
  inv02 U1268 ( .Y(n1171), .A(B[14]) );
  inv02 U1269 ( .Y(n1172), .A(A[14]) );
  inv04 U1270 ( .Y(n1173), .A(carry_14_) );
  nor02 U1271 ( .Y(n1174), .A0(n1171), .A1(n1175) );
  nor02 U1272 ( .Y(n1176), .A0(n1172), .A1(n1177) );
  nor02 U1273 ( .Y(n1178), .A0(n1173), .A1(n1179) );
  nor02 U1274 ( .Y(n1180), .A0(n1173), .A1(n1181) );
  nor02 U1275 ( .Y(n1169), .A0(n1182), .A1(n1183) );
  nor02 U1276 ( .Y(n1184), .A0(n1172), .A1(n1173) );
  nor02 U1277 ( .Y(n1185), .A0(n1171), .A1(n1173) );
  nor02 U1278 ( .Y(n1186), .A0(n1171), .A1(n1172) );
  nor02 U1279 ( .Y(n1170), .A0(n1186), .A1(n1187) );
  nor02 U1280 ( .Y(n1188), .A0(A[14]), .A1(carry_14_) );
  inv01 U1281 ( .Y(n1175), .A(n1188) );
  nor02 U1282 ( .Y(n1189), .A0(B[14]), .A1(carry_14_) );
  inv01 U1283 ( .Y(n1177), .A(n1189) );
  nor02 U1284 ( .Y(n1190), .A0(B[14]), .A1(A[14]) );
  inv01 U1285 ( .Y(n1179), .A(n1190) );
  nor02 U1286 ( .Y(n1191), .A0(n1171), .A1(n1172) );
  inv01 U1287 ( .Y(n1181), .A(n1191) );
  nor02 U1288 ( .Y(n1192), .A0(n1174), .A1(n1176) );
  inv02 U1289 ( .Y(n1182), .A(n1192) );
  nor02 U1290 ( .Y(n1193), .A0(n1178), .A1(n1180) );
  inv02 U1291 ( .Y(n1183), .A(n1193) );
  nor02 U1292 ( .Y(n1194), .A0(n1184), .A1(n1185) );
  inv01 U1293 ( .Y(n1187), .A(n1194) );
  inv02 U1294 ( .Y(carry_3_), .A(n1196) );
  inv02 U1295 ( .Y(n1197), .A(B[2]) );
  inv02 U1296 ( .Y(n1198), .A(A[2]) );
  inv04 U1297 ( .Y(n1199), .A(carry_2_) );
  nor02 U1298 ( .Y(n1200), .A0(n1197), .A1(n1201) );
  nor02 U1299 ( .Y(n1202), .A0(n1198), .A1(n1203) );
  nor02 U1300 ( .Y(n1204), .A0(n1199), .A1(n1205) );
  nor02 U1301 ( .Y(n1206), .A0(n1199), .A1(n1207) );
  nor02 U1302 ( .Y(n1195), .A0(n1208), .A1(n1209) );
  nor02 U1303 ( .Y(n1210), .A0(n1198), .A1(n1199) );
  nor02 U1304 ( .Y(n1211), .A0(n1197), .A1(n1199) );
  nor02 U1305 ( .Y(n1212), .A0(n1197), .A1(n1198) );
  nor02 U1306 ( .Y(n1196), .A0(n1212), .A1(n1213) );
  nor02 U1307 ( .Y(n1214), .A0(A[2]), .A1(carry_2_) );
  inv01 U1308 ( .Y(n1201), .A(n1214) );
  nor02 U1309 ( .Y(n1215), .A0(B[2]), .A1(carry_2_) );
  inv01 U1310 ( .Y(n1203), .A(n1215) );
  nor02 U1311 ( .Y(n1216), .A0(B[2]), .A1(A[2]) );
  inv01 U1312 ( .Y(n1205), .A(n1216) );
  nor02 U1313 ( .Y(n1217), .A0(n1197), .A1(n1198) );
  inv01 U1314 ( .Y(n1207), .A(n1217) );
  nor02 U1315 ( .Y(n1218), .A0(n1200), .A1(n1202) );
  inv02 U1316 ( .Y(n1208), .A(n1218) );
  nor02 U1317 ( .Y(n1219), .A0(n1204), .A1(n1206) );
  inv02 U1318 ( .Y(n1209), .A(n1219) );
  nor02 U1319 ( .Y(n1220), .A0(n1210), .A1(n1211) );
  inv01 U1320 ( .Y(n1213), .A(n1220) );
  inv02 U1321 ( .Y(carry_4_), .A(n1222) );
  inv02 U1322 ( .Y(n1223), .A(B[3]) );
  inv02 U1323 ( .Y(n1224), .A(A[3]) );
  inv04 U1324 ( .Y(n1225), .A(carry_3_) );
  nor02 U1325 ( .Y(n1226), .A0(n1223), .A1(n1227) );
  nor02 U1326 ( .Y(n1228), .A0(n1224), .A1(n1229) );
  nor02 U1327 ( .Y(n1230), .A0(n1225), .A1(n1231) );
  nor02 U1328 ( .Y(n1232), .A0(n1225), .A1(n1233) );
  nor02 U1329 ( .Y(n1221), .A0(n1234), .A1(n1235) );
  nor02 U1330 ( .Y(n1236), .A0(n1224), .A1(n1225) );
  nor02 U1331 ( .Y(n1237), .A0(n1223), .A1(n1225) );
  nor02 U1332 ( .Y(n1238), .A0(n1223), .A1(n1224) );
  nor02 U1333 ( .Y(n1222), .A0(n1238), .A1(n1239) );
  nor02 U1334 ( .Y(n1240), .A0(A[3]), .A1(carry_3_) );
  inv01 U1335 ( .Y(n1227), .A(n1240) );
  nor02 U1336 ( .Y(n1241), .A0(B[3]), .A1(carry_3_) );
  inv01 U1337 ( .Y(n1229), .A(n1241) );
  nor02 U1338 ( .Y(n1242), .A0(B[3]), .A1(A[3]) );
  inv01 U1339 ( .Y(n1231), .A(n1242) );
  nor02 U1340 ( .Y(n1243), .A0(n1223), .A1(n1224) );
  inv01 U1341 ( .Y(n1233), .A(n1243) );
  nor02 U1342 ( .Y(n1244), .A0(n1226), .A1(n1228) );
  inv02 U1343 ( .Y(n1234), .A(n1244) );
  nor02 U1344 ( .Y(n1245), .A0(n1230), .A1(n1232) );
  inv02 U1345 ( .Y(n1235), .A(n1245) );
  nor02 U1346 ( .Y(n1246), .A0(n1236), .A1(n1237) );
  inv01 U1347 ( .Y(n1239), .A(n1246) );
  inv02 U1348 ( .Y(carry_13_), .A(n1248) );
  inv02 U1349 ( .Y(n1249), .A(B[12]) );
  inv02 U1350 ( .Y(n1250), .A(A[12]) );
  inv02 U1351 ( .Y(n1251), .A(carry_12_) );
  nor02 U1352 ( .Y(n1252), .A0(n1249), .A1(n1253) );
  nor02 U1353 ( .Y(n1254), .A0(n1250), .A1(n1255) );
  nor02 U1354 ( .Y(n1256), .A0(n1251), .A1(n1257) );
  nor02 U1355 ( .Y(n1258), .A0(n1251), .A1(n1259) );
  nor02 U1356 ( .Y(n1247), .A0(n1260), .A1(n1261) );
  nor02 U1357 ( .Y(n1262), .A0(n1250), .A1(n1251) );
  nor02 U1358 ( .Y(n1263), .A0(n1249), .A1(n1251) );
  nor02 U1359 ( .Y(n1264), .A0(n1249), .A1(n1250) );
  nor02 U1360 ( .Y(n1248), .A0(n1264), .A1(n1265) );
  nor02 U1361 ( .Y(n1266), .A0(A[12]), .A1(carry_12_) );
  inv01 U1362 ( .Y(n1253), .A(n1266) );
  nor02 U1363 ( .Y(n1267), .A0(B[12]), .A1(carry_12_) );
  inv01 U1364 ( .Y(n1255), .A(n1267) );
  nor02 U1365 ( .Y(n1268), .A0(B[12]), .A1(A[12]) );
  inv01 U1366 ( .Y(n1257), .A(n1268) );
  nor02 U1367 ( .Y(n1269), .A0(n1249), .A1(n1250) );
  inv01 U1368 ( .Y(n1259), .A(n1269) );
  nor02 U1369 ( .Y(n1270), .A0(n1252), .A1(n1254) );
  inv02 U1370 ( .Y(n1260), .A(n1270) );
  nor02 U1371 ( .Y(n1271), .A0(n1256), .A1(n1258) );
  inv02 U1372 ( .Y(n1261), .A(n1271) );
  nor02 U1373 ( .Y(n1272), .A0(n1262), .A1(n1263) );
  inv01 U1374 ( .Y(n1265), .A(n1272) );
  inv02 U1375 ( .Y(carry_18_), .A(n1274) );
  inv02 U1376 ( .Y(n1275), .A(B[17]) );
  inv02 U1377 ( .Y(n1276), .A(A[17]) );
  inv02 U1378 ( .Y(n1277), .A(carry_17_) );
  nor02 U1379 ( .Y(n1278), .A0(n1275), .A1(n1279) );
  nor02 U1380 ( .Y(n1280), .A0(n1276), .A1(n1281) );
  nor02 U1381 ( .Y(n1282), .A0(n1277), .A1(n1283) );
  nor02 U1382 ( .Y(n1284), .A0(n1277), .A1(n1285) );
  nor02 U1383 ( .Y(n1273), .A0(n1286), .A1(n1287) );
  nor02 U1384 ( .Y(n1288), .A0(n1276), .A1(n1277) );
  nor02 U1385 ( .Y(n1289), .A0(n1275), .A1(n1277) );
  nor02 U1386 ( .Y(n1290), .A0(n1275), .A1(n1276) );
  nor02 U1387 ( .Y(n1274), .A0(n1290), .A1(n1291) );
  nor02 U1388 ( .Y(n1292), .A0(A[17]), .A1(carry_17_) );
  inv01 U1389 ( .Y(n1279), .A(n1292) );
  nor02 U1390 ( .Y(n1293), .A0(B[17]), .A1(carry_17_) );
  inv01 U1391 ( .Y(n1281), .A(n1293) );
  nor02 U1392 ( .Y(n1294), .A0(B[17]), .A1(A[17]) );
  inv01 U1393 ( .Y(n1283), .A(n1294) );
  nor02 U1394 ( .Y(n1295), .A0(n1275), .A1(n1276) );
  inv01 U1395 ( .Y(n1285), .A(n1295) );
  nor02 U1396 ( .Y(n1296), .A0(n1278), .A1(n1280) );
  inv02 U1397 ( .Y(n1286), .A(n1296) );
  nor02 U1398 ( .Y(n1297), .A0(n1282), .A1(n1284) );
  inv02 U1399 ( .Y(n1287), .A(n1297) );
  nor02 U1400 ( .Y(n1298), .A0(n1288), .A1(n1289) );
  inv01 U1401 ( .Y(n1291), .A(n1298) );
  inv02 U1402 ( .Y(carry_2_), .A(n1300) );
  inv02 U1403 ( .Y(n1301), .A(B[1]) );
  inv02 U1404 ( .Y(n1302), .A(A[1]) );
  inv02 U1405 ( .Y(n1303), .A(n4) );
  nor02 U1406 ( .Y(n1304), .A0(n1301), .A1(n1305) );
  nor02 U1407 ( .Y(n1306), .A0(n1302), .A1(n1307) );
  nor02 U1408 ( .Y(n1308), .A0(n1303), .A1(n1309) );
  nor02 U1409 ( .Y(n1310), .A0(n1303), .A1(n1311) );
  nor02 U1410 ( .Y(n1299), .A0(n1312), .A1(n1313) );
  nor02 U1411 ( .Y(n1314), .A0(n1302), .A1(n1303) );
  nor02 U1412 ( .Y(n1315), .A0(n1301), .A1(n1303) );
  nor02 U1413 ( .Y(n1316), .A0(n1301), .A1(n1302) );
  nor02 U1414 ( .Y(n1300), .A0(n1316), .A1(n1317) );
  nor02 U1415 ( .Y(n1318), .A0(A[1]), .A1(n4) );
  inv01 U1416 ( .Y(n1305), .A(n1318) );
  nor02 U1417 ( .Y(n1319), .A0(B[1]), .A1(n4) );
  inv01 U1418 ( .Y(n1307), .A(n1319) );
  nor02 U1419 ( .Y(n1320), .A0(B[1]), .A1(A[1]) );
  inv01 U1420 ( .Y(n1309), .A(n1320) );
  nor02 U1421 ( .Y(n1321), .A0(n1301), .A1(n1302) );
  inv01 U1422 ( .Y(n1311), .A(n1321) );
  nor02 U1423 ( .Y(n1322), .A0(n1304), .A1(n1306) );
  inv02 U1424 ( .Y(n1312), .A(n1322) );
  nor02 U1425 ( .Y(n1323), .A0(n1308), .A1(n1310) );
  inv02 U1426 ( .Y(n1313), .A(n1323) );
  nor02 U1427 ( .Y(n1324), .A0(n1314), .A1(n1315) );
  inv01 U1428 ( .Y(n1317), .A(n1324) );
  xor2 U1429 ( .Y(n1325), .A0(B[0]), .A1(A[0]) );
endmodule


module sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_dec_5_1 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   carry_4_, carry_3_, n5, n7, n9, n11, n13, n14, n15;

  xor2 U6 ( .Y(n5), .A0(A[1]), .A1(A[0]) );
  inv01 U7 ( .Y(SUM[1]), .A(n5) );
  xor2 U8 ( .Y(n7), .A0(A[3]), .A1(n15) );
  inv01 U9 ( .Y(SUM[3]), .A(n7) );
  xor2 U10 ( .Y(n9), .A0(carry_4_), .A1(A[4]) );
  inv01 U11 ( .Y(SUM[4]), .A(n9) );
  xor2 U12 ( .Y(n11), .A0(A[2]), .A1(n14) );
  inv01 U13 ( .Y(SUM[2]), .A(n11) );
  nor02 U14 ( .Y(n13), .A0(A[1]), .A1(A[0]) );
  inv02 U15 ( .Y(n14), .A(n13) );
  buf02 U16 ( .Y(n15), .A(carry_3_) );
  inv01 U17 ( .Y(SUM[0]), .A(A[0]) );
  or02 U1_B_2 ( .Y(carry_3_), .A0(A[2]), .A1(n14) );
  or02 U1_B_3 ( .Y(carry_4_), .A0(A[3]), .A1(n15) );
endmodule


module sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_dec_5_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   carry_4_, carry_3_, carry_2_, n5, n7, n9, n11, n13, n14;

  xor2 U6 ( .Y(n5), .A0(carry_4_), .A1(A[4]) );
  inv01 U7 ( .Y(SUM[4]), .A(n5) );
  xor2 U8 ( .Y(n7), .A0(A[2]), .A1(n13) );
  inv01 U9 ( .Y(SUM[2]), .A(n7) );
  xor2 U10 ( .Y(n9), .A0(A[1]), .A1(A[0]) );
  inv01 U11 ( .Y(SUM[1]), .A(n9) );
  xor2 U12 ( .Y(n11), .A0(A[3]), .A1(n14) );
  inv01 U13 ( .Y(SUM[3]), .A(n11) );
  buf02 U14 ( .Y(n13), .A(carry_2_) );
  buf02 U15 ( .Y(n14), .A(carry_3_) );
  inv01 U16 ( .Y(SUM[0]), .A(A[0]) );
  or02 U1_B_1 ( .Y(carry_2_), .A0(A[1]), .A1(A[0]) );
  or02 U1_B_2 ( .Y(carry_3_), .A0(A[2]), .A1(n13) );
  or02 U1_B_3 ( .Y(carry_4_), .A0(A[3]), .A1(n14) );
endmodule


module sqrt_RD_WIDTH52_SQ_WIDTH26 ( clk_i, rad_i, start_i, ready_o, sqr_o, 
        ine_o );
  input [51:0] rad_i;
  output [25:0] sqr_o;
  input clk_i, start_i;
  output ready_o, ine_o;
  wire   s_sqr_o_25_, s_sqr_o_24_, s_sqr_o_23_, s_sqr_o_22_, s_sqr_o_21_,
         s_sqr_o_20_, s_sqr_o_19_, s_sqr_o_18_, s_sqr_o_17_, s_sqr_o_16_,
         s_sqr_o_15_, s_sqr_o_14_, s_sqr_o_13_, s_sqr_o_12_, s_sqr_o_11_,
         s_sqr_o_10_, s_sqr_o_9_, s_sqr_o_8_, s_sqr_o_7_, s_sqr_o_6_,
         s_sqr_o_5_, s_sqr_o_4_, s_sqr_o_3_, s_sqr_o_2_, s_sqr_o_1_,
         s_sqr_o_0_, s_ine_o, s_ready_o, b_25_, b_24_, b_23_, b_22_, b_21_,
         b_20_, b_19_, b_18_, b_17_, b_16_, b_15_, b_14_, b_13_, b_12_, b_11_,
         b_10_, b_9_, b_8_, b_7_, b_6_, b_5_, b_4_, b_3_, b_2_, b_1_, b_0_,
         s_sum2a_25_, s_sum2a_24_, s_sum2a_23_, s_sum2a_22_, s_sum2a_21_,
         s_sum2a_20_, s_sum2a_19_, s_sum2a_18_, s_sum2a_17_, s_sum2a_16_,
         s_sum2a_15_, s_sum2a_14_, s_sum2a_13_, s_sum2a_12_, s_sum2a_11_,
         s_sum2a_10_, s_sum2a_9_, s_sum2a_8_, s_sum2a_7_, s_sum2a_6_,
         s_sum2a_5_, s_sum2a_4_, s_sum2a_3_, s_sum2a_2_, s_sum2a_1_,
         s_sum2a_0_, s_sum1a_25_, s_sum1a_24_, s_sum1a_23_, s_sum1a_22_,
         s_sum1a_21_, s_sum1a_20_, s_sum1a_19_, s_sum1a_18_, s_sum1a_17_,
         s_sum1a_16_, s_sum1a_15_, s_sum1a_14_, s_sum1a_13_, s_sum1a_12_,
         s_sum1a_11_, s_sum1a_10_, s_sum1a_9_, s_sum1a_8_, s_sum1a_7_,
         s_sum1a_6_, s_sum1a_5_, s_sum1a_4_, s_sum1a_3_, s_sum1a_2_,
         s_sum1a_1_, s_sum1a_0_, r1_50_, r1_49_, r1_48_, r1_47_, r1_46_,
         r1_45_, r1_44_, r1_43_, r1_42_, r1_41_, r1_40_, r1_39_, r1_38_,
         r1_37_, r1_36_, r1_35_, r1_34_, r1_33_, r1_32_, r1_31_, r1_30_,
         r1_29_, r1_28_, r1_27_, r1_26_, r1_25_, r1_24_, r1_23_, r1_22_,
         r1_21_, r1_20_, r1_19_, r1_18_, r1_17_, r1_16_, r1_15_, r1_14_,
         r1_13_, r1_12_, r1_11_, r1_10_, r1_9_, r1_8_, r1_7_, r1_6_, r1_5_,
         r1_4_, r1_3_, r1_2_, r1_1_, r1_0_, s_rad_i_51_, s_rad_i_50_,
         s_rad_i_49_, s_rad_i_48_, s_rad_i_47_, s_rad_i_46_, s_rad_i_45_,
         s_rad_i_44_, s_rad_i_43_, s_rad_i_42_, s_rad_i_41_, s_rad_i_40_,
         s_rad_i_39_, s_rad_i_38_, s_rad_i_37_, s_rad_i_36_, s_rad_i_35_,
         s_rad_i_34_, s_rad_i_33_, s_rad_i_32_, s_rad_i_31_, s_rad_i_30_,
         s_rad_i_29_, s_rad_i_28_, s_rad_i_27_, s_rad_i_26_, s_rad_i_25_,
         s_rad_i_24_, s_rad_i_23_, s_rad_i_22_, s_rad_i_21_, s_rad_i_20_,
         s_rad_i_19_, s_rad_i_18_, s_rad_i_17_, s_rad_i_16_, s_rad_i_15_,
         s_rad_i_14_, s_rad_i_13_, s_rad_i_12_, s_rad_i_11_, s_rad_i_10_,
         s_rad_i_9_, s_rad_i_8_, s_rad_i_7_, s_rad_i_6_, s_rad_i_5_,
         s_rad_i_4_, s_rad_i_3_, s_rad_i_2_, s_rad_i_1_, s_rad_i_0_, s_state,
         s_state110, s_count_4_, s_count_3_, s_count_2_, s_count_1_,
         s_count_0_, sum181_4_, sum181_3_, sum181_2_, sum181_1_, sum181_0_,
         b206_25_, c222_4_, c222_3_, c222_2_, c222_1_, c222_0_, c_4_, c_3_,
         c_2_, c_1_, c_0_, ARG260_4_, ARG260_3_, ARG260_2_, ARG260_1_,
         ARG260_0_, s_op1_51_, s_op1_50_, s_op1_49_, s_op1_48_, s_op1_47_,
         s_op1_46_, s_op1_45_, s_op1_44_, s_op1_43_, s_op1_42_, s_op1_41_,
         s_op1_40_, s_op1_39_, s_op1_38_, s_op1_37_, s_op1_36_, s_op1_35_,
         s_op1_34_, s_op1_33_, s_op1_32_, s_op1_31_, s_op1_30_, s_op1_29_,
         s_op1_28_, s_op1_27_, s_op1_26_, s_op1_25_, s_op1_24_, s_op1_23_,
         s_op1_22_, s_op1_21_, s_op1_20_, s_op1_19_, s_op1_18_, s_op1_17_,
         s_op1_16_, s_op1_15_, s_op1_14_, s_op1_13_, s_op1_12_, s_op1_11_,
         s_op1_10_, s_op1_9_, s_op1_8_, s_op1_7_, s_op1_6_, s_op1_5_, s_op1_4_,
         s_op1_3_, s_op1_2_, s_op1_1_, s_op1_0_, r0_2_51_, r0_2_50_, r0_2_49_,
         r0_2_48_, r0_2_47_, r0_2_46_, r0_2_45_, r0_2_44_, r0_2_43_, r0_2_42_,
         r0_2_41_, r0_2_40_, r0_2_39_, r0_2_38_, r0_2_37_, r0_2_36_, r0_2_35_,
         r0_2_34_, r0_2_33_, r0_2_32_, r0_2_31_, r0_2_30_, r0_2_29_, r0_2_28_,
         r0_2_27_, r0_2_26_, r0_2_25_, r0_2_24_, r0_2_23_, r0_2_22_, r0_2_21_,
         r0_2_20_, r0_2_19_, r0_2_18_, r0_2_17_, r0_2_16_, r0_2_15_, r0_2_14_,
         r0_2_13_, r0_2_12_, r0_2_11_, r0_2_10_, r0_2_9_, r0_2_8_, r0_2_7_,
         r0_2_6_, r0_2_5_, r0_2_4_, r0_2_3_, r0_2_2_, r0_2_1_, r0_2_0_,
         result407_50_, s_op2_51_, s_op2_49_, s_op2_48_, s_op2_47_, s_op2_46_,
         s_op2_45_, s_op2_44_, s_op2_43_, s_op2_42_, s_op2_41_, s_op2_40_,
         s_op2_39_, s_op2_38_, s_op2_37_, s_op2_36_, s_op2_23_, s_op2_22_,
         s_op2_21_, s_op2_19_, s_op2_18_, s_op2_17_, s_op2_16_, s_op2_7_,
         s_op2_6_, s_op2_5_, s_op2_4_, s_op2_3_, r0_51_, r0_50_, r0_49_,
         r0_48_, r0_47_, r0_46_, r0_45_, r0_44_, r0_43_, r0_42_, r0_41_,
         r0_40_, r0_39_, r0_38_, r0_37_, r0_36_, r0_35_, r0_34_, r0_33_,
         r0_32_, r0_31_, r0_30_, r0_29_, r0_28_, r0_27_, r0_26_, r0_25_,
         r0_24_, r0_23_, r0_22_, r0_21_, r0_20_, r0_19_, r0_18_, r0_17_,
         r0_16_, r0_15_, r0_14_, r0_13_, r0_12_, r0_11_, r0_10_, r0_9_, r0_8_,
         r0_7_, r0_6_, r0_5_, r0_4_, r0_3_, r0_2_, r0_1_, r0_0_,
         n____return912, r1_2_51_, r1_2_50_, r1_2_49_, r1_2_48_, r1_2_47_,
         r1_2_46_, r1_2_45_, r1_2_44_, r1_2_43_, r1_2_42_, r1_2_41_, r1_2_40_,
         r1_2_39_, r1_2_38_, r1_2_37_, r1_2_36_, r1_2_35_, r1_2_34_, r1_2_33_,
         r1_2_32_, r1_2_31_, r1_2_30_, r1_2_29_, r1_2_28_, r1_2_27_, r1_2_26_,
         r1_2_25_, r1_2_24_, r1_2_23_, r1_2_22_, r1_2_21_, r1_2_20_, r1_2_19_,
         r1_2_18_, r1_2_17_, r1_2_16_, r1_2_15_, r1_2_14_, r1_2_13_, r1_2_12_,
         r1_2_11_, r1_2_10_, r1_2_9_, r1_2_8_, r1_2_7_, r1_2_6_, r1_2_5_,
         r1_2_4_, r1_2_3_, r1_2_2_, r1_2_1_, r1_2_0_, n____return1071,
         ARG1118_25_, ARG1118_24_, ARG1118_23_, ARG1118_22_, ARG1118_21_,
         ARG1118_20_, ARG1118_19_, ARG1118_18_, ARG1118_17_, ARG1118_16_,
         ARG1118_15_, ARG1118_14_, ARG1118_13_, ARG1118_12_, ARG1118_11_,
         ARG1118_10_, ARG1118_9_, ARG1118_8_, ARG1118_7_, ARG1118_6_,
         ARG1118_5_, ARG1118_4_, ARG1118_3_, ARG1118_2_, ARG1118_1_,
         ARG1118_0_, n1384_51_, n1384_49_, n____return1382_50_,
         n____return1382_48_, n____return1382_47_, n____return1382_46_,
         n____return1382_45_, n____return1382_44_, n____return1382_43_,
         n____return1382_42_, n____return1382_41_, n____return1382_40_,
         n____return1382_39_, n____return1382_38_, n____return1382_37_,
         n____return1382_36_, n____return1382_35_, n____return1382_34_,
         n____return1382_33_, n____return1382_32_, n____return1382_31_,
         n____return1382_30_, n____return1382_29_, n____return1382_28_,
         n____return1382_27_, n____return1382_26_, n____return1382_25_,
         n____return1382_24_, n____return1382_23_, n____return1382_22_,
         n____return1382_21_, n____return1382_20_, n____return1382_19_,
         n____return1382_18_, n____return1382_17_, n____return1382_16_,
         n____return1382_15_, n____return1382_14_, n____return1382_13_,
         n____return1382_12_, n____return1382_11_, n____return1382_10_,
         n____return1382_9_, n____return1382_8_, n____return1382_7_,
         n____return1382_6_, n____return1382_5_, n____return1382_4_,
         n____return1382_3_, n____return1382_2_, n____return1382_1_,
         n____return1382_0_, n1346_49_, n____return1344_51_,
         n____return1344_50_, n____return1344_48_, n____return1344_47_,
         n____return1344_46_, n____return1344_45_, n____return1344_44_,
         n____return1344_43_, n____return1344_42_, n____return1344_41_,
         n____return1344_40_, n____return1344_39_, n____return1344_38_,
         n____return1344_37_, n____return1344_36_, n____return1344_35_,
         n____return1344_34_, n____return1344_33_, n____return1344_32_,
         n____return1344_31_, n____return1344_30_, n____return1344_29_,
         n____return1344_28_, n____return1344_27_, n____return1344_26_,
         n____return1344_25_, n____return1344_24_, n____return1344_23_,
         n____return1344_22_, n____return1344_21_, n____return1344_20_,
         n____return1344_19_, n____return1344_18_, n____return1344_17_,
         n____return1344_16_, n____return1344_15_, n____return1344_14_,
         n____return1344_13_, n____return1344_12_, n____return1344_11_,
         n____return1344_10_, n____return1344_9_, n____return1344_8_,
         n____return1344_7_, n____return1344_6_, n____return1344_5_,
         n____return1344_4_, n____return1344_3_, n____return1344_2_,
         n____return1344_1_, n____return1344_0_, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007;
  wire   [51:0] b_2;
  wire   [51:0] s_sum2b;
  wire   [51:0] s_sum1b;

  dff s_count_reg_0_ ( .Q(s_count_0_), .D(n2837), .CLK(clk_i) );
  dff s_count_reg_1_ ( .Q(s_count_1_), .D(n2838), .CLK(clk_i) );
  dff s_count_reg_2_ ( .Q(s_count_2_), .D(n2839), .CLK(clk_i) );
  dff s_count_reg_3_ ( .Q(s_count_3_), .D(n2840), .CLK(clk_i) );
  dff s_count_reg_4_ ( .Q(s_count_4_), .D(n2841), .CLK(clk_i) );
  dff r0_reg_51_ ( .Q(r0_51_), .D(n2842), .CLK(clk_i) );
  dff r0_reg_50_ ( .Q(r0_50_), .D(n2843), .CLK(clk_i) );
  dff r0_reg_49_ ( .Q(r0_49_), .D(n3411), .CLK(clk_i) );
  dff r0_reg_48_ ( .Q(r0_48_), .D(n3087), .CLK(clk_i) );
  dff r0_reg_47_ ( .Q(r0_47_), .D(n3123), .CLK(clk_i) );
  dff r0_reg_46_ ( .Q(r0_46_), .D(n3139), .CLK(clk_i) );
  dff r0_reg_45_ ( .Q(r0_45_), .D(n3147), .CLK(clk_i) );
  dff r0_reg_44_ ( .Q(r0_44_), .D(n3165), .CLK(clk_i) );
  dff r0_reg_43_ ( .Q(r0_43_), .D(n3143), .CLK(clk_i) );
  dff r0_reg_42_ ( .Q(r0_42_), .D(n3097), .CLK(clk_i) );
  dff r0_reg_41_ ( .Q(r0_41_), .D(n3093), .CLK(clk_i) );
  dff r0_reg_40_ ( .Q(r0_40_), .D(n3131), .CLK(clk_i) );
  dff r0_reg_39_ ( .Q(r0_39_), .D(n3163), .CLK(clk_i) );
  dff r0_reg_38_ ( .Q(r0_38_), .D(n3169), .CLK(clk_i) );
  dff r0_reg_37_ ( .Q(r0_37_), .D(n3129), .CLK(clk_i) );
  dff r0_reg_36_ ( .Q(r0_36_), .D(n3105), .CLK(clk_i) );
  dff r0_reg_35_ ( .Q(r0_35_), .D(n3091), .CLK(clk_i) );
  dff r0_reg_34_ ( .Q(r0_34_), .D(n3167), .CLK(clk_i) );
  dff r0_reg_33_ ( .Q(r0_33_), .D(n3095), .CLK(clk_i) );
  dff r0_reg_32_ ( .Q(r0_32_), .D(n3135), .CLK(clk_i) );
  dff r0_reg_31_ ( .Q(r0_31_), .D(n3141), .CLK(clk_i) );
  dff r0_reg_30_ ( .Q(r0_30_), .D(n3133), .CLK(clk_i) );
  dff r0_reg_29_ ( .Q(r0_29_), .D(n3125), .CLK(clk_i) );
  dff r0_reg_28_ ( .Q(r0_28_), .D(n3103), .CLK(clk_i) );
  dff r0_reg_27_ ( .Q(r0_27_), .D(n3137), .CLK(clk_i) );
  dff r0_reg_26_ ( .Q(r0_26_), .D(n3145), .CLK(clk_i) );
  dff r0_reg_25_ ( .Q(r0_25_), .QB(n7144), .D(n2868), .CLK(clk_i) );
  dff r0_reg_24_ ( .Q(r0_24_), .D(n2869), .CLK(clk_i) );
  dff r0_reg_23_ ( .Q(r0_23_), .D(n2870), .CLK(clk_i) );
  dff r0_reg_22_ ( .Q(r0_22_), .D(n2871), .CLK(clk_i) );
  dff r0_reg_21_ ( .Q(r0_21_), .D(n2872), .CLK(clk_i) );
  dff r0_reg_20_ ( .Q(r0_20_), .D(n2873), .CLK(clk_i) );
  dff r0_reg_19_ ( .Q(r0_19_), .D(n2874), .CLK(clk_i) );
  dff r0_reg_18_ ( .Q(r0_18_), .D(n2875), .CLK(clk_i) );
  dff r0_reg_17_ ( .Q(r0_17_), .D(n2876), .CLK(clk_i) );
  dff r0_reg_16_ ( .Q(r0_16_), .D(n2877), .CLK(clk_i) );
  dff r0_reg_15_ ( .Q(r0_15_), .D(n2878), .CLK(clk_i) );
  dff r0_reg_14_ ( .Q(r0_14_), .D(n2879), .CLK(clk_i) );
  dff r0_reg_13_ ( .Q(r0_13_), .D(n2880), .CLK(clk_i) );
  dff r0_reg_12_ ( .Q(r0_12_), .D(n2881), .CLK(clk_i) );
  dff r0_reg_11_ ( .Q(r0_11_), .D(n2882), .CLK(clk_i) );
  dff r0_reg_10_ ( .Q(r0_10_), .D(n2883), .CLK(clk_i) );
  dff r0_reg_9_ ( .Q(r0_9_), .D(n2884), .CLK(clk_i) );
  dff r0_reg_8_ ( .Q(r0_8_), .D(n2885), .CLK(clk_i) );
  dff r0_reg_7_ ( .Q(r0_7_), .D(n2886), .CLK(clk_i) );
  dff r0_reg_6_ ( .Q(r0_6_), .D(n2887), .CLK(clk_i) );
  dff r0_reg_5_ ( .Q(r0_5_), .D(n2888), .CLK(clk_i) );
  dff r0_reg_4_ ( .Q(r0_4_), .QB(n7124), .D(n2889), .CLK(clk_i) );
  dff r0_reg_3_ ( .Q(r0_3_), .D(n2890), .CLK(clk_i) );
  dff r0_reg_2_ ( .Q(r0_2_), .QB(n7120), .D(n2891), .CLK(clk_i) );
  dff r0_reg_1_ ( .Q(r0_1_), .D(n2892), .CLK(clk_i) );
  dff r0_reg_0_ ( .Q(r0_0_), .D(n2893), .CLK(clk_i) );
  dff r0_2_reg_51_ ( .Q(r0_2_51_), .QB(n2778), .D(n2894), .CLK(clk_i) );
  dff r0_2_reg_50_ ( .Q(r0_2_50_), .QB(n2777), .D(n2895), .CLK(clk_i) );
  dff r0_2_reg_49_ ( .Q(r0_2_49_), .QB(n2775), .D(n2896), .CLK(clk_i) );
  dff r0_2_reg_48_ ( .Q(r0_2_48_), .QB(n2774), .D(n2897), .CLK(clk_i) );
  dff r0_2_reg_47_ ( .Q(r0_2_47_), .QB(n2773), .D(n2898), .CLK(clk_i) );
  dff r0_2_reg_46_ ( .Q(r0_2_46_), .QB(n2772), .D(n2899), .CLK(clk_i) );
  dff r0_2_reg_45_ ( .Q(r0_2_45_), .QB(n2771), .D(n2900), .CLK(clk_i) );
  dff r0_2_reg_44_ ( .Q(r0_2_44_), .QB(n2770), .D(n2901), .CLK(clk_i) );
  dff r0_2_reg_43_ ( .Q(r0_2_43_), .QB(n2769), .D(n2902), .CLK(clk_i) );
  dff r0_2_reg_42_ ( .Q(r0_2_42_), .QB(n2768), .D(n2903), .CLK(clk_i) );
  dff r0_2_reg_41_ ( .Q(r0_2_41_), .QB(n2767), .D(n2904), .CLK(clk_i) );
  dff r0_2_reg_40_ ( .Q(r0_2_40_), .QB(n2766), .D(n2905), .CLK(clk_i) );
  dff r0_2_reg_39_ ( .Q(r0_2_39_), .QB(n2764), .D(n2906), .CLK(clk_i) );
  dff r0_2_reg_38_ ( .Q(r0_2_38_), .QB(n2763), .D(n2907), .CLK(clk_i) );
  dff r0_2_reg_37_ ( .Q(r0_2_37_), .QB(n2762), .D(n2908), .CLK(clk_i) );
  dff r0_2_reg_36_ ( .Q(r0_2_36_), .QB(n2761), .D(n2909), .CLK(clk_i) );
  dff r0_2_reg_35_ ( .Q(r0_2_35_), .QB(n2760), .D(n2910), .CLK(clk_i) );
  dff r0_2_reg_34_ ( .Q(r0_2_34_), .QB(n2759), .D(n2911), .CLK(clk_i) );
  dff r0_2_reg_33_ ( .Q(r0_2_33_), .QB(n2758), .D(n2912), .CLK(clk_i) );
  dff r0_2_reg_32_ ( .Q(r0_2_32_), .QB(n2757), .D(n2913), .CLK(clk_i) );
  dff r0_2_reg_31_ ( .Q(r0_2_31_), .QB(n2756), .D(n2914), .CLK(clk_i) );
  dff r0_2_reg_30_ ( .Q(r0_2_30_), .QB(n2755), .D(n2915), .CLK(clk_i) );
  dff r0_2_reg_29_ ( .Q(r0_2_29_), .QB(n2753), .D(n2916), .CLK(clk_i) );
  dff r0_2_reg_28_ ( .Q(r0_2_28_), .QB(n2752), .D(n2917), .CLK(clk_i) );
  dff r0_2_reg_27_ ( .Q(r0_2_27_), .QB(n2751), .D(n2918), .CLK(clk_i) );
  dff r0_2_reg_26_ ( .Q(r0_2_26_), .QB(n2750), .D(n2919), .CLK(clk_i) );
  dff r0_2_reg_25_ ( .Q(r0_2_25_), .QB(n2749), .D(n2920), .CLK(clk_i) );
  dff r0_2_reg_24_ ( .Q(r0_2_24_), .QB(n2748), .D(n2921), .CLK(clk_i) );
  dff r0_2_reg_23_ ( .Q(r0_2_23_), .QB(n2747), .D(n2922), .CLK(clk_i) );
  dff r0_2_reg_22_ ( .Q(r0_2_22_), .QB(n2746), .D(n2923), .CLK(clk_i) );
  dff r0_2_reg_21_ ( .Q(r0_2_21_), .QB(n2745), .D(n2924), .CLK(clk_i) );
  dff r0_2_reg_20_ ( .Q(r0_2_20_), .QB(n2744), .D(n2925), .CLK(clk_i) );
  dff r0_2_reg_19_ ( .Q(r0_2_19_), .QB(n2742), .D(n2926), .CLK(clk_i) );
  dff r0_2_reg_18_ ( .Q(r0_2_18_), .QB(n2741), .D(n2927), .CLK(clk_i) );
  dff r0_2_reg_17_ ( .Q(r0_2_17_), .QB(n2740), .D(n2928), .CLK(clk_i) );
  dff r0_2_reg_16_ ( .Q(r0_2_16_), .QB(n2739), .D(n2929), .CLK(clk_i) );
  dff r0_2_reg_15_ ( .Q(r0_2_15_), .QB(n2738), .D(n2930), .CLK(clk_i) );
  dff r0_2_reg_14_ ( .Q(r0_2_14_), .QB(n2737), .D(n2931), .CLK(clk_i) );
  dff r0_2_reg_13_ ( .Q(r0_2_13_), .QB(n2736), .D(n2932), .CLK(clk_i) );
  dff r0_2_reg_12_ ( .Q(r0_2_12_), .QB(n2735), .D(n2933), .CLK(clk_i) );
  dff r0_2_reg_11_ ( .Q(r0_2_11_), .QB(n2734), .D(n2934), .CLK(clk_i) );
  dff r0_2_reg_10_ ( .Q(r0_2_10_), .QB(n2733), .D(n2935), .CLK(clk_i) );
  dff r0_2_reg_9_ ( .Q(r0_2_9_), .QB(n2783), .D(n2936), .CLK(clk_i) );
  dff r0_2_reg_8_ ( .Q(r0_2_8_), .QB(n2782), .D(n2937), .CLK(clk_i) );
  dff r0_2_reg_7_ ( .Q(r0_2_7_), .QB(n2781), .D(n2938), .CLK(clk_i) );
  dff r0_2_reg_6_ ( .Q(r0_2_6_), .QB(n2780), .D(n2939), .CLK(clk_i) );
  dff r0_2_reg_5_ ( .Q(r0_2_5_), .QB(n2779), .D(n2940), .CLK(clk_i) );
  dff r0_2_reg_4_ ( .Q(r0_2_4_), .QB(n2776), .D(n2941), .CLK(clk_i) );
  dff r0_2_reg_3_ ( .Q(r0_2_3_), .QB(n2765), .D(n2942), .CLK(clk_i) );
  dff r0_2_reg_2_ ( .Q(r0_2_2_), .QB(n2754), .D(n2943), .CLK(clk_i) );
  dff r0_2_reg_1_ ( .Q(r0_2_1_), .QB(n2743), .D(n2944), .CLK(clk_i) );
  dff r0_2_reg_0_ ( .Q(r0_2_0_), .QB(n2732), .D(n2945), .CLK(clk_i) );
  dff r1_reg_50_ ( .Q(r1_50_), .QB(n2808), .D(n3383), .CLK(clk_i) );
  dff r1_reg_49_ ( .Q(r1_49_), .QB(n2807), .D(n3395), .CLK(clk_i) );
  dff r1_reg_48_ ( .Q(r1_48_), .QB(n2806), .D(n3413), .CLK(clk_i) );
  dff r1_reg_47_ ( .Q(r1_47_), .QB(n2805), .D(n3417), .CLK(clk_i) );
  dff r1_reg_46_ ( .Q(r1_46_), .QB(n2804), .D(n3391), .CLK(clk_i) );
  dff r1_reg_45_ ( .Q(r1_45_), .QB(n2803), .D(n3375), .CLK(clk_i) );
  dff r1_reg_44_ ( .Q(r1_44_), .QB(n2802), .D(n3405), .CLK(clk_i) );
  dff r1_reg_43_ ( .Q(r1_43_), .QB(n2801), .D(n3425), .CLK(clk_i) );
  dff r1_reg_42_ ( .Q(r1_42_), .QB(n2800), .D(n3381), .CLK(clk_i) );
  dff r1_reg_41_ ( .Q(r1_41_), .QB(n2799), .D(n3421), .CLK(clk_i) );
  dff r1_reg_40_ ( .Q(r1_40_), .QB(n2798), .D(n3423), .CLK(clk_i) );
  dff r1_reg_39_ ( .Q(r1_39_), .QB(n2797), .D(n3407), .CLK(clk_i) );
  dff r1_reg_38_ ( .Q(r1_38_), .QB(n2796), .D(n3415), .CLK(clk_i) );
  dff r1_reg_37_ ( .Q(r1_37_), .QB(n2795), .D(n3409), .CLK(clk_i) );
  dff r1_reg_36_ ( .Q(r1_36_), .QB(n2794), .D(n3387), .CLK(clk_i) );
  dff r1_reg_35_ ( .Q(r1_35_), .QB(n2793), .D(n3401), .CLK(clk_i) );
  dff r1_reg_34_ ( .Q(r1_34_), .QB(n2792), .D(n3403), .CLK(clk_i) );
  dff r1_reg_33_ ( .Q(r1_33_), .QB(n2791), .D(n3379), .CLK(clk_i) );
  dff r1_reg_32_ ( .Q(r1_32_), .QB(n2790), .D(n3377), .CLK(clk_i) );
  dff r1_reg_31_ ( .Q(r1_31_), .QB(n2789), .D(n3399), .CLK(clk_i) );
  dff r1_reg_30_ ( .Q(r1_30_), .QB(n2788), .D(n3393), .CLK(clk_i) );
  dff r1_reg_29_ ( .Q(r1_29_), .QB(n2787), .D(n3419), .CLK(clk_i) );
  dff r1_reg_28_ ( .Q(r1_28_), .QB(n2786), .D(n3397), .CLK(clk_i) );
  dff r1_reg_27_ ( .Q(r1_27_), .QB(n2785), .D(n3389), .CLK(clk_i) );
  dff r1_reg_26_ ( .Q(r1_26_), .QB(n2784), .D(n3385), .CLK(clk_i) );
  dff r1_reg_25_ ( .Q(r1_25_), .D(n2971), .CLK(clk_i) );
  dff r1_reg_24_ ( .Q(r1_24_), .D(n2972), .CLK(clk_i) );
  dff r1_reg_23_ ( .Q(r1_23_), .D(n2973), .CLK(clk_i) );
  dff r1_reg_22_ ( .Q(r1_22_), .D(n2974), .CLK(clk_i) );
  dff r1_reg_21_ ( .Q(r1_21_), .D(n2975), .CLK(clk_i) );
  dff r1_reg_20_ ( .Q(r1_20_), .D(n2976), .CLK(clk_i) );
  dff r1_reg_19_ ( .Q(r1_19_), .D(n2977), .CLK(clk_i) );
  dff r1_reg_18_ ( .Q(r1_18_), .D(n2978), .CLK(clk_i) );
  dff r1_reg_17_ ( .Q(r1_17_), .D(n2979), .CLK(clk_i) );
  dff r1_reg_16_ ( .Q(r1_16_), .D(n2980), .CLK(clk_i) );
  dff r1_reg_15_ ( .Q(r1_15_), .D(n2981), .CLK(clk_i) );
  dff r1_reg_14_ ( .Q(r1_14_), .D(n2982), .CLK(clk_i) );
  dff r1_reg_13_ ( .Q(r1_13_), .D(n2983), .CLK(clk_i) );
  dff r1_reg_12_ ( .Q(r1_12_), .D(n2984), .CLK(clk_i) );
  dff r1_reg_11_ ( .Q(r1_11_), .D(n2985), .CLK(clk_i) );
  dff r1_reg_10_ ( .Q(r1_10_), .D(n2986), .CLK(clk_i) );
  dff r1_reg_9_ ( .Q(r1_9_), .D(n2987), .CLK(clk_i) );
  dff r1_reg_8_ ( .Q(r1_8_), .D(n2988), .CLK(clk_i) );
  dff r1_reg_7_ ( .Q(r1_7_), .D(n2989), .CLK(clk_i) );
  dff r1_reg_6_ ( .Q(r1_6_), .D(n2990), .CLK(clk_i) );
  dff r1_reg_5_ ( .Q(r1_5_), .D(n2991), .CLK(clk_i) );
  dff r1_reg_4_ ( .Q(r1_4_), .D(n2992), .CLK(clk_i) );
  dff r1_reg_3_ ( .Q(r1_3_), .D(n2993), .CLK(clk_i) );
  dff r1_reg_2_ ( .Q(r1_2_), .D(n2994), .CLK(clk_i) );
  dff r1_reg_1_ ( .Q(r1_1_), .D(n2995), .CLK(clk_i) );
  dff r1_reg_0_ ( .Q(r1_0_), .D(n2996), .CLK(clk_i) );
  dff r1_2_reg_51_ ( .Q(r1_2_51_), .QB(n6947), .D(n2997), .CLK(clk_i) );
  dff r1_2_reg_50_ ( .Q(r1_2_50_), .QB(n6131), .D(n2998), .CLK(clk_i) );
  dff r1_2_reg_49_ ( .Q(r1_2_49_), .QB(n6163), .D(n2999), .CLK(clk_i) );
  dff r1_2_reg_48_ ( .Q(r1_2_48_), .QB(n6890), .D(n3000), .CLK(clk_i) );
  dff r1_2_reg_47_ ( .Q(r1_2_47_), .QB(n6844), .D(n3001), .CLK(clk_i) );
  dff r1_2_reg_46_ ( .Q(r1_2_46_), .QB(n6882), .D(n3002), .CLK(clk_i) );
  dff r1_2_reg_45_ ( .Q(r1_2_45_), .QB(n6830), .D(n3003), .CLK(clk_i) );
  dff r1_2_reg_44_ ( .Q(r1_2_44_), .QB(n6245), .D(n3004), .CLK(clk_i) );
  dff r1_2_reg_43_ ( .Q(r1_2_43_), .QB(n6171), .D(n3005), .CLK(clk_i) );
  dff r1_2_reg_42_ ( .Q(r1_2_42_), .QB(n6239), .D(n3006), .CLK(clk_i) );
  dff r1_2_reg_41_ ( .Q(r1_2_41_), .QB(n6842), .D(n3007), .CLK(clk_i) );
  dff r1_2_reg_40_ ( .Q(r1_2_40_), .QB(n6872), .D(n3008), .CLK(clk_i) );
  dff r1_2_reg_39_ ( .Q(r1_2_39_), .QB(n6179), .D(n3009), .CLK(clk_i) );
  dff r1_2_reg_38_ ( .Q(r1_2_38_), .QB(n6235), .D(n3010), .CLK(clk_i) );
  dff r1_2_reg_37_ ( .Q(r1_2_37_), .QB(n6169), .D(n3011), .CLK(clk_i) );
  dff r1_2_reg_36_ ( .Q(r1_2_36_), .QB(n6892), .D(n3012), .CLK(clk_i) );
  dff r1_2_reg_35_ ( .Q(r1_2_35_), .QB(n6834), .D(n3013), .CLK(clk_i) );
  dff r1_2_reg_34_ ( .Q(r1_2_34_), .QB(n6878), .D(n3014), .CLK(clk_i) );
  dff r1_2_reg_33_ ( .Q(r1_2_33_), .QB(n6848), .D(n3015), .CLK(clk_i) );
  dff r1_2_reg_32_ ( .Q(r1_2_32_), .QB(n6237), .D(n3016), .CLK(clk_i) );
  dff r1_2_reg_31_ ( .Q(r1_2_31_), .QB(n6183), .D(n3017), .CLK(clk_i) );
  dff r1_2_reg_30_ ( .Q(r1_2_30_), .QB(n6249), .D(n3018), .CLK(clk_i) );
  dff r1_2_reg_29_ ( .Q(r1_2_29_), .QB(n6854), .D(n3019), .CLK(clk_i) );
  dff r1_2_reg_28_ ( .Q(r1_2_28_), .QB(n6874), .D(n3020), .CLK(clk_i) );
  dff r1_2_reg_27_ ( .Q(r1_2_27_), .QB(n6175), .D(n3021), .CLK(clk_i) );
  dff r1_2_reg_26_ ( .Q(r1_2_26_), .QB(n6233), .D(n3022), .CLK(clk_i) );
  dff r1_2_reg_25_ ( .Q(r1_2_25_), .QB(n6181), .D(n3023), .CLK(clk_i) );
  dff r1_2_reg_24_ ( .Q(r1_2_24_), .QB(n6886), .D(n3024), .CLK(clk_i) );
  dff r1_2_reg_23_ ( .Q(r1_2_23_), .QB(n6846), .D(n3025), .CLK(clk_i) );
  dff r1_2_reg_22_ ( .Q(r1_2_22_), .QB(n6868), .D(n3026), .CLK(clk_i) );
  dff r1_2_reg_21_ ( .Q(r1_2_21_), .QB(n6836), .D(n3027), .CLK(clk_i) );
  dff r1_2_reg_20_ ( .Q(r1_2_20_), .QB(n6243), .D(n3028), .CLK(clk_i) );
  dff r1_2_reg_19_ ( .Q(r1_2_19_), .QB(n6167), .D(n3029), .CLK(clk_i) );
  dff r1_2_reg_18_ ( .Q(r1_2_18_), .QB(n6880), .D(n3030), .CLK(clk_i) );
  dff r1_2_reg_17_ ( .Q(r1_2_17_), .QB(n6850), .D(n3031), .CLK(clk_i) );
  dff r1_2_reg_16_ ( .Q(r1_2_16_), .QB(n6876), .D(n3032), .CLK(clk_i) );
  dff r1_2_reg_15_ ( .Q(r1_2_15_), .QB(n6173), .D(n3033), .CLK(clk_i) );
  dff r1_2_reg_14_ ( .Q(r1_2_14_), .QB(n6241), .D(n3034), .CLK(clk_i) );
  dff r1_2_reg_13_ ( .Q(r1_2_13_), .QB(n6165), .D(n3035), .CLK(clk_i) );
  dff r1_2_reg_12_ ( .Q(r1_2_12_), .QB(n6888), .D(n3036), .CLK(clk_i) );
  dff r1_2_reg_11_ ( .Q(r1_2_11_), .QB(n6838), .D(n3037), .CLK(clk_i) );
  dff r1_2_reg_10_ ( .Q(r1_2_10_), .QB(n6852), .D(n3038), .CLK(clk_i) );
  dff r1_2_reg_9_ ( .Q(r1_2_9_), .QB(n6231), .D(n3039), .CLK(clk_i) );
  dff r1_2_reg_8_ ( .Q(r1_2_8_), .QB(n6251), .D(n3040), .CLK(clk_i) );
  dff r1_2_reg_7_ ( .Q(r1_2_7_), .QB(n6177), .D(n3041), .CLK(clk_i) );
  dff r1_2_reg_6_ ( .Q(r1_2_6_), .QB(n6884), .D(n3042), .CLK(clk_i) );
  dff r1_2_reg_5_ ( .Q(r1_2_5_), .QB(n6832), .D(n3043), .CLK(clk_i) );
  dff r1_2_reg_4_ ( .Q(r1_2_4_), .QB(n6247), .D(n3044), .CLK(clk_i) );
  dff r1_2_reg_3_ ( .Q(r1_2_3_), .QB(n6840), .D(n3045), .CLK(clk_i) );
  dff r1_2_reg_2_ ( .Q(r1_2_2_), .QB(n6870), .D(n3046), .CLK(clk_i) );
  dff r1_2_reg_1_ ( .Q(r1_2_1_), .D(n3047), .CLK(clk_i) );
  dff r1_2_reg_0_ ( .Q(r1_2_0_), .D(n3048), .CLK(clk_i) );
  dff s_state_reg ( .Q(s_state), .QB(n6949), .D(n3049), .CLK(clk_i) );
  dff s_ready_o_reg ( .Q(s_ready_o), .QB(n2810), .D(n3050), .CLK(clk_i) );
  dff b_reg_51_ ( .QB(n2731), .D(1'b0), .CLK(clk_i) );
  dff b_2_reg_51_ ( .Q(b_2[51]), .QB(n2730), .D(1'b0), .CLK(clk_i) );
  dff s_sqr_o_reg_25_ ( .Q(s_sqr_o_25_), .QB(n2828), .D(n3051), .CLK(clk_i) );
  dff s_sqr_o_reg_24_ ( .Q(s_sqr_o_24_), .QB(n2827), .D(n3052), .CLK(clk_i) );
  dff s_sqr_o_reg_23_ ( .Q(s_sqr_o_23_), .QB(n2826), .D(n3053), .CLK(clk_i) );
  dff s_sqr_o_reg_22_ ( .Q(s_sqr_o_22_), .QB(n2825), .D(n3054), .CLK(clk_i) );
  dff s_sqr_o_reg_21_ ( .Q(s_sqr_o_21_), .QB(n2824), .D(n3055), .CLK(clk_i) );
  dff s_sqr_o_reg_20_ ( .Q(s_sqr_o_20_), .QB(n2823), .D(n3056), .CLK(clk_i) );
  dff s_sqr_o_reg_19_ ( .Q(s_sqr_o_19_), .QB(n2821), .D(n3057), .CLK(clk_i) );
  dff s_sqr_o_reg_18_ ( .Q(s_sqr_o_18_), .QB(n2820), .D(n3058), .CLK(clk_i) );
  dff s_sqr_o_reg_17_ ( .Q(s_sqr_o_17_), .QB(n2819), .D(n3059), .CLK(clk_i) );
  dff s_sqr_o_reg_16_ ( .Q(s_sqr_o_16_), .QB(n2818), .D(n3060), .CLK(clk_i) );
  dff s_sqr_o_reg_15_ ( .Q(s_sqr_o_15_), .QB(n2817), .D(n3061), .CLK(clk_i) );
  dff s_sqr_o_reg_14_ ( .Q(s_sqr_o_14_), .QB(n2816), .D(n3062), .CLK(clk_i) );
  dff s_sqr_o_reg_13_ ( .Q(s_sqr_o_13_), .QB(n2815), .D(n3063), .CLK(clk_i) );
  dff s_sqr_o_reg_12_ ( .Q(s_sqr_o_12_), .QB(n2814), .D(n3064), .CLK(clk_i) );
  dff s_sqr_o_reg_11_ ( .Q(s_sqr_o_11_), .QB(n2813), .D(n3065), .CLK(clk_i) );
  dff s_sqr_o_reg_10_ ( .Q(s_sqr_o_10_), .QB(n2812), .D(n3066), .CLK(clk_i) );
  dff s_sqr_o_reg_9_ ( .Q(s_sqr_o_9_), .QB(n2836), .D(n3067), .CLK(clk_i) );
  dff s_sqr_o_reg_8_ ( .Q(s_sqr_o_8_), .QB(n2835), .D(n3068), .CLK(clk_i) );
  dff s_sqr_o_reg_7_ ( .Q(s_sqr_o_7_), .QB(n2834), .D(n3069), .CLK(clk_i) );
  dff s_sqr_o_reg_6_ ( .Q(s_sqr_o_6_), .QB(n2833), .D(n3070), .CLK(clk_i) );
  dff s_sqr_o_reg_5_ ( .Q(s_sqr_o_5_), .QB(n2832), .D(n3071), .CLK(clk_i) );
  dff s_sqr_o_reg_4_ ( .Q(s_sqr_o_4_), .QB(n2831), .D(n3072), .CLK(clk_i) );
  dff s_sqr_o_reg_3_ ( .Q(s_sqr_o_3_), .QB(n2830), .D(n3073), .CLK(clk_i) );
  dff s_sqr_o_reg_2_ ( .Q(s_sqr_o_2_), .QB(n2829), .D(n3074), .CLK(clk_i) );
  dff s_sqr_o_reg_1_ ( .Q(s_sqr_o_1_), .QB(n2822), .D(n3075), .CLK(clk_i) );
  dff s_sqr_o_reg_0_ ( .Q(s_sqr_o_0_), .QB(n2811), .D(n3076), .CLK(clk_i) );
  dff s_ine_o_reg ( .Q(s_ine_o), .QB(n2809), .D(n3077), .CLK(clk_i) );
  dff s_rad_i_reg_51_ ( .Q(s_rad_i_51_), .D(rad_i[51]), .CLK(clk_i) );
  dff s_rad_i_reg_50_ ( .Q(s_rad_i_50_), .D(rad_i[50]), .CLK(clk_i) );
  dff s_rad_i_reg_49_ ( .Q(s_rad_i_49_), .D(rad_i[49]), .CLK(clk_i) );
  dff s_rad_i_reg_48_ ( .Q(s_rad_i_48_), .D(rad_i[48]), .CLK(clk_i) );
  dff s_rad_i_reg_47_ ( .Q(s_rad_i_47_), .D(rad_i[47]), .CLK(clk_i) );
  dff s_rad_i_reg_46_ ( .Q(s_rad_i_46_), .D(rad_i[46]), .CLK(clk_i) );
  dff s_rad_i_reg_45_ ( .Q(s_rad_i_45_), .D(rad_i[45]), .CLK(clk_i) );
  dff s_rad_i_reg_44_ ( .Q(s_rad_i_44_), .D(rad_i[44]), .CLK(clk_i) );
  dff s_rad_i_reg_43_ ( .Q(s_rad_i_43_), .D(rad_i[43]), .CLK(clk_i) );
  dff s_rad_i_reg_42_ ( .Q(s_rad_i_42_), .D(rad_i[42]), .CLK(clk_i) );
  dff s_rad_i_reg_41_ ( .Q(s_rad_i_41_), .D(rad_i[41]), .CLK(clk_i) );
  dff s_rad_i_reg_40_ ( .Q(s_rad_i_40_), .D(rad_i[40]), .CLK(clk_i) );
  dff s_rad_i_reg_39_ ( .Q(s_rad_i_39_), .D(rad_i[39]), .CLK(clk_i) );
  dff s_rad_i_reg_38_ ( .Q(s_rad_i_38_), .D(rad_i[38]), .CLK(clk_i) );
  dff s_rad_i_reg_37_ ( .Q(s_rad_i_37_), .D(rad_i[37]), .CLK(clk_i) );
  dff s_rad_i_reg_36_ ( .Q(s_rad_i_36_), .D(rad_i[36]), .CLK(clk_i) );
  dff s_rad_i_reg_35_ ( .Q(s_rad_i_35_), .D(rad_i[35]), .CLK(clk_i) );
  dff s_rad_i_reg_34_ ( .Q(s_rad_i_34_), .D(rad_i[34]), .CLK(clk_i) );
  dff s_rad_i_reg_33_ ( .Q(s_rad_i_33_), .D(rad_i[33]), .CLK(clk_i) );
  dff s_rad_i_reg_32_ ( .Q(s_rad_i_32_), .D(rad_i[32]), .CLK(clk_i) );
  dff s_rad_i_reg_31_ ( .Q(s_rad_i_31_), .D(rad_i[31]), .CLK(clk_i) );
  dff s_rad_i_reg_30_ ( .Q(s_rad_i_30_), .D(rad_i[30]), .CLK(clk_i) );
  dff s_rad_i_reg_29_ ( .Q(s_rad_i_29_), .D(rad_i[29]), .CLK(clk_i) );
  dff s_rad_i_reg_28_ ( .Q(s_rad_i_28_), .D(rad_i[28]), .CLK(clk_i) );
  dff s_rad_i_reg_27_ ( .Q(s_rad_i_27_), .D(rad_i[27]), .CLK(clk_i) );
  dff s_rad_i_reg_26_ ( .Q(s_rad_i_26_), .D(rad_i[26]), .CLK(clk_i) );
  dff s_rad_i_reg_25_ ( .Q(s_rad_i_25_), .D(rad_i[25]), .CLK(clk_i) );
  dff s_rad_i_reg_24_ ( .Q(s_rad_i_24_), .D(rad_i[24]), .CLK(clk_i) );
  dff s_rad_i_reg_23_ ( .Q(s_rad_i_23_), .D(rad_i[23]), .CLK(clk_i) );
  dff s_rad_i_reg_22_ ( .Q(s_rad_i_22_), .D(rad_i[22]), .CLK(clk_i) );
  dff s_rad_i_reg_21_ ( .Q(s_rad_i_21_), .D(rad_i[21]), .CLK(clk_i) );
  dff s_rad_i_reg_20_ ( .Q(s_rad_i_20_), .D(rad_i[20]), .CLK(clk_i) );
  dff s_rad_i_reg_19_ ( .Q(s_rad_i_19_), .D(rad_i[19]), .CLK(clk_i) );
  dff s_rad_i_reg_18_ ( .Q(s_rad_i_18_), .D(rad_i[18]), .CLK(clk_i) );
  dff s_rad_i_reg_17_ ( .Q(s_rad_i_17_), .D(rad_i[17]), .CLK(clk_i) );
  dff s_rad_i_reg_16_ ( .Q(s_rad_i_16_), .D(rad_i[16]), .CLK(clk_i) );
  dff s_rad_i_reg_15_ ( .Q(s_rad_i_15_), .D(rad_i[15]), .CLK(clk_i) );
  dff s_rad_i_reg_14_ ( .Q(s_rad_i_14_), .D(rad_i[14]), .CLK(clk_i) );
  dff s_rad_i_reg_13_ ( .Q(s_rad_i_13_), .D(rad_i[13]), .CLK(clk_i) );
  dff s_rad_i_reg_12_ ( .Q(s_rad_i_12_), .D(rad_i[12]), .CLK(clk_i) );
  dff s_rad_i_reg_11_ ( .Q(s_rad_i_11_), .D(rad_i[11]), .CLK(clk_i) );
  dff s_rad_i_reg_10_ ( .Q(s_rad_i_10_), .D(rad_i[10]), .CLK(clk_i) );
  dff s_rad_i_reg_9_ ( .Q(s_rad_i_9_), .D(rad_i[9]), .CLK(clk_i) );
  dff s_rad_i_reg_8_ ( .Q(s_rad_i_8_), .D(rad_i[8]), .CLK(clk_i) );
  dff s_rad_i_reg_7_ ( .Q(s_rad_i_7_), .D(rad_i[7]), .CLK(clk_i) );
  dff s_rad_i_reg_6_ ( .Q(s_rad_i_6_), .D(rad_i[6]), .CLK(clk_i) );
  dff s_rad_i_reg_5_ ( .Q(s_rad_i_5_), .D(rad_i[5]), .CLK(clk_i) );
  dff s_rad_i_reg_4_ ( .Q(s_rad_i_4_), .D(rad_i[4]), .CLK(clk_i) );
  dff s_rad_i_reg_3_ ( .Q(s_rad_i_3_), .D(rad_i[3]), .CLK(clk_i) );
  dff s_rad_i_reg_2_ ( .Q(s_rad_i_2_), .D(rad_i[2]), .CLK(clk_i) );
  dff s_rad_i_reg_1_ ( .Q(s_rad_i_1_), .D(rad_i[1]), .CLK(clk_i) );
  dff s_rad_i_reg_0_ ( .Q(s_rad_i_0_), .D(rad_i[0]), .CLK(clk_i) );
  dff sqr_o_reg_25_ ( .Q(sqr_o[25]), .D(s_sqr_o_25_), .CLK(clk_i) );
  dff sqr_o_reg_24_ ( .Q(sqr_o[24]), .D(s_sqr_o_24_), .CLK(clk_i) );
  dff sqr_o_reg_23_ ( .Q(sqr_o[23]), .D(s_sqr_o_23_), .CLK(clk_i) );
  dff sqr_o_reg_22_ ( .Q(sqr_o[22]), .D(s_sqr_o_22_), .CLK(clk_i) );
  dff sqr_o_reg_21_ ( .Q(sqr_o[21]), .D(s_sqr_o_21_), .CLK(clk_i) );
  dff sqr_o_reg_20_ ( .Q(sqr_o[20]), .D(s_sqr_o_20_), .CLK(clk_i) );
  dff sqr_o_reg_19_ ( .Q(sqr_o[19]), .D(s_sqr_o_19_), .CLK(clk_i) );
  dff sqr_o_reg_18_ ( .Q(sqr_o[18]), .D(s_sqr_o_18_), .CLK(clk_i) );
  dff sqr_o_reg_17_ ( .Q(sqr_o[17]), .D(s_sqr_o_17_), .CLK(clk_i) );
  dff sqr_o_reg_16_ ( .Q(sqr_o[16]), .D(s_sqr_o_16_), .CLK(clk_i) );
  dff sqr_o_reg_15_ ( .Q(sqr_o[15]), .D(s_sqr_o_15_), .CLK(clk_i) );
  dff sqr_o_reg_14_ ( .Q(sqr_o[14]), .D(s_sqr_o_14_), .CLK(clk_i) );
  dff sqr_o_reg_13_ ( .Q(sqr_o[13]), .D(s_sqr_o_13_), .CLK(clk_i) );
  dff sqr_o_reg_12_ ( .Q(sqr_o[12]), .D(s_sqr_o_12_), .CLK(clk_i) );
  dff sqr_o_reg_11_ ( .Q(sqr_o[11]), .D(s_sqr_o_11_), .CLK(clk_i) );
  dff sqr_o_reg_10_ ( .Q(sqr_o[10]), .D(s_sqr_o_10_), .CLK(clk_i) );
  dff sqr_o_reg_9_ ( .Q(sqr_o[9]), .D(s_sqr_o_9_), .CLK(clk_i) );
  dff sqr_o_reg_8_ ( .Q(sqr_o[8]), .D(s_sqr_o_8_), .CLK(clk_i) );
  dff sqr_o_reg_7_ ( .Q(sqr_o[7]), .D(s_sqr_o_7_), .CLK(clk_i) );
  dff sqr_o_reg_6_ ( .Q(sqr_o[6]), .D(s_sqr_o_6_), .CLK(clk_i) );
  dff sqr_o_reg_5_ ( .Q(sqr_o[5]), .D(s_sqr_o_5_), .CLK(clk_i) );
  dff sqr_o_reg_4_ ( .Q(sqr_o[4]), .D(s_sqr_o_4_), .CLK(clk_i) );
  dff sqr_o_reg_3_ ( .Q(sqr_o[3]), .D(s_sqr_o_3_), .CLK(clk_i) );
  dff sqr_o_reg_2_ ( .Q(sqr_o[2]), .D(s_sqr_o_2_), .CLK(clk_i) );
  dff sqr_o_reg_1_ ( .Q(sqr_o[1]), .D(s_sqr_o_1_), .CLK(clk_i) );
  dff sqr_o_reg_0_ ( .Q(sqr_o[0]), .D(s_sqr_o_0_), .CLK(clk_i) );
  dff c_reg_4_ ( .Q(c_4_), .D(c222_4_), .CLK(clk_i) );
  dff c_reg_3_ ( .Q(c_3_), .D(c222_3_), .CLK(clk_i) );
  dff c_reg_2_ ( .Q(c_2_), .D(c222_2_), .CLK(clk_i) );
  dff c_reg_1_ ( .Q(c_1_), .D(c222_1_), .CLK(clk_i) );
  dff c_reg_0_ ( .Q(c_0_), .QB(n6575), .D(c222_0_), .CLK(clk_i) );
  dff s_start_i_reg ( .Q(s_state110), .D(start_i), .CLK(clk_i) );
  dff ine_o_reg ( .Q(ine_o), .D(s_ine_o), .CLK(clk_i) );
  dff ready_o_reg ( .Q(ready_o), .D(s_ready_o), .CLK(clk_i) );
  dff b_reg_50_ ( .QB(n1930), .D(n3966), .CLK(clk_i) );
  dff b_reg_49_ ( .QB(n1929), .D(n3980), .CLK(clk_i) );
  dff b_reg_48_ ( .QB(n1928), .D(n3842), .CLK(clk_i) );
  dff b_reg_47_ ( .QB(n1927), .D(n4024), .CLK(clk_i) );
  dff b_reg_46_ ( .QB(n1926), .D(n3880), .CLK(clk_i) );
  dff b_reg_45_ ( .QB(n1925), .D(n3872), .CLK(clk_i) );
  dff b_reg_44_ ( .QB(n1924), .D(n3988), .CLK(clk_i) );
  dff b_reg_43_ ( .QB(n1923), .D(n3976), .CLK(clk_i) );
  dff b_reg_42_ ( .QB(n1922), .D(n3870), .CLK(clk_i) );
  dff b_reg_41_ ( .QB(n1921), .D(n3990), .CLK(clk_i) );
  dff b_reg_40_ ( .QB(n1920), .D(n3958), .CLK(clk_i) );
  dff b_reg_39_ ( .QB(n1919), .D(n4022), .CLK(clk_i) );
  dff b_reg_38_ ( .QB(n1918), .D(n3876), .CLK(clk_i) );
  dff b_reg_37_ ( .QB(n1917), .D(n3902), .CLK(clk_i) );
  dff b_reg_36_ ( .QB(n1916), .D(n4012), .CLK(clk_i) );
  dff b_reg_35_ ( .QB(n1915), .D(n3908), .CLK(clk_i) );
  dff b_reg_34_ ( .QB(n1914), .D(n3904), .CLK(clk_i) );
  dff b_reg_33_ ( .QB(n1913), .D(n3996), .CLK(clk_i) );
  dff b_reg_32_ ( .QB(n1912), .D(n3926), .CLK(clk_i) );
  dff b_reg_31_ ( .QB(n1911), .D(n3916), .CLK(clk_i) );
  dff b_reg_30_ ( .QB(n1910), .D(n3992), .CLK(clk_i) );
  dff b_reg_29_ ( .QB(n1909), .D(n3974), .CLK(clk_i) );
  dff b_reg_28_ ( .QB(n1908), .D(n3936), .CLK(clk_i) );
  dff b_reg_27_ ( .QB(n1907), .D(n3862), .CLK(clk_i) );
  dff b_reg_26_ ( .QB(n1906), .D(n3948), .CLK(clk_i) );
  dff b_reg_25_ ( .Q(b_25_), .QB(n1905), .D(b206_25_), .CLK(clk_i) );
  dff b_reg_24_ ( .Q(b_24_), .QB(n1904), .D(n4030), .CLK(clk_i) );
  dff b_reg_23_ ( .Q(b_23_), .QB(n1903), .D(n3854), .CLK(clk_i) );
  dff b_reg_22_ ( .Q(b_22_), .QB(n1902), .D(n3932), .CLK(clk_i) );
  dff b_reg_21_ ( .Q(b_21_), .QB(n1901), .D(n3964), .CLK(clk_i) );
  dff b_reg_20_ ( .Q(b_20_), .QB(n1900), .D(n3864), .CLK(clk_i) );
  dff b_reg_19_ ( .Q(b_19_), .QB(n1899), .D(n4018), .CLK(clk_i) );
  dff b_reg_18_ ( .Q(b_18_), .QB(n1898), .D(n3868), .CLK(clk_i) );
  dff b_reg_17_ ( .Q(b_17_), .QB(n1897), .D(n3856), .CLK(clk_i) );
  dff b_reg_16_ ( .Q(b_16_), .QB(n1896), .D(n3994), .CLK(clk_i) );
  dff b_reg_15_ ( .Q(b_15_), .QB(n1895), .D(n3882), .CLK(clk_i) );
  dff b_reg_14_ ( .Q(b_14_), .QB(n1894), .D(n3928), .CLK(clk_i) );
  dff b_reg_13_ ( .Q(b_13_), .QB(n1893), .D(n3962), .CLK(clk_i) );
  dff b_reg_12_ ( .Q(b_12_), .QB(n1892), .D(n3878), .CLK(clk_i) );
  dff b_reg_11_ ( .Q(b_11_), .QB(n1891), .D(n3944), .CLK(clk_i) );
  dff b_reg_10_ ( .Q(b_10_), .QB(n1890), .D(n3950), .CLK(clk_i) );
  dff b_reg_9_ ( .Q(b_9_), .QB(n1889), .D(n4000), .CLK(clk_i) );
  dff b_reg_8_ ( .Q(b_8_), .QB(n1888), .D(n3942), .CLK(clk_i) );
  dff b_reg_7_ ( .Q(b_7_), .QB(n1887), .D(n3898), .CLK(clk_i) );
  dff b_reg_6_ ( .Q(b_6_), .QB(n1886), .D(n4010), .CLK(clk_i) );
  dff b_reg_5_ ( .Q(b_5_), .QB(n1885), .D(n3978), .CLK(clk_i) );
  dff b_reg_4_ ( .Q(b_4_), .QB(n1884), .D(n3934), .CLK(clk_i) );
  dff b_reg_3_ ( .Q(b_3_), .QB(n1883), .D(n3972), .CLK(clk_i) );
  dff b_reg_2_ ( .Q(b_2_), .QB(n1882), .D(n3894), .CLK(clk_i) );
  dff b_reg_1_ ( .Q(b_1_), .QB(n1881), .D(n3924), .CLK(clk_i) );
  dff b_reg_0_ ( .Q(b_0_), .D(n3940), .CLK(clk_i) );
  dff b_2_reg_50_ ( .Q(b_2[50]), .QB(n1880), .D(n7420), .CLK(clk_i) );
  dff b_2_reg_49_ ( .Q(b_2[49]), .QB(n1879), .D(n3896), .CLK(clk_i) );
  dff b_2_reg_48_ ( .Q(b_2[48]), .QB(n1878), .D(n4036), .CLK(clk_i) );
  dff b_2_reg_47_ ( .Q(b_2[47]), .QB(n1877), .D(n4038), .CLK(clk_i) );
  dff b_2_reg_46_ ( .Q(b_2[46]), .QB(n1876), .D(n3850), .CLK(clk_i) );
  dff b_2_reg_45_ ( .Q(b_2[45]), .QB(n1875), .D(n3858), .CLK(clk_i) );
  dff b_2_reg_44_ ( .Q(b_2[44]), .QB(n1874), .D(n4016), .CLK(clk_i) );
  dff b_2_reg_43_ ( .Q(b_2[43]), .QB(n1873), .D(n3892), .CLK(clk_i) );
  dff b_2_reg_42_ ( .Q(b_2[42]), .QB(n1872), .D(n3846), .CLK(clk_i) );
  dff b_2_reg_41_ ( .Q(b_2[41]), .QB(n1871), .D(n4028), .CLK(clk_i) );
  dff b_2_reg_40_ ( .Q(b_2[40]), .QB(n1870), .D(n3918), .CLK(clk_i) );
  dff b_2_reg_39_ ( .Q(b_2[39]), .QB(n1869), .D(n4008), .CLK(clk_i) );
  dff b_2_reg_38_ ( .Q(b_2[38]), .QB(n1868), .D(n3852), .CLK(clk_i) );
  dff b_2_reg_37_ ( .Q(b_2[37]), .QB(n1867), .D(n3900), .CLK(clk_i) );
  dff b_2_reg_36_ ( .Q(b_2[36]), .QB(n1866), .D(n4020), .CLK(clk_i) );
  dff b_2_reg_35_ ( .Q(b_2[35]), .QB(n1865), .D(n3866), .CLK(clk_i) );
  dff b_2_reg_34_ ( .Q(b_2[34]), .QB(n1864), .D(n3884), .CLK(clk_i) );
  dff b_2_reg_33_ ( .Q(b_2[33]), .QB(n1863), .D(n3982), .CLK(clk_i) );
  dff b_2_reg_32_ ( .Q(b_2[32]), .QB(n1862), .D(n3888), .CLK(clk_i) );
  dff b_2_reg_31_ ( .Q(b_2[31]), .QB(n1861), .D(n3848), .CLK(clk_i) );
  dff b_2_reg_30_ ( .Q(b_2[30]), .QB(n1860), .D(n4026), .CLK(clk_i) );
  dff b_2_reg_29_ ( .Q(b_2[29]), .QB(n1859), .D(n3890), .CLK(clk_i) );
  dff b_2_reg_28_ ( .Q(b_2[28]), .QB(n1858), .D(n3986), .CLK(clk_i) );
  dff b_2_reg_27_ ( .Q(b_2[27]), .QB(n1857), .D(n3922), .CLK(clk_i) );
  dff b_2_reg_26_ ( .Q(b_2[26]), .QB(n1856), .D(n3930), .CLK(clk_i) );
  dff b_2_reg_25_ ( .Q(b_2[25]), .QB(n1855), .D(n4014), .CLK(clk_i) );
  dff b_2_reg_24_ ( .Q(b_2[24]), .QB(n1854), .D(n3956), .CLK(clk_i) );
  dff b_2_reg_23_ ( .Q(b_2[23]), .QB(n1853), .D(n3970), .CLK(clk_i) );
  dff b_2_reg_22_ ( .Q(b_2[22]), .QB(n1852), .D(n4032), .CLK(clk_i) );
  dff b_2_reg_21_ ( .Q(b_2[21]), .QB(n1851), .D(n3952), .CLK(clk_i) );
  dff b_2_reg_20_ ( .Q(b_2[20]), .QB(n1850), .D(n3860), .CLK(clk_i) );
  dff b_2_reg_19_ ( .Q(b_2[19]), .QB(n1849), .D(n3954), .CLK(clk_i) );
  dff b_2_reg_18_ ( .Q(b_2[18]), .QB(n1848), .D(n3912), .CLK(clk_i) );
  dff b_2_reg_17_ ( .Q(b_2[17]), .QB(n1847), .D(n4034), .CLK(clk_i) );
  dff b_2_reg_16_ ( .Q(b_2[16]), .QB(n1846), .D(n3938), .CLK(clk_i) );
  dff b_2_reg_15_ ( .Q(b_2[15]), .QB(n1845), .D(n3840), .CLK(clk_i) );
  dff b_2_reg_14_ ( .Q(b_2[14]), .QB(n1844), .D(n3968), .CLK(clk_i) );
  dff b_2_reg_13_ ( .Q(b_2[13]), .QB(n1843), .D(n3910), .CLK(clk_i) );
  dff b_2_reg_12_ ( .Q(b_2[12]), .QB(n1842), .D(n3914), .CLK(clk_i) );
  dff b_2_reg_11_ ( .Q(b_2[11]), .QB(n1841), .D(n4004), .CLK(clk_i) );
  dff b_2_reg_10_ ( .Q(b_2[10]), .QB(n1840), .D(n3920), .CLK(clk_i) );
  dff b_2_reg_9_ ( .Q(b_2[9]), .QB(n1839), .D(n4006), .CLK(clk_i) );
  dff b_2_reg_8_ ( .Q(b_2[8]), .QB(n1838), .D(n3886), .CLK(clk_i) );
  dff b_2_reg_7_ ( .Q(b_2[7]), .QB(n1837), .D(n3960), .CLK(clk_i) );
  dff b_2_reg_6_ ( .Q(b_2[6]), .QB(n1836), .D(n3998), .CLK(clk_i) );
  dff b_2_reg_5_ ( .Q(b_2[5]), .QB(n1835), .D(n3874), .CLK(clk_i) );
  dff b_2_reg_4_ ( .Q(b_2[4]), .QB(n1834), .D(n3984), .CLK(clk_i) );
  dff b_2_reg_3_ ( .Q(b_2[3]), .QB(n1833), .D(n3946), .CLK(clk_i) );
  dff b_2_reg_2_ ( .Q(b_2[2]), .QB(n1832), .D(n3906), .CLK(clk_i) );
  dff b_2_reg_1_ ( .Q(b_2[1]), .D(n4002), .CLK(clk_i) );
  dff b_2_reg_0_ ( .Q(b_2[0]), .D(n3844), .CLK(clk_i) );
  buf12 U1467 ( .Y(n7369), .A(n7448) );
  inv04 U1468 ( .Y(n6906), .A(n7658) );
  ao22 U1469 ( .Y(n3078), .A0(n7600), .A1(c_2_), .B0(n7599), .B1(n7651) );
  inv01 U1470 ( .Y(n3079), .A(n3078) );
  inv01 U1471 ( .Y(s_op2_6_), .A(n3080) );
  nor02 U1472 ( .Y(n3081), .A0(n7364), .A1(n7439) );
  nor02 U1473 ( .Y(n3082), .A0(n7440), .A1(n7437) );
  nor02 U1474 ( .Y(n3080), .A0(n3081), .A1(n3082) );
  inv01 U1475 ( .Y(s_op2_5_), .A(n3083) );
  nor02 U1476 ( .Y(n3084), .A0(n7366), .A1(n7439) );
  nor02 U1477 ( .Y(n3085), .A0(n7442), .A1(n7437) );
  nor02 U1478 ( .Y(n3083), .A0(n3084), .A1(n3085) );
  or02 U1479 ( .Y(n3086), .A0(n7453), .A1(n7433) );
  inv01 U1480 ( .Y(n3087), .A(n3086) );
  xor2 U1481 ( .Y(n3088), .A0(s_rad_i_7_), .A1(n7742) );
  inv01 U1482 ( .Y(n3089), .A(n3088) );
  or02 U1483 ( .Y(n3090), .A0(n7535), .A1(n7433) );
  inv01 U1484 ( .Y(n3091), .A(n3090) );
  or02 U1485 ( .Y(n3092), .A0(n7498), .A1(n7433) );
  inv01 U1486 ( .Y(n3093), .A(n3092) );
  or02 U1487 ( .Y(n3094), .A0(n7541), .A1(n7433) );
  inv01 U1488 ( .Y(n3095), .A(n3094) );
  or02 U1489 ( .Y(n3096), .A0(n7492), .A1(n7433) );
  inv01 U1490 ( .Y(n3097), .A(n3096) );
  xor2 U1491 ( .Y(n3098), .A0(s_rad_i_15_), .A1(n7752) );
  inv01 U1492 ( .Y(n3099), .A(n3098) );
  xor2 U1493 ( .Y(n3100), .A0(s_rad_i_13_), .A1(n7751) );
  inv01 U1494 ( .Y(n3101), .A(n3100) );
  or02 U1495 ( .Y(n3102), .A0(n7563), .A1(n7433) );
  inv01 U1496 ( .Y(n3103), .A(n3102) );
  or02 U1497 ( .Y(n3104), .A0(n7524), .A1(n7433) );
  inv01 U1498 ( .Y(n3105), .A(n3104) );
  xor2 U1499 ( .Y(n3106), .A0(s_rad_i_43_), .A1(n7732) );
  inv01 U1500 ( .Y(n3107), .A(n3106) );
  xor2 U1501 ( .Y(n3108), .A0(s_rad_i_27_), .A1(n7762) );
  inv01 U1502 ( .Y(n3109), .A(n3108) );
  xor2 U1503 ( .Y(n3110), .A0(s_rad_i_31_), .A1(n7768) );
  inv01 U1504 ( .Y(n3111), .A(n3110) );
  xor2 U1505 ( .Y(n3112), .A0(s_rad_i_25_), .A1(n7761) );
  inv01 U1506 ( .Y(n3113), .A(n3112) );
  xor2 U1507 ( .Y(n3114), .A0(s_rad_i_39_), .A1(n7725) );
  inv01 U1508 ( .Y(n3115), .A(n3114) );
  xor2 U1509 ( .Y(n3116), .A0(s_rad_i_19_), .A1(n7756) );
  inv01 U1510 ( .Y(n3117), .A(n3116) );
  xor2 U1511 ( .Y(n3118), .A0(s_rad_i_37_), .A1(n7724) );
  inv01 U1512 ( .Y(n3119), .A(n3118) );
  xor2 U1513 ( .Y(n3120), .A0(s_rad_i_49_), .A1(n7736) );
  inv01 U1514 ( .Y(n3121), .A(n3120) );
  or02 U1515 ( .Y(n3122), .A0(n7465), .A1(n7432) );
  inv01 U1516 ( .Y(n3123), .A(n3122) );
  or02 U1517 ( .Y(n3124), .A0(n7559), .A1(n7432) );
  inv01 U1518 ( .Y(n3125), .A(n3124) );
  ao22 U1519 ( .Y(n3126), .A0(ARG1118_1_), .A1(n7771), .B0(r1_1_), .B1(n7389)
         );
  inv01 U1520 ( .Y(n3127), .A(n3126) );
  or02 U1521 ( .Y(n3128), .A0(n7520), .A1(n7432) );
  inv01 U1522 ( .Y(n3129), .A(n3128) );
  or02 U1523 ( .Y(n3130), .A0(n7504), .A1(n7432) );
  inv01 U1524 ( .Y(n3131), .A(n3130) );
  or02 U1525 ( .Y(n3132), .A0(n7555), .A1(n7432) );
  inv01 U1526 ( .Y(n3133), .A(n3132) );
  or02 U1527 ( .Y(n3134), .A0(n7550), .A1(n7432) );
  inv01 U1528 ( .Y(n3135), .A(n3134) );
  or02 U1529 ( .Y(n3136), .A0(n7574), .A1(n7432) );
  inv01 U1530 ( .Y(n3137), .A(n3136) );
  or02 U1531 ( .Y(n3138), .A0(n7464), .A1(n7432) );
  inv01 U1532 ( .Y(n3139), .A(n3138) );
  or02 U1533 ( .Y(n3140), .A0(n7556), .A1(n7431) );
  inv01 U1534 ( .Y(n3141), .A(n3140) );
  or02 U1535 ( .Y(n3142), .A0(n7493), .A1(n7431) );
  inv01 U1536 ( .Y(n3143), .A(n3142) );
  or02 U1537 ( .Y(n3144), .A0(n7573), .A1(n7431) );
  inv01 U1538 ( .Y(n3145), .A(n3144) );
  or02 U1539 ( .Y(n3146), .A0(n7474), .A1(n7431) );
  inv01 U1540 ( .Y(n3147), .A(n3146) );
  nand02 U1541 ( .Y(n7786), .A0(n3148), .A1(n3149) );
  inv01 U1542 ( .Y(n3150), .A(n7389) );
  inv01 U1543 ( .Y(n3151), .A(n7771) );
  inv01 U1544 ( .Y(n3152), .A(ARG1118_23_) );
  inv01 U1545 ( .Y(n3153), .A(r1_23_) );
  nand02 U1546 ( .Y(n3154), .A0(n3150), .A1(n3151) );
  nand02 U1547 ( .Y(n3155), .A0(n3150), .A1(n3152) );
  nand02 U1548 ( .Y(n3156), .A0(n3151), .A1(n3153) );
  nand02 U1549 ( .Y(n3157), .A0(n3152), .A1(n3153) );
  nand02 U1550 ( .Y(n3158), .A0(n3154), .A1(n3155) );
  inv01 U1551 ( .Y(n3148), .A(n3158) );
  nand02 U1552 ( .Y(n3159), .A0(n3156), .A1(n3157) );
  inv01 U1553 ( .Y(n3149), .A(n3159) );
  ao22 U1554 ( .Y(n3160), .A0(ARG1118_15_), .A1(n7771), .B0(r1_15_), .B1(n7389) );
  inv01 U1555 ( .Y(n3161), .A(n3160) );
  or02 U1556 ( .Y(n3162), .A0(n7515), .A1(n7431) );
  inv01 U1557 ( .Y(n3163), .A(n3162) );
  or02 U1558 ( .Y(n3164), .A0(n7480), .A1(n7431) );
  inv01 U1559 ( .Y(n3165), .A(n3164) );
  or02 U1560 ( .Y(n3166), .A0(n7534), .A1(n7431) );
  inv01 U1561 ( .Y(n3167), .A(n3166) );
  or02 U1562 ( .Y(n3168), .A0(n7514), .A1(n7431) );
  inv01 U1563 ( .Y(n3169), .A(n3168) );
  nand02 U1564 ( .Y(n7770), .A0(n3170), .A1(n3171) );
  inv01 U1565 ( .Y(n3172), .A(n7389) );
  inv01 U1566 ( .Y(n3173), .A(n7771) );
  inv01 U1567 ( .Y(n3174), .A(ARG1118_0_) );
  inv01 U1568 ( .Y(n3175), .A(r1_0_) );
  nand02 U1569 ( .Y(n3176), .A0(n3172), .A1(n3173) );
  nand02 U1570 ( .Y(n3177), .A0(n3172), .A1(n3174) );
  nand02 U1571 ( .Y(n3178), .A0(n3173), .A1(n3175) );
  nand02 U1572 ( .Y(n3179), .A0(n3174), .A1(n3175) );
  nand02 U1573 ( .Y(n3180), .A0(n3176), .A1(n3177) );
  inv01 U1574 ( .Y(n3170), .A(n3180) );
  nand02 U1575 ( .Y(n3181), .A0(n3178), .A1(n3179) );
  inv01 U1576 ( .Y(n3171), .A(n3181) );
  nand02 U1577 ( .Y(n7776), .A0(n3182), .A1(n3183) );
  inv01 U1578 ( .Y(n3184), .A(n7389) );
  inv01 U1579 ( .Y(n3185), .A(n7771) );
  inv01 U1580 ( .Y(n3186), .A(ARG1118_9_) );
  inv01 U1581 ( .Y(n3187), .A(r1_9_) );
  nand02 U1582 ( .Y(n3188), .A0(n3184), .A1(n3185) );
  nand02 U1583 ( .Y(n3189), .A0(n3184), .A1(n3186) );
  nand02 U1584 ( .Y(n3190), .A0(n3185), .A1(n3187) );
  nand02 U1585 ( .Y(n3191), .A0(n3186), .A1(n3187) );
  nand02 U1586 ( .Y(n3192), .A0(n3188), .A1(n3189) );
  inv01 U1587 ( .Y(n3182), .A(n3192) );
  nand02 U1588 ( .Y(n3193), .A0(n3190), .A1(n3191) );
  inv01 U1589 ( .Y(n3183), .A(n3193) );
  nand02 U1590 ( .Y(n7778), .A0(n3194), .A1(n3195) );
  inv01 U1591 ( .Y(n3196), .A(n7389) );
  inv01 U1592 ( .Y(n3197), .A(n7771) );
  inv01 U1593 ( .Y(n3198), .A(ARG1118_11_) );
  inv01 U1594 ( .Y(n3199), .A(r1_11_) );
  nand02 U1595 ( .Y(n3200), .A0(n3196), .A1(n3197) );
  nand02 U1596 ( .Y(n3201), .A0(n3196), .A1(n3198) );
  nand02 U1597 ( .Y(n3202), .A0(n3197), .A1(n3199) );
  nand02 U1598 ( .Y(n3203), .A0(n3198), .A1(n3199) );
  nand02 U1599 ( .Y(n3204), .A0(n3200), .A1(n3201) );
  inv01 U1600 ( .Y(n3194), .A(n3204) );
  nand02 U1601 ( .Y(n3205), .A0(n3202), .A1(n3203) );
  inv01 U1602 ( .Y(n3195), .A(n3205) );
  ao22 U1603 ( .Y(n3206), .A0(ARG1118_7_), .A1(n7771), .B0(r1_7_), .B1(n7389)
         );
  inv01 U1604 ( .Y(n3207), .A(n3206) );
  ao22 U1605 ( .Y(n3208), .A0(ARG1118_12_), .A1(n7771), .B0(r1_12_), .B1(n7389) );
  inv01 U1606 ( .Y(n3209), .A(n3208) );
  nand02 U1607 ( .Y(n7777), .A0(n3210), .A1(n3211) );
  inv01 U1608 ( .Y(n3212), .A(n7389) );
  inv01 U1609 ( .Y(n3213), .A(n7771) );
  inv01 U1610 ( .Y(n3214), .A(ARG1118_10_) );
  inv01 U1611 ( .Y(n3215), .A(r1_10_) );
  nand02 U1612 ( .Y(n3216), .A0(n3212), .A1(n3213) );
  nand02 U1613 ( .Y(n3217), .A0(n3212), .A1(n3214) );
  nand02 U1614 ( .Y(n3218), .A0(n3213), .A1(n3215) );
  nand02 U1615 ( .Y(n3219), .A0(n3214), .A1(n3215) );
  nand02 U1616 ( .Y(n3220), .A0(n3216), .A1(n3217) );
  inv01 U1617 ( .Y(n3210), .A(n3220) );
  nand02 U1618 ( .Y(n3221), .A0(n3218), .A1(n3219) );
  inv01 U1619 ( .Y(n3211), .A(n3221) );
  nand02 U1620 ( .Y(n7781), .A0(n3222), .A1(n3223) );
  inv01 U1621 ( .Y(n3224), .A(n7389) );
  inv01 U1622 ( .Y(n3225), .A(n7771) );
  inv01 U1623 ( .Y(n3226), .A(ARG1118_17_) );
  inv01 U1624 ( .Y(n3227), .A(r1_17_) );
  nand02 U1625 ( .Y(n3228), .A0(n3224), .A1(n3225) );
  nand02 U1626 ( .Y(n3229), .A0(n3224), .A1(n3226) );
  nand02 U1627 ( .Y(n3230), .A0(n3225), .A1(n3227) );
  nand02 U1628 ( .Y(n3231), .A0(n3226), .A1(n3227) );
  nand02 U1629 ( .Y(n3232), .A0(n3228), .A1(n3229) );
  inv01 U1630 ( .Y(n3222), .A(n3232) );
  nand02 U1631 ( .Y(n3233), .A0(n3230), .A1(n3231) );
  inv01 U1632 ( .Y(n3223), .A(n3233) );
  nand02 U1633 ( .Y(n7782), .A0(n3234), .A1(n3235) );
  inv01 U1634 ( .Y(n3236), .A(n7389) );
  inv01 U1635 ( .Y(n3237), .A(n7771) );
  inv01 U1636 ( .Y(n3238), .A(ARG1118_18_) );
  inv01 U1637 ( .Y(n3239), .A(r1_18_) );
  nand02 U1638 ( .Y(n3240), .A0(n3236), .A1(n3237) );
  nand02 U1639 ( .Y(n3241), .A0(n3236), .A1(n3238) );
  nand02 U1640 ( .Y(n3242), .A0(n3237), .A1(n3239) );
  nand02 U1641 ( .Y(n3243), .A0(n3238), .A1(n3239) );
  nand02 U1642 ( .Y(n3244), .A0(n3240), .A1(n3241) );
  inv01 U1643 ( .Y(n3234), .A(n3244) );
  nand02 U1644 ( .Y(n3245), .A0(n3242), .A1(n3243) );
  inv01 U1645 ( .Y(n3235), .A(n3245) );
  ao22 U1646 ( .Y(n3246), .A0(ARG1118_6_), .A1(n7771), .B0(r1_6_), .B1(n7389)
         );
  inv01 U1647 ( .Y(n3247), .A(n3246) );
  nand02 U1648 ( .Y(n7783), .A0(n3248), .A1(n3249) );
  inv01 U1649 ( .Y(n3250), .A(n7389) );
  inv01 U1650 ( .Y(n3251), .A(n7771) );
  inv01 U1651 ( .Y(n3252), .A(ARG1118_19_) );
  inv01 U1652 ( .Y(n3253), .A(r1_19_) );
  nand02 U1653 ( .Y(n3254), .A0(n3250), .A1(n3251) );
  nand02 U1654 ( .Y(n3255), .A0(n3250), .A1(n3252) );
  nand02 U1655 ( .Y(n3256), .A0(n3251), .A1(n3253) );
  nand02 U1656 ( .Y(n3257), .A0(n3252), .A1(n3253) );
  nand02 U1657 ( .Y(n3258), .A0(n3254), .A1(n3255) );
  inv01 U1658 ( .Y(n3248), .A(n3258) );
  nand02 U1659 ( .Y(n3259), .A0(n3256), .A1(n3257) );
  inv01 U1660 ( .Y(n3249), .A(n3259) );
  nand02 U1661 ( .Y(n7773), .A0(n3260), .A1(n3261) );
  inv01 U1662 ( .Y(n3262), .A(n7389) );
  inv01 U1663 ( .Y(n3263), .A(n7771) );
  inv01 U1664 ( .Y(n3264), .A(ARG1118_3_) );
  inv01 U1665 ( .Y(n3265), .A(r1_3_) );
  nand02 U1666 ( .Y(n3266), .A0(n3262), .A1(n3263) );
  nand02 U1667 ( .Y(n3267), .A0(n3262), .A1(n3264) );
  nand02 U1668 ( .Y(n3268), .A0(n3263), .A1(n3265) );
  nand02 U1669 ( .Y(n3269), .A0(n3264), .A1(n3265) );
  nand02 U1670 ( .Y(n3270), .A0(n3266), .A1(n3267) );
  inv01 U1671 ( .Y(n3260), .A(n3270) );
  nand02 U1672 ( .Y(n3271), .A0(n3268), .A1(n3269) );
  inv01 U1673 ( .Y(n3261), .A(n3271) );
  nand02 U1674 ( .Y(n7784), .A0(n3272), .A1(n3273) );
  inv01 U1675 ( .Y(n3274), .A(n7389) );
  inv01 U1676 ( .Y(n3275), .A(n7771) );
  inv01 U1677 ( .Y(n3276), .A(ARG1118_20_) );
  inv01 U1678 ( .Y(n3277), .A(r1_20_) );
  nand02 U1679 ( .Y(n3278), .A0(n3274), .A1(n3275) );
  nand02 U1680 ( .Y(n3279), .A0(n3274), .A1(n3276) );
  nand02 U1681 ( .Y(n3280), .A0(n3275), .A1(n3277) );
  nand02 U1682 ( .Y(n3281), .A0(n3276), .A1(n3277) );
  nand02 U1683 ( .Y(n3282), .A0(n3278), .A1(n3279) );
  inv01 U1684 ( .Y(n3272), .A(n3282) );
  nand02 U1685 ( .Y(n3283), .A0(n3280), .A1(n3281) );
  inv01 U1686 ( .Y(n3273), .A(n3283) );
  ao22 U1687 ( .Y(n3284), .A0(ARG1118_22_), .A1(n7771), .B0(r1_22_), .B1(n7389) );
  inv01 U1688 ( .Y(n3285), .A(n3284) );
  ao22 U1689 ( .Y(n3286), .A0(ARG1118_25_), .A1(n7771), .B0(r1_25_), .B1(n7389) );
  inv01 U1690 ( .Y(n3287), .A(n3286) );
  nand02 U1691 ( .Y(n7774), .A0(n3288), .A1(n3289) );
  inv01 U1692 ( .Y(n3290), .A(n7389) );
  inv01 U1693 ( .Y(n3291), .A(n7771) );
  inv01 U1694 ( .Y(n3292), .A(ARG1118_4_) );
  inv01 U1695 ( .Y(n3293), .A(r1_4_) );
  nand02 U1696 ( .Y(n3294), .A0(n3290), .A1(n3291) );
  nand02 U1697 ( .Y(n3295), .A0(n3290), .A1(n3292) );
  nand02 U1698 ( .Y(n3296), .A0(n3291), .A1(n3293) );
  nand02 U1699 ( .Y(n3297), .A0(n3292), .A1(n3293) );
  nand02 U1700 ( .Y(n3298), .A0(n3294), .A1(n3295) );
  inv01 U1701 ( .Y(n3288), .A(n3298) );
  nand02 U1702 ( .Y(n3299), .A0(n3296), .A1(n3297) );
  inv01 U1703 ( .Y(n3289), .A(n3299) );
  nand02 U1704 ( .Y(n7785), .A0(n3300), .A1(n3301) );
  inv01 U1705 ( .Y(n3302), .A(n7389) );
  inv01 U1706 ( .Y(n3303), .A(n7771) );
  inv01 U1707 ( .Y(n3304), .A(ARG1118_21_) );
  inv01 U1708 ( .Y(n3305), .A(r1_21_) );
  nand02 U1709 ( .Y(n3306), .A0(n3302), .A1(n3303) );
  nand02 U1710 ( .Y(n3307), .A0(n3302), .A1(n3304) );
  nand02 U1711 ( .Y(n3308), .A0(n3303), .A1(n3305) );
  nand02 U1712 ( .Y(n3309), .A0(n3304), .A1(n3305) );
  nand02 U1713 ( .Y(n3310), .A0(n3306), .A1(n3307) );
  inv01 U1714 ( .Y(n3300), .A(n3310) );
  nand02 U1715 ( .Y(n3311), .A0(n3308), .A1(n3309) );
  inv01 U1716 ( .Y(n3301), .A(n3311) );
  nand02 U1717 ( .Y(n7775), .A0(n3312), .A1(n3313) );
  inv01 U1718 ( .Y(n3314), .A(n7389) );
  inv01 U1719 ( .Y(n3315), .A(n7771) );
  inv01 U1720 ( .Y(n3316), .A(ARG1118_5_) );
  inv01 U1721 ( .Y(n3317), .A(r1_5_) );
  nand02 U1722 ( .Y(n3318), .A0(n3314), .A1(n3315) );
  nand02 U1723 ( .Y(n3319), .A0(n3314), .A1(n3316) );
  nand02 U1724 ( .Y(n3320), .A0(n3315), .A1(n3317) );
  nand02 U1725 ( .Y(n3321), .A0(n3316), .A1(n3317) );
  nand02 U1726 ( .Y(n3322), .A0(n3318), .A1(n3319) );
  inv01 U1727 ( .Y(n3312), .A(n3322) );
  nand02 U1728 ( .Y(n3323), .A0(n3320), .A1(n3321) );
  inv01 U1729 ( .Y(n3313), .A(n3323) );
  ao22 U1730 ( .Y(n3324), .A0(ARG1118_13_), .A1(n7771), .B0(r1_13_), .B1(n7389) );
  inv01 U1731 ( .Y(n3325), .A(n3324) );
  ao22 U1732 ( .Y(n3326), .A0(ARG1118_24_), .A1(n7771), .B0(r1_24_), .B1(n7389) );
  inv01 U1733 ( .Y(n3327), .A(n3326) );
  ao22 U1734 ( .Y(n3328), .A0(n7374), .A1(n7569), .B0(n7384), .B1(n7570) );
  inv01 U1735 ( .Y(n3329), .A(n3328) );
  xor2 U1736 ( .Y(n3330), .A0(s_rad_i_30_), .A1(n7766) );
  inv01 U1737 ( .Y(n3331), .A(n3330) );
  xor2 U1738 ( .Y(n3332), .A0(s_rad_i_1_), .A1(n7758) );
  inv01 U1739 ( .Y(n3333), .A(n3332) );
  ao22 U1740 ( .Y(n3334), .A0(n7384), .A1(n7569), .B0(n7374), .B1(n7587) );
  inv01 U1741 ( .Y(n3335), .A(n3334) );
  nand02 U1742 ( .Y(n7780), .A0(n3336), .A1(n3337) );
  inv01 U1743 ( .Y(n3338), .A(n7389) );
  inv01 U1744 ( .Y(n3339), .A(n7771) );
  inv01 U1745 ( .Y(n3340), .A(ARG1118_16_) );
  inv01 U1746 ( .Y(n3341), .A(r1_16_) );
  nand02 U1747 ( .Y(n3342), .A0(n3338), .A1(n3339) );
  nand02 U1748 ( .Y(n3343), .A0(n3338), .A1(n3340) );
  nand02 U1749 ( .Y(n3344), .A0(n3339), .A1(n3341) );
  nand02 U1750 ( .Y(n3345), .A0(n3340), .A1(n3341) );
  nand02 U1751 ( .Y(n3346), .A0(n3342), .A1(n3343) );
  inv01 U1752 ( .Y(n3336), .A(n3346) );
  nand02 U1753 ( .Y(n3347), .A0(n3344), .A1(n3345) );
  inv01 U1754 ( .Y(n3337), .A(n3347) );
  nand02 U1755 ( .Y(n7772), .A0(n3348), .A1(n3349) );
  inv01 U1756 ( .Y(n3350), .A(n7389) );
  inv01 U1757 ( .Y(n3351), .A(n7771) );
  inv01 U1758 ( .Y(n3352), .A(ARG1118_2_) );
  inv01 U1759 ( .Y(n3353), .A(r1_2_) );
  nand02 U1760 ( .Y(n3354), .A0(n3350), .A1(n3351) );
  nand02 U1761 ( .Y(n3355), .A0(n3350), .A1(n3352) );
  nand02 U1762 ( .Y(n3356), .A0(n3351), .A1(n3353) );
  nand02 U1763 ( .Y(n3357), .A0(n3352), .A1(n3353) );
  nand02 U1764 ( .Y(n3358), .A0(n3354), .A1(n3355) );
  inv01 U1765 ( .Y(n3348), .A(n3358) );
  nand02 U1766 ( .Y(n3359), .A0(n3356), .A1(n3357) );
  inv01 U1767 ( .Y(n3349), .A(n3359) );
  nand02 U1768 ( .Y(n7779), .A0(n3360), .A1(n3361) );
  inv01 U1769 ( .Y(n3362), .A(n7389) );
  inv01 U1770 ( .Y(n3363), .A(n7771) );
  inv01 U1771 ( .Y(n3364), .A(ARG1118_14_) );
  inv01 U1772 ( .Y(n3365), .A(r1_14_) );
  nand02 U1773 ( .Y(n3366), .A0(n3362), .A1(n3363) );
  nand02 U1774 ( .Y(n3367), .A0(n3362), .A1(n3364) );
  nand02 U1775 ( .Y(n3368), .A0(n3363), .A1(n3365) );
  nand02 U1776 ( .Y(n3369), .A0(n3364), .A1(n3365) );
  nand02 U1777 ( .Y(n3370), .A0(n3366), .A1(n3367) );
  inv01 U1778 ( .Y(n3360), .A(n3370) );
  nand02 U1779 ( .Y(n3371), .A0(n3368), .A1(n3369) );
  inv01 U1780 ( .Y(n3361), .A(n3371) );
  ao22 U1781 ( .Y(n3372), .A0(ARG1118_8_), .A1(n7771), .B0(r1_8_), .B1(n7389)
         );
  inv01 U1782 ( .Y(n3373), .A(n3372) );
  or02 U1783 ( .Y(n3374), .A0(n7429), .A1(n2803) );
  inv01 U1784 ( .Y(n3375), .A(n3374) );
  or02 U1785 ( .Y(n3376), .A0(n7429), .A1(n2790) );
  inv01 U1786 ( .Y(n3377), .A(n3376) );
  or02 U1787 ( .Y(n3378), .A0(n7429), .A1(n2791) );
  inv01 U1788 ( .Y(n3379), .A(n3378) );
  or02 U1789 ( .Y(n3380), .A0(n7429), .A1(n2800) );
  inv01 U1790 ( .Y(n3381), .A(n3380) );
  or02 U1791 ( .Y(n3382), .A0(n7429), .A1(n2808) );
  inv01 U1792 ( .Y(n3383), .A(n3382) );
  or02 U1793 ( .Y(n3384), .A0(n7429), .A1(n2784) );
  inv01 U1794 ( .Y(n3385), .A(n3384) );
  or02 U1795 ( .Y(n3386), .A0(n7429), .A1(n2794) );
  inv01 U1796 ( .Y(n3387), .A(n3386) );
  or02 U1797 ( .Y(n3388), .A0(n7429), .A1(n2785) );
  inv01 U1798 ( .Y(n3389), .A(n3388) );
  or02 U1799 ( .Y(n3390), .A0(n7429), .A1(n2804) );
  inv01 U1800 ( .Y(n3391), .A(n3390) );
  or02 U1801 ( .Y(n3392), .A0(n7427), .A1(n2788) );
  inv01 U1802 ( .Y(n3393), .A(n3392) );
  or02 U1803 ( .Y(n3394), .A0(n7427), .A1(n2807) );
  inv01 U1804 ( .Y(n3395), .A(n3394) );
  or02 U1805 ( .Y(n3396), .A0(n7427), .A1(n2786) );
  inv01 U1806 ( .Y(n3397), .A(n3396) );
  or02 U1807 ( .Y(n3398), .A0(n7427), .A1(n2789) );
  inv01 U1808 ( .Y(n3399), .A(n3398) );
  or02 U1809 ( .Y(n3400), .A0(n7427), .A1(n2793) );
  inv01 U1810 ( .Y(n3401), .A(n3400) );
  or02 U1811 ( .Y(n3402), .A0(n7427), .A1(n2792) );
  inv01 U1812 ( .Y(n3403), .A(n3402) );
  or02 U1813 ( .Y(n3404), .A0(n7427), .A1(n2802) );
  inv01 U1814 ( .Y(n3405), .A(n3404) );
  or02 U1815 ( .Y(n3406), .A0(n7427), .A1(n2797) );
  inv01 U1816 ( .Y(n3407), .A(n3406) );
  or02 U1817 ( .Y(n3408), .A0(n7427), .A1(n2795) );
  inv01 U1818 ( .Y(n3409), .A(n3408) );
  or02 U1819 ( .Y(n3410), .A0(n7455), .A1(n7432) );
  inv01 U1820 ( .Y(n3411), .A(n3410) );
  or02 U1821 ( .Y(n3412), .A0(n7428), .A1(n2806) );
  inv01 U1822 ( .Y(n3413), .A(n3412) );
  or02 U1823 ( .Y(n3414), .A0(n7428), .A1(n2796) );
  inv01 U1824 ( .Y(n3415), .A(n3414) );
  or02 U1825 ( .Y(n3416), .A0(n7428), .A1(n2805) );
  inv01 U1826 ( .Y(n3417), .A(n3416) );
  or02 U1827 ( .Y(n3418), .A0(n7428), .A1(n2787) );
  inv01 U1828 ( .Y(n3419), .A(n3418) );
  or02 U1829 ( .Y(n3420), .A0(n7428), .A1(n2799) );
  inv01 U1830 ( .Y(n3421), .A(n3420) );
  or02 U1831 ( .Y(n3422), .A0(n7428), .A1(n2798) );
  inv01 U1832 ( .Y(n3423), .A(n3422) );
  or02 U1833 ( .Y(n3424), .A0(n7428), .A1(n2801) );
  inv01 U1834 ( .Y(n3425), .A(n3424) );
  nand02 U1835 ( .Y(n7670), .A0(n3426), .A1(n3427) );
  inv01 U1836 ( .Y(n3428), .A(n7399) );
  inv01 U1837 ( .Y(n3429), .A(n7401) );
  inv01 U1838 ( .Y(n3430), .A(r0_25_) );
  inv01 U1839 ( .Y(n3431), .A(r0_26_) );
  nand02 U1840 ( .Y(n3432), .A0(n3428), .A1(n3429) );
  nand02 U1841 ( .Y(n3433), .A0(n3428), .A1(n3430) );
  nand02 U1842 ( .Y(n3434), .A0(n3429), .A1(n3431) );
  nand02 U1843 ( .Y(n3435), .A0(n3430), .A1(n3431) );
  nand02 U1844 ( .Y(n3436), .A0(n3432), .A1(n3433) );
  inv01 U1845 ( .Y(n3426), .A(n3436) );
  nand02 U1846 ( .Y(n3437), .A0(n3434), .A1(n3435) );
  inv01 U1847 ( .Y(n3427), .A(n3437) );
  nand02 U1848 ( .Y(n7650), .A0(n3438), .A1(n3439) );
  inv01 U1849 ( .Y(n3440), .A(n7398) );
  inv01 U1850 ( .Y(n3441), .A(n7401) );
  inv01 U1851 ( .Y(n3442), .A(r0_7_) );
  inv01 U1852 ( .Y(n3443), .A(r0_8_) );
  nand02 U1853 ( .Y(n3444), .A0(n3440), .A1(n3441) );
  nand02 U1854 ( .Y(n3445), .A0(n3440), .A1(n3442) );
  nand02 U1855 ( .Y(n3446), .A0(n3441), .A1(n3443) );
  nand02 U1856 ( .Y(n3447), .A0(n3442), .A1(n3443) );
  nand02 U1857 ( .Y(n3448), .A0(n3444), .A1(n3445) );
  inv01 U1858 ( .Y(n3438), .A(n3448) );
  nand02 U1859 ( .Y(n3449), .A0(n3446), .A1(n3447) );
  inv01 U1860 ( .Y(n3439), .A(n3449) );
  nand02 U1861 ( .Y(n7456), .A0(n3450), .A1(n3451) );
  inv01 U1862 ( .Y(n3452), .A(n7398) );
  inv01 U1863 ( .Y(n3453), .A(n7401) );
  inv01 U1864 ( .Y(n3454), .A(r0_50_) );
  inv01 U1865 ( .Y(n3455), .A(r0_51_) );
  nand02 U1866 ( .Y(n3456), .A0(n3452), .A1(n3453) );
  nand02 U1867 ( .Y(n3457), .A0(n3452), .A1(n3454) );
  nand02 U1868 ( .Y(n3458), .A0(n3453), .A1(n3455) );
  nand02 U1869 ( .Y(n3459), .A0(n3454), .A1(n3455) );
  nand02 U1870 ( .Y(n3460), .A0(n3456), .A1(n3457) );
  inv01 U1871 ( .Y(n3450), .A(n3460) );
  nand02 U1872 ( .Y(n3461), .A0(n3458), .A1(n3459) );
  inv01 U1873 ( .Y(n3451), .A(n3461) );
  ao22 U1874 ( .Y(n3462), .A0(r0_44_), .A1(n7401), .B0(r0_45_), .B1(n7400) );
  inv01 U1875 ( .Y(n3463), .A(n3462) );
  nand02 U1876 ( .Y(n7499), .A0(n3464), .A1(n3465) );
  inv01 U1877 ( .Y(n3466), .A(n7399) );
  inv01 U1878 ( .Y(n3467), .A(n7401) );
  inv01 U1879 ( .Y(n3468), .A(r0_43_) );
  inv01 U1880 ( .Y(n3469), .A(r0_44_) );
  nand02 U1881 ( .Y(n3470), .A0(n3466), .A1(n3467) );
  nand02 U1882 ( .Y(n3471), .A0(n3466), .A1(n3468) );
  nand02 U1883 ( .Y(n3472), .A0(n3467), .A1(n3469) );
  nand02 U1884 ( .Y(n3473), .A0(n3468), .A1(n3469) );
  nand02 U1885 ( .Y(n3474), .A0(n3470), .A1(n3471) );
  inv01 U1886 ( .Y(n3464), .A(n3474) );
  nand02 U1887 ( .Y(n3475), .A0(n3472), .A1(n3473) );
  inv01 U1888 ( .Y(n3465), .A(n3475) );
  nand02 U1889 ( .Y(n7564), .A0(n3476), .A1(n3477) );
  inv01 U1890 ( .Y(n3478), .A(n7398) );
  inv01 U1891 ( .Y(n3479), .A(n7401) );
  inv01 U1892 ( .Y(n3480), .A(r0_30_) );
  inv01 U1893 ( .Y(n3481), .A(r0_31_) );
  nand02 U1894 ( .Y(n3482), .A0(n3478), .A1(n3479) );
  nand02 U1895 ( .Y(n3483), .A0(n3478), .A1(n3480) );
  nand02 U1896 ( .Y(n3484), .A0(n3479), .A1(n3481) );
  nand02 U1897 ( .Y(n3485), .A0(n3480), .A1(n3481) );
  nand02 U1898 ( .Y(n3486), .A0(n3482), .A1(n3483) );
  inv01 U1899 ( .Y(n3476), .A(n3486) );
  nand02 U1900 ( .Y(n3487), .A0(n3484), .A1(n3485) );
  inv01 U1901 ( .Y(n3477), .A(n3487) );
  nand02 U1902 ( .Y(n7505), .A0(n3488), .A1(n3489) );
  inv01 U1903 ( .Y(n3490), .A(n7398) );
  inv01 U1904 ( .Y(n3491), .A(n7401) );
  inv01 U1905 ( .Y(n3492), .A(r0_42_) );
  inv01 U1906 ( .Y(n3493), .A(r0_43_) );
  nand02 U1907 ( .Y(n3494), .A0(n3490), .A1(n3491) );
  nand02 U1908 ( .Y(n3495), .A0(n3490), .A1(n3492) );
  nand02 U1909 ( .Y(n3496), .A0(n3491), .A1(n3493) );
  nand02 U1910 ( .Y(n3497), .A0(n3492), .A1(n3493) );
  nand02 U1911 ( .Y(n3498), .A0(n3494), .A1(n3495) );
  inv01 U1912 ( .Y(n3488), .A(n3498) );
  nand02 U1913 ( .Y(n3499), .A0(n3496), .A1(n3497) );
  inv01 U1914 ( .Y(n3489), .A(n3499) );
  ao22 U1915 ( .Y(n3500), .A0(r0_28_), .A1(n7401), .B0(r0_29_), .B1(n7400) );
  inv01 U1916 ( .Y(n3501), .A(n3500) );
  buf04 U1917 ( .Y(n7399), .A(n7396) );
  ao22 U1918 ( .Y(n3502), .A0(r0_32_), .A1(n7401), .B0(r0_33_), .B1(n7400) );
  inv01 U1919 ( .Y(n3503), .A(n3502) );
  nand02 U1920 ( .Y(n7583), .A0(n3504), .A1(n3505) );
  inv01 U1921 ( .Y(n3506), .A(n7398) );
  inv01 U1922 ( .Y(n3507), .A(n7401) );
  inv01 U1923 ( .Y(n3508), .A(r0_26_) );
  inv01 U1924 ( .Y(n3509), .A(r0_27_) );
  nand02 U1925 ( .Y(n3510), .A0(n3506), .A1(n3507) );
  nand02 U1926 ( .Y(n3511), .A0(n3506), .A1(n3508) );
  nand02 U1927 ( .Y(n3512), .A0(n3507), .A1(n3509) );
  nand02 U1928 ( .Y(n3513), .A0(n3508), .A1(n3509) );
  nand02 U1929 ( .Y(n3514), .A0(n3510), .A1(n3511) );
  inv01 U1930 ( .Y(n3504), .A(n3514) );
  nand02 U1931 ( .Y(n3515), .A0(n3512), .A1(n3513) );
  inv01 U1932 ( .Y(n3505), .A(n3515) );
  ao22 U1933 ( .Y(n3516), .A0(r0_18_), .A1(n7401), .B0(r0_19_), .B1(n7398) );
  inv01 U1934 ( .Y(n3517), .A(n3516) );
  nand02 U1935 ( .Y(n7637), .A0(n3518), .A1(n3519) );
  inv01 U1936 ( .Y(n3520), .A(n7399) );
  inv01 U1937 ( .Y(n3521), .A(n7401) );
  inv01 U1938 ( .Y(n3522), .A(r0_13_) );
  inv01 U1939 ( .Y(n3523), .A(r0_14_) );
  nand02 U1940 ( .Y(n3524), .A0(n3520), .A1(n3521) );
  nand02 U1941 ( .Y(n3525), .A0(n3520), .A1(n3522) );
  nand02 U1942 ( .Y(n3526), .A0(n3521), .A1(n3523) );
  nand02 U1943 ( .Y(n3527), .A0(n3522), .A1(n3523) );
  nand02 U1944 ( .Y(n3528), .A0(n3524), .A1(n3525) );
  inv01 U1945 ( .Y(n3518), .A(n3528) );
  nand02 U1946 ( .Y(n3529), .A0(n3526), .A1(n3527) );
  inv01 U1947 ( .Y(n3519), .A(n3529) );
  nand02 U1948 ( .Y(n7655), .A0(n3530), .A1(n3531) );
  inv01 U1949 ( .Y(n3532), .A(n7399) );
  inv01 U1950 ( .Y(n3533), .A(n7401) );
  inv01 U1951 ( .Y(n3534), .A(r0_11_) );
  inv01 U1952 ( .Y(n3535), .A(r0_12_) );
  nand02 U1953 ( .Y(n3536), .A0(n3532), .A1(n3533) );
  nand02 U1954 ( .Y(n3537), .A0(n3532), .A1(n3534) );
  nand02 U1955 ( .Y(n3538), .A0(n3533), .A1(n3535) );
  nand02 U1956 ( .Y(n3539), .A0(n3534), .A1(n3535) );
  nand02 U1957 ( .Y(n3540), .A0(n3536), .A1(n3537) );
  inv01 U1958 ( .Y(n3530), .A(n3540) );
  nand02 U1959 ( .Y(n3541), .A0(n3538), .A1(n3539) );
  inv01 U1960 ( .Y(n3531), .A(n3541) );
  ao22 U1961 ( .Y(n3542), .A0(r0_27_), .A1(n7401), .B0(r0_28_), .B1(n7399) );
  inv01 U1962 ( .Y(n3543), .A(n3542) );
  nand02 U1963 ( .Y(n7648), .A0(n3544), .A1(n3545) );
  inv01 U1964 ( .Y(n3546), .A(n7399) );
  inv01 U1965 ( .Y(n3547), .A(n7401) );
  inv01 U1966 ( .Y(n3548), .A(r0_8_) );
  inv01 U1967 ( .Y(n3549), .A(r0_9_) );
  nand02 U1968 ( .Y(n3550), .A0(n3546), .A1(n3547) );
  nand02 U1969 ( .Y(n3551), .A0(n3546), .A1(n3548) );
  nand02 U1970 ( .Y(n3552), .A0(n3547), .A1(n3549) );
  nand02 U1971 ( .Y(n3553), .A0(n3548), .A1(n3549) );
  nand02 U1972 ( .Y(n3554), .A0(n3550), .A1(n3551) );
  inv01 U1973 ( .Y(n3544), .A(n3554) );
  nand02 U1974 ( .Y(n3555), .A0(n3552), .A1(n3553) );
  inv01 U1975 ( .Y(n3545), .A(n3555) );
  ao22 U1976 ( .Y(n3556), .A0(r0_46_), .A1(n7401), .B0(r0_47_), .B1(n7398) );
  inv01 U1977 ( .Y(n3557), .A(n3556) );
  nand02 U1978 ( .Y(n7662), .A0(n3558), .A1(n3559) );
  inv01 U1979 ( .Y(n3560), .A(n7398) );
  inv01 U1980 ( .Y(n3561), .A(n7401) );
  inv01 U1981 ( .Y(n3562), .A(r0_9_) );
  inv01 U1982 ( .Y(n3563), .A(r0_10_) );
  nand02 U1983 ( .Y(n3564), .A0(n3560), .A1(n3561) );
  nand02 U1984 ( .Y(n3565), .A0(n3560), .A1(n3562) );
  nand02 U1985 ( .Y(n3566), .A0(n3561), .A1(n3563) );
  nand02 U1986 ( .Y(n3567), .A0(n3562), .A1(n3563) );
  nand02 U1987 ( .Y(n3568), .A0(n3564), .A1(n3565) );
  inv01 U1988 ( .Y(n3558), .A(n3568) );
  nand02 U1989 ( .Y(n3569), .A0(n3566), .A1(n3567) );
  inv01 U1990 ( .Y(n3559), .A(n3569) );
  ao22 U1991 ( .Y(n3570), .A0(r0_34_), .A1(n7401), .B0(r0_35_), .B1(n7398) );
  inv01 U1992 ( .Y(n3571), .A(n3570) );
  nand02 U1993 ( .Y(n7645), .A0(n3572), .A1(n3573) );
  inv01 U1994 ( .Y(n3574), .A(n7400) );
  inv01 U1995 ( .Y(n3575), .A(n7401) );
  inv01 U1996 ( .Y(n3576), .A(r0_12_) );
  inv01 U1997 ( .Y(n3577), .A(r0_13_) );
  nand02 U1998 ( .Y(n3578), .A0(n3574), .A1(n3575) );
  nand02 U1999 ( .Y(n3579), .A0(n3574), .A1(n3576) );
  nand02 U2000 ( .Y(n3580), .A0(n3575), .A1(n3577) );
  nand02 U2001 ( .Y(n3581), .A0(n3576), .A1(n3577) );
  nand02 U2002 ( .Y(n3582), .A0(n3578), .A1(n3579) );
  inv01 U2003 ( .Y(n3572), .A(n3582) );
  nand02 U2004 ( .Y(n3583), .A0(n3580), .A1(n3581) );
  inv01 U2005 ( .Y(n3573), .A(n3583) );
  nand02 U2006 ( .Y(n7542), .A0(n3584), .A1(n3585) );
  inv01 U2007 ( .Y(n3586), .A(n7399) );
  inv01 U2008 ( .Y(n3587), .A(n7401) );
  inv01 U2009 ( .Y(n3588), .A(r0_35_) );
  inv01 U2010 ( .Y(n3589), .A(r0_36_) );
  nand02 U2011 ( .Y(n3590), .A0(n3586), .A1(n3587) );
  nand02 U2012 ( .Y(n3591), .A0(n3586), .A1(n3588) );
  nand02 U2013 ( .Y(n3592), .A0(n3587), .A1(n3589) );
  nand02 U2014 ( .Y(n3593), .A0(n3588), .A1(n3589) );
  nand02 U2015 ( .Y(n3594), .A0(n3590), .A1(n3591) );
  inv01 U2016 ( .Y(n3584), .A(n3594) );
  nand02 U2017 ( .Y(n3595), .A0(n3592), .A1(n3593) );
  inv01 U2018 ( .Y(n3585), .A(n3595) );
  ao22 U2019 ( .Y(n3596), .A0(r0_23_), .A1(n7401), .B0(r0_24_), .B1(n7399) );
  inv01 U2020 ( .Y(n3597), .A(n3596) );
  nand02 U2021 ( .Y(n7560), .A0(n3598), .A1(n3599) );
  inv01 U2022 ( .Y(n3600), .A(n7399) );
  inv01 U2023 ( .Y(n3601), .A(n7401) );
  inv01 U2024 ( .Y(n3602), .A(r0_31_) );
  inv01 U2025 ( .Y(n3603), .A(r0_32_) );
  nand02 U2026 ( .Y(n3604), .A0(n3600), .A1(n3601) );
  nand02 U2027 ( .Y(n3605), .A0(n3600), .A1(n3602) );
  nand02 U2028 ( .Y(n3606), .A0(n3601), .A1(n3603) );
  nand02 U2029 ( .Y(n3607), .A0(n3602), .A1(n3603) );
  nand02 U2030 ( .Y(n3608), .A0(n3604), .A1(n3605) );
  inv01 U2031 ( .Y(n3598), .A(n3608) );
  nand02 U2032 ( .Y(n3609), .A0(n3606), .A1(n3607) );
  inv01 U2033 ( .Y(n3599), .A(n3609) );
  nand02 U2034 ( .Y(n7466), .A0(n3610), .A1(n3611) );
  inv01 U2035 ( .Y(n3612), .A(n7400) );
  inv01 U2036 ( .Y(n3613), .A(n7401) );
  inv01 U2037 ( .Y(n3614), .A(r0_48_) );
  inv01 U2038 ( .Y(n3615), .A(r0_49_) );
  nand02 U2039 ( .Y(n3616), .A0(n3612), .A1(n3613) );
  nand02 U2040 ( .Y(n3617), .A0(n3612), .A1(n3614) );
  nand02 U2041 ( .Y(n3618), .A0(n3613), .A1(n3615) );
  nand02 U2042 ( .Y(n3619), .A0(n3614), .A1(n3615) );
  nand02 U2043 ( .Y(n3620), .A0(n3616), .A1(n3617) );
  inv01 U2044 ( .Y(n3610), .A(n3620) );
  nand02 U2045 ( .Y(n3621), .A0(n3618), .A1(n3619) );
  inv01 U2046 ( .Y(n3611), .A(n3621) );
  nand02 U2047 ( .Y(n7661), .A0(n3622), .A1(n3623) );
  inv01 U2048 ( .Y(n3624), .A(n7399) );
  inv01 U2049 ( .Y(n3625), .A(n7401) );
  inv01 U2050 ( .Y(n3626), .A(r0_6_) );
  inv01 U2051 ( .Y(n3627), .A(r0_7_) );
  nand02 U2052 ( .Y(n3628), .A0(n3624), .A1(n3625) );
  nand02 U2053 ( .Y(n3629), .A0(n3624), .A1(n3626) );
  nand02 U2054 ( .Y(n3630), .A0(n3625), .A1(n3627) );
  nand02 U2055 ( .Y(n3631), .A0(n3626), .A1(n3627) );
  nand02 U2056 ( .Y(n3632), .A0(n3628), .A1(n3629) );
  inv01 U2057 ( .Y(n3622), .A(n3632) );
  nand02 U2058 ( .Y(n3633), .A0(n3630), .A1(n3631) );
  inv01 U2059 ( .Y(n3623), .A(n3633) );
  ao22 U2060 ( .Y(n3634), .A0(r0_20_), .A1(n7401), .B0(r0_21_), .B1(n7400) );
  inv01 U2061 ( .Y(n3635), .A(n3634) );
  ao22 U2062 ( .Y(n3636), .A0(r0_40_), .A1(n7401), .B0(r0_41_), .B1(n7400) );
  inv01 U2063 ( .Y(n3637), .A(n3636) );
  nand02 U2064 ( .Y(n7633), .A0(n3638), .A1(n3639) );
  inv01 U2065 ( .Y(n3640), .A(n7400) );
  inv01 U2066 ( .Y(n3641), .A(n7401) );
  inv01 U2067 ( .Y(n3642), .A(r0_14_) );
  inv01 U2068 ( .Y(n3643), .A(r0_15_) );
  nand02 U2069 ( .Y(n3644), .A0(n3640), .A1(n3641) );
  nand02 U2070 ( .Y(n3645), .A0(n3640), .A1(n3642) );
  nand02 U2071 ( .Y(n3646), .A0(n3641), .A1(n3643) );
  nand02 U2072 ( .Y(n3647), .A0(n3642), .A1(n3643) );
  nand02 U2073 ( .Y(n3648), .A0(n3644), .A1(n3645) );
  inv01 U2074 ( .Y(n3638), .A(n3648) );
  nand02 U2075 ( .Y(n3649), .A0(n3646), .A1(n3647) );
  inv01 U2076 ( .Y(n3639), .A(n3649) );
  nand02 U2077 ( .Y(n7673), .A0(n3650), .A1(n3651) );
  inv01 U2078 ( .Y(n3652), .A(n7399) );
  inv01 U2079 ( .Y(n3653), .A(n7401) );
  inv01 U2080 ( .Y(n3654), .A(r0_29_) );
  inv01 U2081 ( .Y(n3655), .A(r0_30_) );
  nand02 U2082 ( .Y(n3656), .A0(n3652), .A1(n3653) );
  nand02 U2083 ( .Y(n3657), .A0(n3652), .A1(n3654) );
  nand02 U2084 ( .Y(n3658), .A0(n3653), .A1(n3655) );
  nand02 U2085 ( .Y(n3659), .A0(n3654), .A1(n3655) );
  nand02 U2086 ( .Y(n3660), .A0(n3656), .A1(n3657) );
  inv01 U2087 ( .Y(n3650), .A(n3660) );
  nand02 U2088 ( .Y(n3661), .A0(n3658), .A1(n3659) );
  inv01 U2089 ( .Y(n3651), .A(n3661) );
  ao22 U2090 ( .Y(n3662), .A0(r0_37_), .A1(n7401), .B0(r0_38_), .B1(n7400) );
  inv01 U2091 ( .Y(n3663), .A(n3662) );
  nand02 U2092 ( .Y(n7475), .A0(n3664), .A1(n3665) );
  inv01 U2093 ( .Y(n3666), .A(n7399) );
  inv01 U2094 ( .Y(n3667), .A(n7401) );
  inv01 U2095 ( .Y(n3668), .A(r0_47_) );
  inv01 U2096 ( .Y(n3669), .A(r0_48_) );
  nand02 U2097 ( .Y(n3670), .A0(n3666), .A1(n3667) );
  nand02 U2098 ( .Y(n3671), .A0(n3666), .A1(n3668) );
  nand02 U2099 ( .Y(n3672), .A0(n3667), .A1(n3669) );
  nand02 U2100 ( .Y(n3673), .A0(n3668), .A1(n3669) );
  nand02 U2101 ( .Y(n3674), .A0(n3670), .A1(n3671) );
  inv01 U2102 ( .Y(n3664), .A(n3674) );
  nand02 U2103 ( .Y(n3675), .A0(n3672), .A1(n3673) );
  inv01 U2104 ( .Y(n3665), .A(n3675) );
  nand02 U2105 ( .Y(n7659), .A0(n3676), .A1(n3677) );
  inv01 U2106 ( .Y(n3678), .A(n7400) );
  inv01 U2107 ( .Y(n3679), .A(n7401) );
  inv01 U2108 ( .Y(n3680), .A(r0_2_) );
  inv01 U2109 ( .Y(n3681), .A(r0_3_) );
  nand02 U2110 ( .Y(n3682), .A0(n3678), .A1(n3679) );
  nand02 U2111 ( .Y(n3683), .A0(n3678), .A1(n3680) );
  nand02 U2112 ( .Y(n3684), .A0(n3679), .A1(n3681) );
  nand02 U2113 ( .Y(n3685), .A0(n3680), .A1(n3681) );
  nand02 U2114 ( .Y(n3686), .A0(n3682), .A1(n3683) );
  inv01 U2115 ( .Y(n3676), .A(n3686) );
  nand02 U2116 ( .Y(n3687), .A0(n3684), .A1(n3685) );
  inv01 U2117 ( .Y(n3677), .A(n3687) );
  nand02 U2118 ( .Y(n7657), .A0(n3688), .A1(n3689) );
  inv01 U2119 ( .Y(n3690), .A(n7398) );
  inv01 U2120 ( .Y(n3691), .A(n7401) );
  inv01 U2121 ( .Y(n3692), .A(r0_10_) );
  inv01 U2122 ( .Y(n3693), .A(r0_11_) );
  nand02 U2123 ( .Y(n3694), .A0(n3690), .A1(n3691) );
  nand02 U2124 ( .Y(n3695), .A0(n3690), .A1(n3692) );
  nand02 U2125 ( .Y(n3696), .A0(n3691), .A1(n3693) );
  nand02 U2126 ( .Y(n3697), .A0(n3692), .A1(n3693) );
  nand02 U2127 ( .Y(n3698), .A0(n3694), .A1(n3695) );
  inv01 U2128 ( .Y(n3688), .A(n3698) );
  nand02 U2129 ( .Y(n3699), .A0(n3696), .A1(n3697) );
  inv01 U2130 ( .Y(n3689), .A(n3699) );
  ao22 U2131 ( .Y(n3700), .A0(r0_19_), .A1(n7401), .B0(r0_20_), .B1(n7399) );
  inv01 U2132 ( .Y(n3701), .A(n3700) );
  inv01 U2133 ( .Y(n7675), .A(n3702) );
  nor02 U2134 ( .Y(n3703), .A0(n4048), .A1(n4049) );
  nor02 U2135 ( .Y(n3704), .A0(n7678), .A1(n7679) );
  nor02 U2136 ( .Y(n3702), .A0(n3703), .A1(n3704) );
  nand02 U2137 ( .Y(n7664), .A0(n3705), .A1(n3706) );
  inv01 U2138 ( .Y(n3707), .A(n7400) );
  inv01 U2139 ( .Y(n3708), .A(n7401) );
  inv01 U2140 ( .Y(n3709), .A(r0_5_) );
  inv01 U2141 ( .Y(n3710), .A(r0_6_) );
  nand02 U2142 ( .Y(n3711), .A0(n3707), .A1(n3708) );
  nand02 U2143 ( .Y(n3712), .A0(n3707), .A1(n3709) );
  nand02 U2144 ( .Y(n3713), .A0(n3708), .A1(n3710) );
  nand02 U2145 ( .Y(n3714), .A0(n3709), .A1(n3710) );
  nand02 U2146 ( .Y(n3715), .A0(n3711), .A1(n3712) );
  inv01 U2147 ( .Y(n3705), .A(n3715) );
  nand02 U2148 ( .Y(n3716), .A0(n3713), .A1(n3714) );
  inv01 U2149 ( .Y(n3706), .A(n3716) );
  nand02 U2150 ( .Y(n7672), .A0(n3717), .A1(n3718) );
  inv01 U2151 ( .Y(n3719), .A(n7400) );
  inv01 U2152 ( .Y(n3720), .A(n7401) );
  inv01 U2153 ( .Y(n3721), .A(r0_33_) );
  inv01 U2154 ( .Y(n3722), .A(r0_34_) );
  nand02 U2155 ( .Y(n3723), .A0(n3719), .A1(n3720) );
  nand02 U2156 ( .Y(n3724), .A0(n3719), .A1(n3721) );
  nand02 U2157 ( .Y(n3725), .A0(n3720), .A1(n3722) );
  nand02 U2158 ( .Y(n3726), .A0(n3721), .A1(n3722) );
  nand02 U2159 ( .Y(n3727), .A0(n3723), .A1(n3724) );
  inv01 U2160 ( .Y(n3717), .A(n3727) );
  nand02 U2161 ( .Y(n3728), .A0(n3725), .A1(n3726) );
  inv01 U2162 ( .Y(n3718), .A(n3728) );
  ao22 U2163 ( .Y(n3729), .A0(r0_38_), .A1(n7401), .B0(r0_39_), .B1(n7398) );
  inv01 U2164 ( .Y(n3730), .A(n3729) );
  nand02 U2165 ( .Y(n7671), .A0(n3731), .A1(n3732) );
  inv01 U2166 ( .Y(n3733), .A(n7398) );
  inv01 U2167 ( .Y(n3734), .A(n7401) );
  inv01 U2168 ( .Y(n3735), .A(r0_21_) );
  inv01 U2169 ( .Y(n3736), .A(r0_22_) );
  nand02 U2170 ( .Y(n3737), .A0(n3733), .A1(n3734) );
  nand02 U2171 ( .Y(n3738), .A0(n3733), .A1(n3735) );
  nand02 U2172 ( .Y(n3739), .A0(n3734), .A1(n3736) );
  nand02 U2173 ( .Y(n3740), .A0(n3735), .A1(n3736) );
  nand02 U2174 ( .Y(n3741), .A0(n3737), .A1(n3738) );
  inv01 U2175 ( .Y(n3731), .A(n3741) );
  nand02 U2176 ( .Y(n3742), .A0(n3739), .A1(n3740) );
  inv01 U2177 ( .Y(n3732), .A(n3742) );
  nand02 U2178 ( .Y(n7653), .A0(n3743), .A1(n3744) );
  inv01 U2179 ( .Y(n3745), .A(n7400) );
  inv01 U2180 ( .Y(n3746), .A(n7401) );
  inv01 U2181 ( .Y(n3747), .A(r0_3_) );
  inv01 U2182 ( .Y(n3748), .A(r0_4_) );
  nand02 U2183 ( .Y(n3749), .A0(n3745), .A1(n3746) );
  nand02 U2184 ( .Y(n3750), .A0(n3745), .A1(n3747) );
  nand02 U2185 ( .Y(n3751), .A0(n3746), .A1(n3748) );
  nand02 U2186 ( .Y(n3752), .A0(n3747), .A1(n3748) );
  nand02 U2187 ( .Y(n3753), .A0(n3749), .A1(n3750) );
  inv01 U2188 ( .Y(n3743), .A(n3753) );
  nand02 U2189 ( .Y(n3754), .A0(n3751), .A1(n3752) );
  inv01 U2190 ( .Y(n3744), .A(n3754) );
  ao22 U2191 ( .Y(n3755), .A0(r0_39_), .A1(n7401), .B0(r0_40_), .B1(n7399) );
  inv01 U2192 ( .Y(n3756), .A(n3755) );
  nand02 U2193 ( .Y(n7592), .A0(n3757), .A1(n3758) );
  inv01 U2194 ( .Y(n3759), .A(n7400) );
  inv01 U2195 ( .Y(n3760), .A(n7401) );
  inv01 U2196 ( .Y(n3761), .A(r0_24_) );
  inv01 U2197 ( .Y(n3762), .A(r0_25_) );
  nand02 U2198 ( .Y(n3763), .A0(n3759), .A1(n3760) );
  nand02 U2199 ( .Y(n3764), .A0(n3759), .A1(n3761) );
  nand02 U2200 ( .Y(n3765), .A0(n3760), .A1(n3762) );
  nand02 U2201 ( .Y(n3766), .A0(n3761), .A1(n3762) );
  nand02 U2202 ( .Y(n3767), .A0(n3763), .A1(n3764) );
  inv01 U2203 ( .Y(n3757), .A(n3767) );
  nand02 U2204 ( .Y(n3768), .A0(n3765), .A1(n3766) );
  inv01 U2205 ( .Y(n3758), .A(n3768) );
  nand02 U2206 ( .Y(n7536), .A0(n3769), .A1(n3770) );
  inv01 U2207 ( .Y(n3771), .A(n7400) );
  inv01 U2208 ( .Y(n3772), .A(n7401) );
  inv01 U2209 ( .Y(n3773), .A(r0_36_) );
  inv01 U2210 ( .Y(n3774), .A(r0_37_) );
  nand02 U2211 ( .Y(n3775), .A0(n3771), .A1(n3772) );
  nand02 U2212 ( .Y(n3776), .A0(n3771), .A1(n3773) );
  nand02 U2213 ( .Y(n3777), .A0(n3772), .A1(n3774) );
  nand02 U2214 ( .Y(n3778), .A0(n3773), .A1(n3774) );
  nand02 U2215 ( .Y(n3779), .A0(n3775), .A1(n3776) );
  inv01 U2216 ( .Y(n3769), .A(n3779) );
  nand02 U2217 ( .Y(n3780), .A0(n3777), .A1(n3778) );
  inv01 U2218 ( .Y(n3770), .A(n3780) );
  nand02 U2219 ( .Y(n7668), .A0(n3781), .A1(n3782) );
  inv01 U2220 ( .Y(n3783), .A(n7399) );
  inv01 U2221 ( .Y(n3784), .A(n7401) );
  inv01 U2222 ( .Y(n3785), .A(r0_45_) );
  inv01 U2223 ( .Y(n3786), .A(r0_46_) );
  nand02 U2224 ( .Y(n3787), .A0(n3783), .A1(n3784) );
  nand02 U2225 ( .Y(n3788), .A0(n3783), .A1(n3785) );
  nand02 U2226 ( .Y(n3789), .A0(n3784), .A1(n3786) );
  nand02 U2227 ( .Y(n3790), .A0(n3785), .A1(n3786) );
  nand02 U2228 ( .Y(n3791), .A0(n3787), .A1(n3788) );
  inv01 U2229 ( .Y(n3781), .A(n3791) );
  nand02 U2230 ( .Y(n3792), .A0(n3789), .A1(n3790) );
  inv01 U2231 ( .Y(n3782), .A(n3792) );
  ao22 U2232 ( .Y(n3793), .A0(r0_41_), .A1(n7401), .B0(r0_42_), .B1(n7398) );
  inv01 U2233 ( .Y(n3794), .A(n3793) );
  ao22 U2234 ( .Y(n3795), .A0(r0_17_), .A1(n7401), .B0(r0_18_), .B1(n7400) );
  inv01 U2235 ( .Y(n3796), .A(n3795) );
  ao22 U2236 ( .Y(n3797), .A0(r0_22_), .A1(n7401), .B0(r0_23_), .B1(n7398) );
  inv01 U2237 ( .Y(n3798), .A(n3797) );
  xor2 U2238 ( .Y(n3799), .A0(n6781), .A1(r1_2_51_) );
  inv01 U2239 ( .Y(n3800), .A(n3799) );
  nand02 U2240 ( .Y(n7626), .A0(n3801), .A1(n3802) );
  inv01 U2241 ( .Y(n3803), .A(n7399) );
  inv01 U2242 ( .Y(n3804), .A(n7401) );
  inv01 U2243 ( .Y(n3805), .A(r0_16_) );
  inv01 U2244 ( .Y(n3806), .A(r0_17_) );
  nand02 U2245 ( .Y(n3807), .A0(n3803), .A1(n3804) );
  nand02 U2246 ( .Y(n3808), .A0(n3803), .A1(n3805) );
  nand02 U2247 ( .Y(n3809), .A0(n3804), .A1(n3806) );
  nand02 U2248 ( .Y(n3810), .A0(n3805), .A1(n3806) );
  nand02 U2249 ( .Y(n3811), .A0(n3807), .A1(n3808) );
  inv01 U2250 ( .Y(n3801), .A(n3811) );
  nand02 U2251 ( .Y(n3812), .A0(n3809), .A1(n3810) );
  inv01 U2252 ( .Y(n3802), .A(n3812) );
  nand02 U2253 ( .Y(n7630), .A0(n3813), .A1(n3814) );
  inv01 U2254 ( .Y(n3815), .A(n7398) );
  inv01 U2255 ( .Y(n3816), .A(n7401) );
  inv01 U2256 ( .Y(n3817), .A(r0_15_) );
  inv01 U2257 ( .Y(n3818), .A(r0_16_) );
  nand02 U2258 ( .Y(n3819), .A0(n3815), .A1(n3816) );
  nand02 U2259 ( .Y(n3820), .A0(n3815), .A1(n3817) );
  nand02 U2260 ( .Y(n3821), .A0(n3816), .A1(n3818) );
  nand02 U2261 ( .Y(n3822), .A0(n3817), .A1(n3818) );
  nand02 U2262 ( .Y(n3823), .A0(n3819), .A1(n3820) );
  inv01 U2263 ( .Y(n3813), .A(n3823) );
  nand02 U2264 ( .Y(n3824), .A0(n3821), .A1(n3822) );
  inv01 U2265 ( .Y(n3814), .A(n3824) );
  nand02 U2266 ( .Y(n7643), .A0(n3825), .A1(n3826) );
  inv01 U2267 ( .Y(n3827), .A(n7398) );
  inv01 U2268 ( .Y(n3828), .A(n7401) );
  inv01 U2269 ( .Y(n3829), .A(r0_4_) );
  inv01 U2270 ( .Y(n3830), .A(r0_5_) );
  nand02 U2271 ( .Y(n3831), .A0(n3827), .A1(n3828) );
  nand02 U2272 ( .Y(n3832), .A0(n3827), .A1(n3829) );
  nand02 U2273 ( .Y(n3833), .A0(n3828), .A1(n3830) );
  nand02 U2274 ( .Y(n3834), .A0(n3829), .A1(n3830) );
  nand02 U2275 ( .Y(n3835), .A0(n3831), .A1(n3832) );
  inv01 U2276 ( .Y(n3825), .A(n3835) );
  nand02 U2277 ( .Y(n3836), .A0(n3833), .A1(n3834) );
  inv01 U2278 ( .Y(n3826), .A(n3836) );
  ao22 U2279 ( .Y(n3837), .A0(r0_49_), .A1(n7401), .B0(r0_50_), .B1(n7398) );
  inv01 U2280 ( .Y(n3838), .A(n3837) );
  or02 U2281 ( .Y(n3839), .A0(n7419), .A1(n1847) );
  inv01 U2282 ( .Y(n3840), .A(n3839) );
  or02 U2283 ( .Y(n3841), .A0(n7419), .A1(n1929) );
  inv01 U2284 ( .Y(n3842), .A(n3841) );
  or02 U2285 ( .Y(n3843), .A0(n7419), .A1(n1832) );
  inv01 U2286 ( .Y(n3844), .A(n3843) );
  or02 U2287 ( .Y(n3845), .A0(n7419), .A1(n1874) );
  inv01 U2288 ( .Y(n3846), .A(n3845) );
  or02 U2289 ( .Y(n3847), .A0(n7419), .A1(n1863) );
  inv01 U2290 ( .Y(n3848), .A(n3847) );
  or02 U2291 ( .Y(n3849), .A0(n7421), .A1(n1878) );
  inv01 U2292 ( .Y(n3850), .A(n3849) );
  or02 U2293 ( .Y(n3851), .A0(n7421), .A1(n1870) );
  inv01 U2294 ( .Y(n3852), .A(n3851) );
  or02 U2295 ( .Y(n3853), .A0(n7421), .A1(n1904) );
  inv01 U2296 ( .Y(n3854), .A(n3853) );
  or02 U2297 ( .Y(n3855), .A0(n7419), .A1(n1898) );
  inv01 U2298 ( .Y(n3856), .A(n3855) );
  or02 U2299 ( .Y(n3857), .A0(n7419), .A1(n1877) );
  inv01 U2300 ( .Y(n3858), .A(n3857) );
  or02 U2301 ( .Y(n3859), .A0(n7419), .A1(n1852) );
  inv01 U2302 ( .Y(n3860), .A(n3859) );
  or02 U2303 ( .Y(n3861), .A0(n7421), .A1(n1908) );
  inv01 U2304 ( .Y(n3862), .A(n3861) );
  or02 U2305 ( .Y(n3863), .A0(n7421), .A1(n1901) );
  inv01 U2306 ( .Y(n3864), .A(n3863) );
  or02 U2307 ( .Y(n3865), .A0(n7421), .A1(n1867) );
  inv01 U2308 ( .Y(n3866), .A(n3865) );
  or02 U2309 ( .Y(n3867), .A0(n7421), .A1(n1899) );
  inv01 U2310 ( .Y(n3868), .A(n3867) );
  or02 U2311 ( .Y(n3869), .A0(n7419), .A1(n1923) );
  inv01 U2312 ( .Y(n3870), .A(n3869) );
  or02 U2313 ( .Y(n3871), .A0(n7419), .A1(n1926) );
  inv01 U2314 ( .Y(n3872), .A(n3871) );
  or02 U2315 ( .Y(n3873), .A0(n7419), .A1(n1837) );
  inv01 U2316 ( .Y(n3874), .A(n3873) );
  or02 U2317 ( .Y(n3875), .A0(n7421), .A1(n1919) );
  inv01 U2318 ( .Y(n3876), .A(n3875) );
  or02 U2319 ( .Y(n3877), .A0(n7421), .A1(n1893) );
  inv01 U2320 ( .Y(n3878), .A(n3877) );
  or02 U2321 ( .Y(n3879), .A0(n7421), .A1(n1927) );
  inv01 U2322 ( .Y(n3880), .A(n3879) );
  or02 U2323 ( .Y(n3881), .A0(n7421), .A1(n1896) );
  inv01 U2324 ( .Y(n3882), .A(n3881) );
  or02 U2325 ( .Y(n3883), .A0(n7419), .A1(n1866) );
  inv01 U2326 ( .Y(n3884), .A(n3883) );
  or02 U2327 ( .Y(n3885), .A0(n7419), .A1(n1840) );
  inv01 U2328 ( .Y(n3886), .A(n3885) );
  or02 U2329 ( .Y(n3887), .A0(n7419), .A1(n1864) );
  inv01 U2330 ( .Y(n3888), .A(n3887) );
  or02 U2331 ( .Y(n3889), .A0(n7419), .A1(n1861) );
  inv01 U2332 ( .Y(n3890), .A(n3889) );
  or02 U2333 ( .Y(n3891), .A0(n7421), .A1(n1875) );
  inv01 U2334 ( .Y(n3892), .A(n3891) );
  or02 U2335 ( .Y(n3893), .A0(n7421), .A1(n1883) );
  inv01 U2336 ( .Y(n3894), .A(n3893) );
  or02 U2337 ( .Y(n3895), .A0(n7421), .A1(n2730) );
  inv01 U2338 ( .Y(n3896), .A(n3895) );
  or02 U2339 ( .Y(n3897), .A0(n7419), .A1(n1888) );
  inv01 U2340 ( .Y(n3898), .A(n3897) );
  or02 U2341 ( .Y(n3899), .A0(n7419), .A1(n1869) );
  inv01 U2342 ( .Y(n3900), .A(n3899) );
  or02 U2343 ( .Y(n3901), .A0(n7419), .A1(n1918) );
  inv01 U2344 ( .Y(n3902), .A(n3901) );
  or02 U2345 ( .Y(n3903), .A0(n7419), .A1(n1915) );
  inv01 U2346 ( .Y(n3904), .A(n3903) );
  or02 U2347 ( .Y(n3905), .A0(n7421), .A1(n1834) );
  inv01 U2348 ( .Y(n3906), .A(n3905) );
  or02 U2349 ( .Y(n3907), .A0(n7421), .A1(n1916) );
  inv01 U2350 ( .Y(n3908), .A(n3907) );
  or02 U2351 ( .Y(n3909), .A0(n7421), .A1(n1845) );
  inv01 U2352 ( .Y(n3910), .A(n3909) );
  or02 U2353 ( .Y(n3911), .A0(n7419), .A1(n1850) );
  inv01 U2354 ( .Y(n3912), .A(n3911) );
  or02 U2355 ( .Y(n3913), .A0(n7419), .A1(n1844) );
  inv01 U2356 ( .Y(n3914), .A(n3913) );
  or02 U2357 ( .Y(n3915), .A0(n7419), .A1(n1912) );
  inv01 U2358 ( .Y(n3916), .A(n3915) );
  or02 U2359 ( .Y(n3917), .A0(n7419), .A1(n1872) );
  inv01 U2360 ( .Y(n3918), .A(n3917) );
  or02 U2361 ( .Y(n3919), .A0(n7421), .A1(n1842) );
  inv01 U2362 ( .Y(n3920), .A(n3919) );
  or02 U2363 ( .Y(n3921), .A0(n7421), .A1(n1859) );
  inv01 U2364 ( .Y(n3922), .A(n3921) );
  or02 U2365 ( .Y(n3923), .A0(n7421), .A1(n1882) );
  inv01 U2366 ( .Y(n3924), .A(n3923) );
  or02 U2367 ( .Y(n3925), .A0(n7421), .A1(n1913) );
  inv01 U2368 ( .Y(n3926), .A(n3925) );
  or02 U2369 ( .Y(n3927), .A0(n7419), .A1(n1895) );
  inv01 U2370 ( .Y(n3928), .A(n3927) );
  or02 U2371 ( .Y(n3929), .A0(n7419), .A1(n1858) );
  inv01 U2372 ( .Y(n3930), .A(n3929) );
  or02 U2373 ( .Y(n3931), .A0(n7419), .A1(n1903) );
  inv01 U2374 ( .Y(n3932), .A(n3931) );
  or02 U2375 ( .Y(n3933), .A0(n7419), .A1(n1885) );
  inv01 U2376 ( .Y(n3934), .A(n3933) );
  or02 U2377 ( .Y(n3935), .A0(n7420), .A1(n1909) );
  inv01 U2378 ( .Y(n3936), .A(n3935) );
  or02 U2379 ( .Y(n3937), .A0(n7421), .A1(n1848) );
  inv01 U2380 ( .Y(n3938), .A(n3937) );
  or02 U2381 ( .Y(n3939), .A0(n7421), .A1(n1881) );
  inv01 U2382 ( .Y(n3940), .A(n3939) );
  or02 U2383 ( .Y(n3941), .A0(n7421), .A1(n1889) );
  inv01 U2384 ( .Y(n3942), .A(n3941) );
  or02 U2385 ( .Y(n3943), .A0(n7419), .A1(n1892) );
  inv01 U2386 ( .Y(n3944), .A(n3943) );
  or02 U2387 ( .Y(n3945), .A0(n7419), .A1(n1835) );
  inv01 U2388 ( .Y(n3946), .A(n3945) );
  or02 U2389 ( .Y(n3947), .A0(n7419), .A1(n1907) );
  inv01 U2390 ( .Y(n3948), .A(n3947) );
  or02 U2391 ( .Y(n3949), .A0(n7419), .A1(n1891) );
  inv01 U2392 ( .Y(n3950), .A(n3949) );
  or02 U2393 ( .Y(n3951), .A0(n7421), .A1(n1853) );
  inv01 U2394 ( .Y(n3952), .A(n3951) );
  or02 U2395 ( .Y(n3953), .A0(n7421), .A1(n1851) );
  inv01 U2396 ( .Y(n3954), .A(n3953) );
  or02 U2397 ( .Y(n3955), .A0(n7421), .A1(n1856) );
  inv01 U2398 ( .Y(n3956), .A(n3955) );
  or02 U2399 ( .Y(n3957), .A0(n7421), .A1(n1921) );
  inv01 U2400 ( .Y(n3958), .A(n3957) );
  or02 U2401 ( .Y(n3959), .A0(n7420), .A1(n1839) );
  inv01 U2402 ( .Y(n3960), .A(n3959) );
  or02 U2403 ( .Y(n3961), .A0(n7420), .A1(n1894) );
  inv01 U2404 ( .Y(n3962), .A(n3961) );
  or02 U2405 ( .Y(n3963), .A0(n7420), .A1(n1902) );
  inv01 U2406 ( .Y(n3964), .A(n3963) );
  or02 U2407 ( .Y(n3965), .A0(n7420), .A1(n2731) );
  inv01 U2408 ( .Y(n3966), .A(n3965) );
  or02 U2409 ( .Y(n3967), .A0(n7419), .A1(n1846) );
  inv01 U2410 ( .Y(n3968), .A(n3967) );
  or02 U2411 ( .Y(n3969), .A0(n7419), .A1(n1855) );
  inv01 U2412 ( .Y(n3970), .A(n3969) );
  or02 U2413 ( .Y(n3971), .A0(n7419), .A1(n1884) );
  inv01 U2414 ( .Y(n3972), .A(n3971) );
  or02 U2415 ( .Y(n3973), .A0(n7419), .A1(n1910) );
  inv01 U2416 ( .Y(n3974), .A(n3973) );
  or02 U2417 ( .Y(n3975), .A0(n7421), .A1(n1924) );
  inv01 U2418 ( .Y(n3976), .A(n3975) );
  or02 U2419 ( .Y(n3977), .A0(n7421), .A1(n1886) );
  inv01 U2420 ( .Y(n3978), .A(n3977) );
  or02 U2421 ( .Y(n3979), .A0(n7421), .A1(n1930) );
  inv01 U2422 ( .Y(n3980), .A(n3979) );
  or02 U2423 ( .Y(n3981), .A0(n7421), .A1(n1865) );
  inv01 U2424 ( .Y(n3982), .A(n3981) );
  or02 U2425 ( .Y(n3983), .A0(n7420), .A1(n1836) );
  inv01 U2426 ( .Y(n3984), .A(n3983) );
  or02 U2427 ( .Y(n3985), .A0(n7420), .A1(n1860) );
  inv01 U2428 ( .Y(n3986), .A(n3985) );
  or02 U2429 ( .Y(n3987), .A0(n7420), .A1(n1925) );
  inv01 U2430 ( .Y(n3988), .A(n3987) );
  or02 U2431 ( .Y(n3989), .A0(n7420), .A1(n1922) );
  inv01 U2432 ( .Y(n3990), .A(n3989) );
  or02 U2433 ( .Y(n3991), .A0(n7420), .A1(n1911) );
  inv01 U2434 ( .Y(n3992), .A(n3991) );
  or02 U2435 ( .Y(n3993), .A0(n7420), .A1(n1897) );
  inv01 U2436 ( .Y(n3994), .A(n3993) );
  or02 U2437 ( .Y(n3995), .A0(n7420), .A1(n1914) );
  inv01 U2438 ( .Y(n3996), .A(n3995) );
  or02 U2439 ( .Y(n3997), .A0(n7420), .A1(n1838) );
  inv01 U2440 ( .Y(n3998), .A(n3997) );
  or02 U2441 ( .Y(n3999), .A0(n7420), .A1(n1890) );
  inv01 U2442 ( .Y(n4000), .A(n3999) );
  or02 U2443 ( .Y(n4001), .A0(n7420), .A1(n1833) );
  inv01 U2444 ( .Y(n4002), .A(n4001) );
  or02 U2445 ( .Y(n4003), .A0(n7420), .A1(n1843) );
  inv01 U2446 ( .Y(n4004), .A(n4003) );
  or02 U2447 ( .Y(n4005), .A0(n7420), .A1(n1841) );
  inv01 U2448 ( .Y(n4006), .A(n4005) );
  or02 U2449 ( .Y(n4007), .A0(n7420), .A1(n1871) );
  inv01 U2450 ( .Y(n4008), .A(n4007) );
  or02 U2451 ( .Y(n4009), .A0(n7420), .A1(n1887) );
  inv01 U2452 ( .Y(n4010), .A(n4009) );
  or02 U2453 ( .Y(n4011), .A0(n7420), .A1(n1917) );
  inv01 U2454 ( .Y(n4012), .A(n4011) );
  or02 U2455 ( .Y(n4013), .A0(n7420), .A1(n1857) );
  inv01 U2456 ( .Y(n4014), .A(n4013) );
  or02 U2457 ( .Y(n4015), .A0(n7420), .A1(n1876) );
  inv01 U2458 ( .Y(n4016), .A(n4015) );
  or02 U2459 ( .Y(n4017), .A0(n7420), .A1(n1900) );
  inv01 U2460 ( .Y(n4018), .A(n4017) );
  or02 U2461 ( .Y(n4019), .A0(n7420), .A1(n1868) );
  inv01 U2462 ( .Y(n4020), .A(n4019) );
  or02 U2463 ( .Y(n4021), .A0(n7420), .A1(n1920) );
  inv01 U2464 ( .Y(n4022), .A(n4021) );
  or02 U2465 ( .Y(n4023), .A0(n7420), .A1(n1928) );
  inv01 U2466 ( .Y(n4024), .A(n4023) );
  or02 U2467 ( .Y(n4025), .A0(n7420), .A1(n1862) );
  inv01 U2468 ( .Y(n4026), .A(n4025) );
  or02 U2469 ( .Y(n4027), .A0(n7420), .A1(n1873) );
  inv01 U2470 ( .Y(n4028), .A(n4027) );
  or02 U2471 ( .Y(n4029), .A0(n7420), .A1(n1905) );
  inv01 U2472 ( .Y(n4030), .A(n4029) );
  or02 U2473 ( .Y(n4031), .A0(n7420), .A1(n1854) );
  inv01 U2474 ( .Y(n4032), .A(n4031) );
  or02 U2475 ( .Y(n4033), .A0(n7420), .A1(n1849) );
  inv01 U2476 ( .Y(n4034), .A(n4033) );
  or02 U2477 ( .Y(n4035), .A0(n7420), .A1(n1880) );
  inv01 U2478 ( .Y(n4036), .A(n4035) );
  or02 U2479 ( .Y(n4037), .A0(n7420), .A1(n1879) );
  inv01 U2480 ( .Y(n4038), .A(n4037) );
  nand02 U2481 ( .Y(n7638), .A0(n4039), .A1(n4040) );
  inv01 U2482 ( .Y(n4041), .A(n7442) );
  inv01 U2483 ( .Y(n4042), .A(n7640) );
  inv01 U2484 ( .Y(n4043), .A(n7366) );
  inv01 U2485 ( .Y(n4044), .A(n7639) );
  nand02 U2486 ( .Y(n4039), .A0(n4041), .A1(n4042) );
  nand02 U2487 ( .Y(n4040), .A0(n4043), .A1(n4044) );
  inv01 U2488 ( .Y(n7669), .A(n4045) );
  nor02 U2489 ( .Y(n4046), .A0(n7640), .A1(n7566) );
  nor02 U2490 ( .Y(n4047), .A0(n7639), .A1(n7586) );
  nor02 U2491 ( .Y(n4045), .A0(n4046), .A1(n4047) );
  buf02 U2492 ( .Y(n4048), .A(n7680) );
  buf02 U2493 ( .Y(n4049), .A(n7681) );
  xor2 U2494 ( .Y(n4050), .A0(n6254), .A1(n____return1382_8_) );
  inv01 U2495 ( .Y(n4051), .A(n4050) );
  xor2 U2496 ( .Y(n4052), .A0(s_rad_i_3_), .A1(n____return1382_3_) );
  inv01 U2497 ( .Y(n4053), .A(n4052) );
  xor2 U2498 ( .Y(n4054), .A0(s_rad_i_3_), .A1(r1_2_3_) );
  inv01 U2499 ( .Y(n4055), .A(n4054) );
  inv08 U2500 ( .Y(n7387), .A(n7386) );
  xor2 U2501 ( .Y(n4056), .A0(s_rad_i_16_), .A1(r1_2_16_) );
  inv01 U2502 ( .Y(n4057), .A(n4056) );
  xor2 U2503 ( .Y(n4058), .A0(s_rad_i_6_), .A1(n____return1382_6_) );
  inv01 U2504 ( .Y(n4059), .A(n4058) );
  xor2 U2505 ( .Y(n4060), .A0(s_rad_i_16_), .A1(n____return1382_16_) );
  inv01 U2506 ( .Y(n4061), .A(n4060) );
  xor2 U2507 ( .Y(n4062), .A0(s_rad_i_28_), .A1(r1_2_28_) );
  inv01 U2508 ( .Y(n4063), .A(n4062) );
  xor2 U2509 ( .Y(n4064), .A0(s_rad_i_28_), .A1(n____return1382_28_) );
  inv01 U2510 ( .Y(n4065), .A(n4064) );
  xor2 U2511 ( .Y(n4066), .A0(s_rad_i_41_), .A1(r1_2_41_) );
  inv01 U2512 ( .Y(n4067), .A(n4066) );
  xor2 U2513 ( .Y(n4068), .A0(s_rad_i_41_), .A1(n____return1382_41_) );
  inv01 U2514 ( .Y(n4069), .A(n4068) );
  xor2 U2515 ( .Y(n4070), .A0(s_rad_i_6_), .A1(r1_2_6_) );
  inv01 U2516 ( .Y(n4071), .A(n4070) );
  xor2 U2517 ( .Y(n4072), .A0(s_rad_i_2_), .A1(n____return1382_2_) );
  inv01 U2518 ( .Y(n4073), .A(n4072) );
  xor2 U2519 ( .Y(n4074), .A0(s_rad_i_2_), .A1(r1_2_2_) );
  inv01 U2520 ( .Y(n4075), .A(n4074) );
  xor2 U2521 ( .Y(n4076), .A0(s_rad_i_18_), .A1(r1_2_18_) );
  inv01 U2522 ( .Y(n4077), .A(n4076) );
  xor2 U2523 ( .Y(n4078), .A0(s_rad_i_18_), .A1(n____return1382_18_) );
  inv01 U2524 ( .Y(n4079), .A(n4078) );
  xor2 U2525 ( .Y(n4080), .A0(n6263), .A1(r1_2_24_) );
  inv01 U2526 ( .Y(n4081), .A(n4080) );
  xor2 U2527 ( .Y(n4082), .A0(n6258), .A1(n____return1382_12_) );
  inv01 U2528 ( .Y(n4083), .A(n4082) );
  xor2 U2529 ( .Y(n4084), .A0(n6262), .A1(n____return1382_24_) );
  inv01 U2530 ( .Y(n4085), .A(n4084) );
  xor2 U2531 ( .Y(n4086), .A0(n6259), .A1(r1_2_12_) );
  inv01 U2532 ( .Y(n4087), .A(n4086) );
  xor2 U2533 ( .Y(n4088), .A0(s_rad_i_29_), .A1(n____return1382_29_) );
  inv01 U2534 ( .Y(n4089), .A(n4088) );
  xor2 U2535 ( .Y(n4090), .A0(s_rad_i_7_), .A1(n____return1382_7_) );
  inv01 U2536 ( .Y(n4091), .A(n4090) );
  xor2 U2537 ( .Y(n4092), .A0(s_rad_i_17_), .A1(n____return1382_17_) );
  inv01 U2538 ( .Y(n4093), .A(n4092) );
  xor2 U2539 ( .Y(n4094), .A0(s_rad_i_29_), .A1(r1_2_29_) );
  inv01 U2540 ( .Y(n4095), .A(n4094) );
  xor2 U2541 ( .Y(n4096), .A0(s_rad_i_17_), .A1(r1_2_17_) );
  inv01 U2542 ( .Y(n4097), .A(n4096) );
  xor2 U2543 ( .Y(n4098), .A0(s_rad_i_5_), .A1(r1_2_5_) );
  inv01 U2544 ( .Y(n4099), .A(n4098) );
  xor2 U2545 ( .Y(n4100), .A0(s_rad_i_40_), .A1(n____return1382_40_) );
  inv01 U2546 ( .Y(n4101), .A(n4100) );
  xor2 U2547 ( .Y(n4102), .A0(s_rad_i_40_), .A1(r1_2_40_) );
  inv01 U2548 ( .Y(n4103), .A(n4102) );
  xor2 U2549 ( .Y(n4104), .A0(s_rad_i_36_), .A1(n____return1382_36_) );
  inv01 U2550 ( .Y(n4105), .A(n4104) );
  xor2 U2551 ( .Y(n4106), .A0(s_rad_i_48_), .A1(n____return1382_48_) );
  inv01 U2552 ( .Y(n4107), .A(n4106) );
  xor2 U2553 ( .Y(n4108), .A0(s_rad_i_36_), .A1(r1_2_36_) );
  inv01 U2554 ( .Y(n4109), .A(n4108) );
  xor2 U2555 ( .Y(n4110), .A0(s_rad_i_48_), .A1(r1_2_48_) );
  inv01 U2556 ( .Y(n4111), .A(n4110) );
  xor2 U2557 ( .Y(n4112), .A0(s_rad_i_11_), .A1(n____return1382_11_) );
  inv01 U2558 ( .Y(n4113), .A(n4112) );
  xor2 U2559 ( .Y(n4114), .A0(s_rad_i_35_), .A1(n____return1382_35_) );
  inv01 U2560 ( .Y(n4115), .A(n4114) );
  xor2 U2561 ( .Y(n4116), .A0(s_rad_i_23_), .A1(r1_2_23_) );
  inv01 U2562 ( .Y(n4117), .A(n4116) );
  xor2 U2563 ( .Y(n4118), .A0(s_rad_i_47_), .A1(n____return1382_47_) );
  inv01 U2564 ( .Y(n4119), .A(n4118) );
  xor2 U2565 ( .Y(n4120), .A0(s_rad_i_35_), .A1(r1_2_35_) );
  inv01 U2566 ( .Y(n4121), .A(n4120) );
  xor2 U2567 ( .Y(n4122), .A0(s_rad_i_11_), .A1(r1_2_11_) );
  inv01 U2568 ( .Y(n4123), .A(n4122) );
  xor2 U2569 ( .Y(n4124), .A0(s_rad_i_47_), .A1(r1_2_47_) );
  inv01 U2570 ( .Y(n4125), .A(n4124) );
  xor2 U2571 ( .Y(n4126), .A0(s_rad_i_23_), .A1(n____return1382_23_) );
  inv01 U2572 ( .Y(n4127), .A(n4126) );
  xor2 U2573 ( .Y(n4128), .A0(s_rad_i_10_), .A1(n____return1382_10_) );
  inv01 U2574 ( .Y(n4129), .A(n4128) );
  xor2 U2575 ( .Y(n4130), .A0(s_rad_i_10_), .A1(r1_2_10_) );
  inv01 U2576 ( .Y(n4131), .A(n4130) );
  xor2 U2577 ( .Y(n4132), .A0(s_rad_i_46_), .A1(n____return1382_46_) );
  inv01 U2578 ( .Y(n4133), .A(n4132) );
  xor2 U2579 ( .Y(n4134), .A0(s_rad_i_46_), .A1(r1_2_46_) );
  inv01 U2580 ( .Y(n4135), .A(n4134) );
  xor2 U2581 ( .Y(n4136), .A0(s_rad_i_34_), .A1(n____return1382_34_) );
  inv01 U2582 ( .Y(n4137), .A(n4136) );
  xor2 U2583 ( .Y(n4138), .A0(s_rad_i_22_), .A1(n____return1382_22_) );
  inv01 U2584 ( .Y(n4139), .A(n4138) );
  xor2 U2585 ( .Y(n4140), .A0(s_rad_i_34_), .A1(r1_2_34_) );
  inv01 U2586 ( .Y(n4141), .A(n4140) );
  xor2 U2587 ( .Y(n4142), .A0(s_rad_i_22_), .A1(r1_2_22_) );
  inv01 U2588 ( .Y(n4143), .A(n4142) );
  inv02 U2589 ( .Y(n7651), .A(c_2_) );
  xor2 U2590 ( .Y(n4144), .A0(s_rad_i_33_), .A1(r1_2_33_) );
  inv01 U2591 ( .Y(n4145), .A(n4144) );
  xor2 U2592 ( .Y(n4146), .A0(s_rad_i_33_), .A1(n____return1382_33_) );
  inv01 U2593 ( .Y(n4147), .A(n4146) );
  xor2 U2594 ( .Y(n4148), .A0(s_rad_i_45_), .A1(n____return1382_45_) );
  inv01 U2595 ( .Y(n4149), .A(n4148) );
  xor2 U2596 ( .Y(n4150), .A0(s_rad_i_45_), .A1(r1_2_45_) );
  inv01 U2597 ( .Y(n4151), .A(n4150) );
  xor2 U2598 ( .Y(n4152), .A0(s_rad_i_21_), .A1(r1_2_21_) );
  inv01 U2599 ( .Y(n4153), .A(n4152) );
  xor2 U2600 ( .Y(n4154), .A0(s_rad_i_21_), .A1(n____return1382_21_) );
  inv01 U2601 ( .Y(n4155), .A(n4154) );
  xor2 U2602 ( .Y(n4156), .A0(s_rad_i_0_), .A1(r1_2_0_) );
  inv01 U2603 ( .Y(n4157), .A(n4156) );
  xor2 U2604 ( .Y(n4158), .A0(s_rad_i_0_), .A1(n____return1382_0_) );
  inv01 U2605 ( .Y(n4159), .A(n4158) );
  or02 U2606 ( .Y(n4160), .A0(n7674), .A1(n6945) );
  inv01 U2607 ( .Y(n4161), .A(n4160) );
  inv08 U2608 ( .Y(n7403), .A(n7402) );
  inv08 U2609 ( .Y(n7404), .A(n7402) );
  inv01 U2610 ( .Y(n3050), .A(n4162) );
  nor02 U2611 ( .Y(n4163), .A0(n7677), .A1(n7788) );
  nor02 U2612 ( .Y(n4164), .A0(n7362), .A1(n2810) );
  nor02 U2613 ( .Y(n4162), .A0(n4163), .A1(n4164) );
  nand02 U2614 ( .Y(n3077), .A0(n4165), .A1(n4166) );
  inv01 U2615 ( .Y(n4167), .A(n7677) );
  inv01 U2616 ( .Y(n4168), .A(n7676) );
  inv01 U2617 ( .Y(n4169), .A(n7675) );
  inv01 U2618 ( .Y(n4170), .A(n2809) );
  nand02 U2619 ( .Y(n4171), .A0(n4167), .A1(n4168) );
  nand02 U2620 ( .Y(n4172), .A0(n4167), .A1(n4169) );
  nand02 U2621 ( .Y(n4173), .A0(n4168), .A1(n4170) );
  nand02 U2622 ( .Y(n4174), .A0(n4169), .A1(n4170) );
  nand02 U2623 ( .Y(n4175), .A0(n4171), .A1(n4172) );
  inv01 U2624 ( .Y(n4165), .A(n4175) );
  nand02 U2625 ( .Y(n4176), .A0(n4173), .A1(n4174) );
  inv01 U2626 ( .Y(n4166), .A(n4176) );
  inv02 U2627 ( .Y(n7676), .A(n7348) );
  inv04 U2628 ( .Y(n4177), .A(n7618) );
  inv04 U2629 ( .Y(n7618), .A(c_3_) );
  inv01 U2630 ( .Y(n3076), .A(n4178) );
  nor02 U2631 ( .Y(n4179), .A0(n7385), .A1(n2811) );
  inv01 U2632 ( .Y(n4180), .A(n7770) );
  nor02 U2633 ( .Y(n4178), .A0(n4179), .A1(n4180) );
  inv01 U2634 ( .Y(n3054), .A(n4181) );
  nor02 U2635 ( .Y(n4182), .A0(n7385), .A1(n2825) );
  inv01 U2636 ( .Y(n4183), .A(n3285) );
  nor02 U2637 ( .Y(n4181), .A0(n4182), .A1(n4183) );
  inv01 U2638 ( .Y(n3071), .A(n4184) );
  nor02 U2639 ( .Y(n4185), .A0(n7385), .A1(n2832) );
  inv01 U2640 ( .Y(n4186), .A(n7775) );
  nor02 U2641 ( .Y(n4184), .A0(n4185), .A1(n4186) );
  inv01 U2642 ( .Y(n3052), .A(n4187) );
  nor02 U2643 ( .Y(n4188), .A0(n7385), .A1(n2827) );
  inv01 U2644 ( .Y(n4189), .A(n3327) );
  nor02 U2645 ( .Y(n4187), .A0(n4188), .A1(n4189) );
  inv01 U2646 ( .Y(n3061), .A(n4190) );
  nor02 U2647 ( .Y(n4191), .A0(n7385), .A1(n2817) );
  inv01 U2648 ( .Y(n4192), .A(n3161) );
  nor02 U2649 ( .Y(n4190), .A0(n4191), .A1(n4192) );
  inv01 U2650 ( .Y(n3074), .A(n4193) );
  nor02 U2651 ( .Y(n4194), .A0(n7385), .A1(n2829) );
  inv01 U2652 ( .Y(n4195), .A(n7772) );
  nor02 U2653 ( .Y(n4193), .A0(n4194), .A1(n4195) );
  inv01 U2654 ( .Y(n3060), .A(n4196) );
  nor02 U2655 ( .Y(n4197), .A0(n7385), .A1(n2818) );
  inv01 U2656 ( .Y(n4198), .A(n7780) );
  nor02 U2657 ( .Y(n4196), .A0(n4197), .A1(n4198) );
  inv01 U2658 ( .Y(n3066), .A(n4199) );
  nor02 U2659 ( .Y(n4200), .A0(n7385), .A1(n2812) );
  inv01 U2660 ( .Y(n4201), .A(n7777) );
  nor02 U2661 ( .Y(n4199), .A0(n4200), .A1(n4201) );
  inv01 U2662 ( .Y(n3072), .A(n4202) );
  nor02 U2663 ( .Y(n4203), .A0(n7385), .A1(n2831) );
  inv01 U2664 ( .Y(n4204), .A(n7774) );
  nor02 U2665 ( .Y(n4202), .A0(n4203), .A1(n4204) );
  inv01 U2666 ( .Y(n3067), .A(n4205) );
  nor02 U2667 ( .Y(n4206), .A0(n7385), .A1(n2836) );
  inv01 U2668 ( .Y(n4207), .A(n7776) );
  nor02 U2669 ( .Y(n4205), .A0(n4206), .A1(n4207) );
  inv01 U2670 ( .Y(n3065), .A(n4208) );
  nor02 U2671 ( .Y(n4209), .A0(n7385), .A1(n2813) );
  inv01 U2672 ( .Y(n4210), .A(n7778) );
  nor02 U2673 ( .Y(n4208), .A0(n4209), .A1(n4210) );
  inv01 U2674 ( .Y(n3053), .A(n4211) );
  nor02 U2675 ( .Y(n4212), .A0(n7385), .A1(n2826) );
  inv01 U2676 ( .Y(n4213), .A(n7786) );
  nor02 U2677 ( .Y(n4211), .A0(n4212), .A1(n4213) );
  inv01 U2678 ( .Y(n3056), .A(n4214) );
  nor02 U2679 ( .Y(n4215), .A0(n7385), .A1(n2823) );
  inv01 U2680 ( .Y(n4216), .A(n7784) );
  nor02 U2681 ( .Y(n4214), .A0(n4215), .A1(n4216) );
  inv01 U2682 ( .Y(n3055), .A(n4217) );
  nor02 U2683 ( .Y(n4218), .A0(n7385), .A1(n2824) );
  inv01 U2684 ( .Y(n4219), .A(n7785) );
  nor02 U2685 ( .Y(n4217), .A0(n4218), .A1(n4219) );
  inv01 U2686 ( .Y(n3062), .A(n4220) );
  nor02 U2687 ( .Y(n4221), .A0(n7385), .A1(n2816) );
  inv01 U2688 ( .Y(n4222), .A(n7779) );
  nor02 U2689 ( .Y(n4220), .A0(n4221), .A1(n4222) );
  inv01 U2690 ( .Y(n3057), .A(n4223) );
  nor02 U2691 ( .Y(n4224), .A0(n7385), .A1(n2821) );
  inv01 U2692 ( .Y(n4225), .A(n7783) );
  nor02 U2693 ( .Y(n4223), .A0(n4224), .A1(n4225) );
  inv01 U2694 ( .Y(n3075), .A(n4226) );
  nor02 U2695 ( .Y(n4227), .A0(n7385), .A1(n2822) );
  inv01 U2696 ( .Y(n4228), .A(n3127) );
  nor02 U2697 ( .Y(n4226), .A0(n4227), .A1(n4228) );
  inv01 U2698 ( .Y(n3059), .A(n4229) );
  nor02 U2699 ( .Y(n4230), .A0(n7385), .A1(n2819) );
  inv01 U2700 ( .Y(n4231), .A(n7781) );
  nor02 U2701 ( .Y(n4229), .A0(n4230), .A1(n4231) );
  inv01 U2702 ( .Y(n3070), .A(n4232) );
  nor02 U2703 ( .Y(n4233), .A0(n7385), .A1(n2833) );
  inv01 U2704 ( .Y(n4234), .A(n3247) );
  nor02 U2705 ( .Y(n4232), .A0(n4233), .A1(n4234) );
  inv01 U2706 ( .Y(n3058), .A(n4235) );
  nor02 U2707 ( .Y(n4236), .A0(n7385), .A1(n2820) );
  inv01 U2708 ( .Y(n4237), .A(n7782) );
  nor02 U2709 ( .Y(n4235), .A0(n4236), .A1(n4237) );
  inv01 U2710 ( .Y(n3068), .A(n4238) );
  nor02 U2711 ( .Y(n4239), .A0(n7385), .A1(n2835) );
  inv01 U2712 ( .Y(n4240), .A(n3373) );
  nor02 U2713 ( .Y(n4238), .A0(n4239), .A1(n4240) );
  inv01 U2714 ( .Y(n3069), .A(n4241) );
  nor02 U2715 ( .Y(n4242), .A0(n7385), .A1(n2834) );
  inv01 U2716 ( .Y(n4243), .A(n3207) );
  nor02 U2717 ( .Y(n4241), .A0(n4242), .A1(n4243) );
  inv01 U2718 ( .Y(n3051), .A(n4244) );
  nor02 U2719 ( .Y(n4245), .A0(n7385), .A1(n2828) );
  inv01 U2720 ( .Y(n4246), .A(n3287) );
  nor02 U2721 ( .Y(n4244), .A0(n4245), .A1(n4246) );
  inv01 U2722 ( .Y(n3063), .A(n4247) );
  nor02 U2723 ( .Y(n4248), .A0(n7385), .A1(n2815) );
  inv01 U2724 ( .Y(n4249), .A(n3325) );
  nor02 U2725 ( .Y(n4247), .A0(n4248), .A1(n4249) );
  inv01 U2726 ( .Y(n3073), .A(n4250) );
  nor02 U2727 ( .Y(n4251), .A0(n7385), .A1(n2830) );
  inv01 U2728 ( .Y(n4252), .A(n7773) );
  nor02 U2729 ( .Y(n4250), .A0(n4251), .A1(n4252) );
  inv01 U2730 ( .Y(n3064), .A(n4253) );
  nor02 U2731 ( .Y(n4254), .A0(n7385), .A1(n2814) );
  inv01 U2732 ( .Y(n4255), .A(n3209) );
  nor02 U2733 ( .Y(n4253), .A0(n4254), .A1(n4255) );
  or03 U2734 ( .Y(n4256), .A0(n____return1071), .A1(n7421), .A2(n6952) );
  inv01 U2735 ( .Y(n4257), .A(n4256) );
  inv01 U2736 ( .Y(n7529), .A(n4258) );
  nor02 U2737 ( .Y(n4259), .A0(n7439), .A1(n7482) );
  nor02 U2738 ( .Y(n4260), .A0(n7387), .A1(n6829) );
  nor02 U2739 ( .Y(n4261), .A0(n7437), .A1(n7483) );
  nor02 U2740 ( .Y(n4258), .A0(n4261), .A1(n4262) );
  nor02 U2741 ( .Y(n4263), .A0(n4259), .A1(n4260) );
  inv01 U2742 ( .Y(n4262), .A(n4263) );
  inv02 U2743 ( .Y(n7439), .A(n7370) );
  inv02 U2744 ( .Y(n4391), .A(n7925) );
  inv01 U2745 ( .Y(n2976), .A(n4264) );
  nor02 U2746 ( .Y(n4265), .A0(n7429), .A1(n7985) );
  nor02 U2747 ( .Y(n4266), .A0(n7423), .A1(n7984) );
  nor02 U2748 ( .Y(n4267), .A0(n7409), .A1(n7983) );
  nor02 U2749 ( .Y(n4264), .A0(n4267), .A1(n4268) );
  nor02 U2750 ( .Y(n4269), .A0(n4265), .A1(n4266) );
  inv01 U2751 ( .Y(n4268), .A(n4269) );
  nand02 U2752 ( .Y(n2977), .A0(n4270), .A1(n4271) );
  inv01 U2753 ( .Y(n4272), .A(n7982) );
  inv01 U2754 ( .Y(n4273), .A(n7427) );
  inv01 U2755 ( .Y(n4274), .A(n7981) );
  inv01 U2756 ( .Y(n4275), .A(n7425) );
  inv01 U2757 ( .Y(n4276), .A(n7980) );
  inv01 U2758 ( .Y(n4277), .A(n7407) );
  nand02 U2759 ( .Y(n4278), .A0(n4272), .A1(n4273) );
  nand02 U2760 ( .Y(n4279), .A0(n4274), .A1(n4275) );
  nand02 U2761 ( .Y(n4270), .A0(n4276), .A1(n4277) );
  nand02 U2762 ( .Y(n4280), .A0(n4278), .A1(n4279) );
  inv01 U2763 ( .Y(n4271), .A(n4280) );
  inv01 U2764 ( .Y(n2980), .A(n4281) );
  nor02 U2765 ( .Y(n4282), .A0(n7427), .A1(n7973) );
  nor02 U2766 ( .Y(n4283), .A0(n7425), .A1(n7972) );
  nor02 U2767 ( .Y(n4284), .A0(n7407), .A1(n7971) );
  nor02 U2768 ( .Y(n4281), .A0(n4284), .A1(n4285) );
  nor02 U2769 ( .Y(n4286), .A0(n4282), .A1(n4283) );
  inv01 U2770 ( .Y(n4285), .A(n4286) );
  inv01 U2771 ( .Y(n3024), .A(n4287) );
  nor02 U2772 ( .Y(n4288), .A0(n7429), .A1(n7855) );
  nor02 U2773 ( .Y(n4289), .A0(n7423), .A1(n7854) );
  nor02 U2774 ( .Y(n4290), .A0(n7409), .A1(n7853) );
  nor02 U2775 ( .Y(n4287), .A0(n4290), .A1(n4291) );
  nor02 U2776 ( .Y(n4292), .A0(n4288), .A1(n4289) );
  inv01 U2777 ( .Y(n4291), .A(n4292) );
  nand02 U2778 ( .Y(n2978), .A0(n4293), .A1(n4294) );
  inv01 U2779 ( .Y(n4295), .A(n7979) );
  inv01 U2780 ( .Y(n4296), .A(n7428) );
  inv01 U2781 ( .Y(n4297), .A(n7978) );
  inv01 U2782 ( .Y(n4298), .A(n7424) );
  inv01 U2783 ( .Y(n4299), .A(n7977) );
  inv01 U2784 ( .Y(n4300), .A(n7408) );
  nand02 U2785 ( .Y(n4301), .A0(n4295), .A1(n4296) );
  nand02 U2786 ( .Y(n4302), .A0(n4297), .A1(n4298) );
  nand02 U2787 ( .Y(n4293), .A0(n4299), .A1(n4300) );
  nand02 U2788 ( .Y(n4303), .A0(n4301), .A1(n4302) );
  inv01 U2789 ( .Y(n4294), .A(n4303) );
  inv01 U2790 ( .Y(n2993), .A(n4304) );
  nor02 U2791 ( .Y(n4305), .A0(n7428), .A1(n7934) );
  nor02 U2792 ( .Y(n4306), .A0(n7424), .A1(n7933) );
  nor02 U2793 ( .Y(n4307), .A0(n7408), .A1(n7932) );
  nor02 U2794 ( .Y(n4304), .A0(n4307), .A1(n4308) );
  nor02 U2795 ( .Y(n4309), .A0(n4305), .A1(n4306) );
  inv01 U2796 ( .Y(n4308), .A(n4309) );
  nand02 U2797 ( .Y(n3046), .A0(n4310), .A1(n4311) );
  inv01 U2798 ( .Y(n4312), .A(n7798) );
  inv01 U2799 ( .Y(n4313), .A(n7427) );
  inv01 U2800 ( .Y(n4314), .A(n7797) );
  inv01 U2801 ( .Y(n4315), .A(n7425) );
  inv01 U2802 ( .Y(n4316), .A(n7796) );
  inv01 U2803 ( .Y(n4317), .A(n7407) );
  nand02 U2804 ( .Y(n4318), .A0(n4312), .A1(n4313) );
  nand02 U2805 ( .Y(n4319), .A0(n4314), .A1(n4315) );
  nand02 U2806 ( .Y(n4310), .A0(n4316), .A1(n4317) );
  nand02 U2807 ( .Y(n4320), .A0(n4318), .A1(n4319) );
  inv01 U2808 ( .Y(n4311), .A(n4320) );
  inv01 U2809 ( .Y(n3010), .A(n4321) );
  nor02 U2810 ( .Y(n4322), .A0(n7429), .A1(n7726) );
  nor02 U2811 ( .Y(n4323), .A0(n7425), .A1(n7889) );
  nor02 U2812 ( .Y(n4324), .A0(n7407), .A1(n7888) );
  nor02 U2813 ( .Y(n4321), .A0(n4324), .A1(n4325) );
  nor02 U2814 ( .Y(n4326), .A0(n4322), .A1(n4323) );
  inv01 U2815 ( .Y(n4325), .A(n4326) );
  inv01 U2816 ( .Y(n2983), .A(n4327) );
  nor02 U2817 ( .Y(n4328), .A0(n7427), .A1(n7964) );
  nor02 U2818 ( .Y(n4329), .A0(n7425), .A1(n7963) );
  nor02 U2819 ( .Y(n4330), .A0(n7407), .A1(n7962) );
  nor02 U2820 ( .Y(n4327), .A0(n4330), .A1(n4331) );
  nor02 U2821 ( .Y(n4332), .A0(n4328), .A1(n4329) );
  inv01 U2822 ( .Y(n4331), .A(n4332) );
  nand02 U2823 ( .Y(n3030), .A0(n4333), .A1(n4334) );
  inv01 U2824 ( .Y(n4335), .A(n7839) );
  inv01 U2825 ( .Y(n4336), .A(n7429) );
  inv01 U2826 ( .Y(n4337), .A(n7838) );
  inv01 U2827 ( .Y(n4338), .A(n7423) );
  inv01 U2828 ( .Y(n4339), .A(n7837) );
  inv01 U2829 ( .Y(n4340), .A(n7409) );
  nand02 U2830 ( .Y(n4341), .A0(n4335), .A1(n4336) );
  nand02 U2831 ( .Y(n4342), .A0(n4337), .A1(n4338) );
  nand02 U2832 ( .Y(n4333), .A0(n4339), .A1(n4340) );
  nand02 U2833 ( .Y(n4343), .A0(n4341), .A1(n4342) );
  inv01 U2834 ( .Y(n4334), .A(n4343) );
  nand02 U2835 ( .Y(n2972), .A0(n4344), .A1(n4345) );
  inv01 U2836 ( .Y(n4346), .A(n7997) );
  inv01 U2837 ( .Y(n4347), .A(n7429) );
  inv01 U2838 ( .Y(n4348), .A(n7996) );
  inv01 U2839 ( .Y(n4349), .A(n7424) );
  inv01 U2840 ( .Y(n4350), .A(n7995) );
  inv01 U2841 ( .Y(n4351), .A(n7408) );
  nand02 U2842 ( .Y(n4352), .A0(n4346), .A1(n4347) );
  nand02 U2843 ( .Y(n4353), .A0(n4348), .A1(n4349) );
  nand02 U2844 ( .Y(n4344), .A0(n4350), .A1(n4351) );
  nand02 U2845 ( .Y(n4354), .A0(n4352), .A1(n4353) );
  inv01 U2846 ( .Y(n4345), .A(n4354) );
  inv01 U2847 ( .Y(n3035), .A(n4355) );
  nor02 U2848 ( .Y(n4356), .A0(n7429), .A1(n7751) );
  nor02 U2849 ( .Y(n4357), .A0(n7424), .A1(n7826) );
  nor02 U2850 ( .Y(n4358), .A0(n7408), .A1(n7825) );
  nor02 U2851 ( .Y(n4355), .A0(n4358), .A1(n4359) );
  nor02 U2852 ( .Y(n4360), .A0(n4356), .A1(n4357) );
  inv01 U2853 ( .Y(n4359), .A(n4360) );
  nand02 U2854 ( .Y(n2988), .A0(n4361), .A1(n4362) );
  inv01 U2855 ( .Y(n4363), .A(n7949) );
  inv01 U2856 ( .Y(n4364), .A(n7429) );
  inv01 U2857 ( .Y(n4365), .A(n7948) );
  inv01 U2858 ( .Y(n4366), .A(n7423) );
  inv01 U2859 ( .Y(n4367), .A(n7947) );
  inv01 U2860 ( .Y(n4368), .A(n7409) );
  nand02 U2861 ( .Y(n4369), .A0(n4363), .A1(n4364) );
  nand02 U2862 ( .Y(n4370), .A0(n4365), .A1(n4366) );
  nand02 U2863 ( .Y(n4361), .A0(n4367), .A1(n4368) );
  nand02 U2864 ( .Y(n4371), .A0(n4369), .A1(n4370) );
  inv01 U2865 ( .Y(n4362), .A(n4371) );
  nand02 U2866 ( .Y(n3015), .A0(n4372), .A1(n4373) );
  inv01 U2867 ( .Y(n4374), .A(n7876) );
  inv01 U2868 ( .Y(n4375), .A(n7429) );
  inv01 U2869 ( .Y(n4376), .A(n7875) );
  inv01 U2870 ( .Y(n4377), .A(n7423) );
  inv01 U2871 ( .Y(n4378), .A(n7874) );
  inv01 U2872 ( .Y(n4379), .A(n7409) );
  nand02 U2873 ( .Y(n4380), .A0(n4374), .A1(n4375) );
  nand02 U2874 ( .Y(n4381), .A0(n4376), .A1(n4377) );
  nand02 U2875 ( .Y(n4372), .A0(n4378), .A1(n4379) );
  nand02 U2876 ( .Y(n4382), .A0(n4380), .A1(n4381) );
  inv01 U2877 ( .Y(n4373), .A(n4382) );
  inv01 U2878 ( .Y(n3048), .A(n4383) );
  nor02 U2879 ( .Y(n4384), .A0(n7428), .A1(n7793) );
  nor02 U2880 ( .Y(n4385), .A0(n7423), .A1(n7792) );
  nor02 U2881 ( .Y(n4386), .A0(n7409), .A1(n7790) );
  nor02 U2882 ( .Y(n4383), .A0(n4386), .A1(n4387) );
  nor02 U2883 ( .Y(n4388), .A0(n4384), .A1(n4385) );
  inv01 U2884 ( .Y(n4387), .A(n4388) );
  nand02 U2885 ( .Y(n2996), .A0(n4389), .A1(n4390) );
  inv01 U2886 ( .Y(n4392), .A(n7428) );
  inv01 U2887 ( .Y(n4393), .A(n7924) );
  inv01 U2888 ( .Y(n4394), .A(n7424) );
  inv01 U2889 ( .Y(n4395), .A(n7923) );
  inv01 U2890 ( .Y(n4396), .A(n7408) );
  nand02 U2891 ( .Y(n4397), .A0(n4391), .A1(n4392) );
  nand02 U2892 ( .Y(n4398), .A0(n4393), .A1(n4394) );
  nand02 U2893 ( .Y(n4389), .A0(n4395), .A1(n4396) );
  nand02 U2894 ( .Y(n4399), .A0(n4397), .A1(n4398) );
  inv01 U2895 ( .Y(n4390), .A(n4399) );
  nand02 U2896 ( .Y(n3038), .A0(n4400), .A1(n4401) );
  inv01 U2897 ( .Y(n4402), .A(n7818) );
  inv01 U2898 ( .Y(n4403), .A(n7428) );
  inv01 U2899 ( .Y(n4404), .A(n7817) );
  inv01 U2900 ( .Y(n4405), .A(n7424) );
  inv01 U2901 ( .Y(n4406), .A(n7816) );
  inv01 U2902 ( .Y(n4407), .A(n7408) );
  nand02 U2903 ( .Y(n4408), .A0(n4402), .A1(n4403) );
  nand02 U2904 ( .Y(n4409), .A0(n4404), .A1(n4405) );
  nand02 U2905 ( .Y(n4400), .A0(n4406), .A1(n4407) );
  nand02 U2906 ( .Y(n4410), .A0(n4408), .A1(n4409) );
  inv01 U2907 ( .Y(n4401), .A(n4410) );
  inv01 U2908 ( .Y(n3020), .A(n4411) );
  nor02 U2909 ( .Y(n4412), .A0(n7427), .A1(n7864) );
  nor02 U2910 ( .Y(n4413), .A0(n7424), .A1(n7863) );
  nor02 U2911 ( .Y(n4414), .A0(n7408), .A1(n7862) );
  nor02 U2912 ( .Y(n4411), .A0(n4414), .A1(n4415) );
  nor02 U2913 ( .Y(n4416), .A0(n4412), .A1(n4413) );
  inv01 U2914 ( .Y(n4415), .A(n4416) );
  nand02 U2915 ( .Y(n3037), .A0(n4417), .A1(n4418) );
  inv01 U2916 ( .Y(n4419), .A(n7821) );
  inv01 U2917 ( .Y(n4420), .A(n7428) );
  inv01 U2918 ( .Y(n4421), .A(n7820) );
  inv01 U2919 ( .Y(n4422), .A(n7425) );
  inv01 U2920 ( .Y(n4423), .A(n7819) );
  inv01 U2921 ( .Y(n4424), .A(n7407) );
  nand02 U2922 ( .Y(n4425), .A0(n4419), .A1(n4420) );
  nand02 U2923 ( .Y(n4426), .A0(n4421), .A1(n4422) );
  nand02 U2924 ( .Y(n4417), .A0(n4423), .A1(n4424) );
  nand02 U2925 ( .Y(n4427), .A0(n4425), .A1(n4426) );
  inv01 U2926 ( .Y(n4418), .A(n4427) );
  nand02 U2927 ( .Y(n2974), .A0(n4428), .A1(n4429) );
  inv01 U2928 ( .Y(n4430), .A(n7991) );
  inv01 U2929 ( .Y(n4431), .A(n7427) );
  inv01 U2930 ( .Y(n4432), .A(n7990) );
  inv01 U2931 ( .Y(n4433), .A(n7425) );
  inv01 U2932 ( .Y(n4434), .A(n7989) );
  inv01 U2933 ( .Y(n4435), .A(n7407) );
  nand02 U2934 ( .Y(n4436), .A0(n4430), .A1(n4431) );
  nand02 U2935 ( .Y(n4437), .A0(n4432), .A1(n4433) );
  nand02 U2936 ( .Y(n4428), .A0(n4434), .A1(n4435) );
  nand02 U2937 ( .Y(n4438), .A0(n4436), .A1(n4437) );
  inv01 U2938 ( .Y(n4429), .A(n4438) );
  inv01 U2939 ( .Y(n3007), .A(n4439) );
  nor02 U2940 ( .Y(n4440), .A0(n7427), .A1(n7897) );
  nor02 U2941 ( .Y(n4441), .A0(n7425), .A1(n7896) );
  nor02 U2942 ( .Y(n4442), .A0(n7407), .A1(n7895) );
  nor02 U2943 ( .Y(n4439), .A0(n4442), .A1(n4443) );
  nor02 U2944 ( .Y(n4444), .A0(n4440), .A1(n4441) );
  inv01 U2945 ( .Y(n4443), .A(n4444) );
  nand02 U2946 ( .Y(n2987), .A0(n4445), .A1(n4446) );
  inv01 U2947 ( .Y(n4447), .A(n7952) );
  inv01 U2948 ( .Y(n4448), .A(n7428) );
  inv01 U2949 ( .Y(n4449), .A(n7951) );
  inv01 U2950 ( .Y(n4450), .A(n7424) );
  inv01 U2951 ( .Y(n4451), .A(n7950) );
  inv01 U2952 ( .Y(n4452), .A(n7408) );
  nand02 U2953 ( .Y(n4453), .A0(n4447), .A1(n4448) );
  nand02 U2954 ( .Y(n4454), .A0(n4449), .A1(n4450) );
  nand02 U2955 ( .Y(n4445), .A0(n4451), .A1(n4452) );
  nand02 U2956 ( .Y(n4455), .A0(n4453), .A1(n4454) );
  inv01 U2957 ( .Y(n4446), .A(n4455) );
  inv01 U2958 ( .Y(n2984), .A(n4456) );
  nor02 U2959 ( .Y(n4457), .A0(n7428), .A1(n7961) );
  nor02 U2960 ( .Y(n4458), .A0(n7424), .A1(n7960) );
  nor02 U2961 ( .Y(n4459), .A0(n7408), .A1(n7959) );
  nor02 U2962 ( .Y(n4456), .A0(n4459), .A1(n4460) );
  nor02 U2963 ( .Y(n4461), .A0(n4457), .A1(n4458) );
  inv01 U2964 ( .Y(n4460), .A(n4461) );
  nand02 U2965 ( .Y(n3012), .A0(n4462), .A1(n4463) );
  inv01 U2966 ( .Y(n4464), .A(n7885) );
  inv01 U2967 ( .Y(n4465), .A(n7429) );
  inv01 U2968 ( .Y(n4466), .A(n7884) );
  inv01 U2969 ( .Y(n4467), .A(n7423) );
  inv01 U2970 ( .Y(n4468), .A(n7883) );
  inv01 U2971 ( .Y(n4469), .A(n7409) );
  nand02 U2972 ( .Y(n4470), .A0(n4464), .A1(n4465) );
  nand02 U2973 ( .Y(n4471), .A0(n4466), .A1(n4467) );
  nand02 U2974 ( .Y(n4462), .A0(n4468), .A1(n4469) );
  nand02 U2975 ( .Y(n4472), .A0(n4470), .A1(n4471) );
  inv01 U2976 ( .Y(n4463), .A(n4472) );
  nand02 U2977 ( .Y(n3006), .A0(n4473), .A1(n4474) );
  inv01 U2978 ( .Y(n4475), .A(n7730) );
  inv01 U2979 ( .Y(n4476), .A(n7429) );
  inv01 U2980 ( .Y(n4477), .A(n7899) );
  inv01 U2981 ( .Y(n4478), .A(n7423) );
  inv01 U2982 ( .Y(n4479), .A(n7898) );
  inv01 U2983 ( .Y(n4480), .A(n7409) );
  nand02 U2984 ( .Y(n4481), .A0(n4475), .A1(n4476) );
  nand02 U2985 ( .Y(n4482), .A0(n4477), .A1(n4478) );
  nand02 U2986 ( .Y(n4473), .A0(n4479), .A1(n4480) );
  nand02 U2987 ( .Y(n4483), .A0(n4481), .A1(n4482) );
  inv01 U2988 ( .Y(n4474), .A(n4483) );
  inv01 U2989 ( .Y(n2991), .A(n4484) );
  nor02 U2990 ( .Y(n4485), .A0(n7429), .A1(n7940) );
  nor02 U2991 ( .Y(n4486), .A0(n7423), .A1(n7939) );
  nor02 U2992 ( .Y(n4487), .A0(n7409), .A1(n7938) );
  nor02 U2993 ( .Y(n4484), .A0(n4487), .A1(n4488) );
  nor02 U2994 ( .Y(n4489), .A0(n4485), .A1(n4486) );
  inv01 U2995 ( .Y(n4488), .A(n4489) );
  nand02 U2996 ( .Y(n2989), .A0(n4490), .A1(n4491) );
  inv01 U2997 ( .Y(n4492), .A(n7946) );
  inv01 U2998 ( .Y(n4493), .A(n7427) );
  inv01 U2999 ( .Y(n4494), .A(n7945) );
  inv01 U3000 ( .Y(n4495), .A(n7425) );
  inv01 U3001 ( .Y(n4496), .A(n7944) );
  inv01 U3002 ( .Y(n4497), .A(n7407) );
  nand02 U3003 ( .Y(n4498), .A0(n4492), .A1(n4493) );
  nand02 U3004 ( .Y(n4499), .A0(n4494), .A1(n4495) );
  nand02 U3005 ( .Y(n4490), .A0(n4496), .A1(n4497) );
  nand02 U3006 ( .Y(n4500), .A0(n4498), .A1(n4499) );
  inv01 U3007 ( .Y(n4491), .A(n4500) );
  inv01 U3008 ( .Y(n3043), .A(n4501) );
  nor02 U3009 ( .Y(n4502), .A0(n7429), .A1(n7806) );
  nor02 U3010 ( .Y(n4503), .A0(n7425), .A1(n7805) );
  nor02 U3011 ( .Y(n4504), .A0(n7407), .A1(n7804) );
  nor02 U3012 ( .Y(n4501), .A0(n4504), .A1(n4505) );
  nor02 U3013 ( .Y(n4506), .A0(n4502), .A1(n4503) );
  inv01 U3014 ( .Y(n4505), .A(n4506) );
  inv01 U3015 ( .Y(n3025), .A(n4507) );
  nor02 U3016 ( .Y(n4508), .A0(n7428), .A1(n7852) );
  nor02 U3017 ( .Y(n4509), .A0(n7425), .A1(n7851) );
  nor02 U3018 ( .Y(n4510), .A0(n7407), .A1(n7850) );
  nor02 U3019 ( .Y(n4507), .A0(n4510), .A1(n4511) );
  nor02 U3020 ( .Y(n4512), .A0(n4508), .A1(n4509) );
  inv01 U3021 ( .Y(n4511), .A(n4512) );
  nand02 U3022 ( .Y(n3026), .A0(n4513), .A1(n4514) );
  inv01 U3023 ( .Y(n4515), .A(n7849) );
  inv01 U3024 ( .Y(n4516), .A(n7428) );
  inv01 U3025 ( .Y(n4517), .A(n7848) );
  inv01 U3026 ( .Y(n4518), .A(n7424) );
  inv01 U3027 ( .Y(n4519), .A(n7847) );
  inv01 U3028 ( .Y(n4520), .A(n7408) );
  nand02 U3029 ( .Y(n4521), .A0(n4515), .A1(n4516) );
  nand02 U3030 ( .Y(n4522), .A0(n4517), .A1(n4518) );
  nand02 U3031 ( .Y(n4513), .A0(n4519), .A1(n4520) );
  nand02 U3032 ( .Y(n4523), .A0(n4521), .A1(n4522) );
  inv01 U3033 ( .Y(n4514), .A(n4523) );
  inv01 U3034 ( .Y(n3017), .A(n4524) );
  nor02 U3035 ( .Y(n4525), .A0(n7427), .A1(n7768) );
  nor02 U3036 ( .Y(n4526), .A0(n7424), .A1(n7871) );
  nor02 U3037 ( .Y(n4527), .A0(n7408), .A1(n7870) );
  nor02 U3038 ( .Y(n4524), .A0(n4527), .A1(n4528) );
  nor02 U3039 ( .Y(n4529), .A0(n4525), .A1(n4526) );
  inv01 U3040 ( .Y(n4528), .A(n4529) );
  nand02 U3041 ( .Y(n3036), .A0(n4530), .A1(n4531) );
  inv01 U3042 ( .Y(n4532), .A(n7824) );
  inv01 U3043 ( .Y(n4533), .A(n7427) );
  inv01 U3044 ( .Y(n4534), .A(n7823) );
  inv01 U3045 ( .Y(n4535), .A(n7423) );
  inv01 U3046 ( .Y(n4536), .A(n7822) );
  inv01 U3047 ( .Y(n4537), .A(n7409) );
  nand02 U3048 ( .Y(n4538), .A0(n4532), .A1(n4533) );
  nand02 U3049 ( .Y(n4539), .A0(n4534), .A1(n4535) );
  nand02 U3050 ( .Y(n4530), .A0(n4536), .A1(n4537) );
  nand02 U3051 ( .Y(n4540), .A0(n4538), .A1(n4539) );
  inv01 U3052 ( .Y(n4531), .A(n4540) );
  nand02 U3053 ( .Y(n3018), .A0(n4541), .A1(n4542) );
  inv01 U3054 ( .Y(n4543), .A(n7766) );
  inv01 U3055 ( .Y(n4544), .A(n7428) );
  inv01 U3056 ( .Y(n4545), .A(n7869) );
  inv01 U3057 ( .Y(n4546), .A(n7423) );
  inv01 U3058 ( .Y(n4547), .A(n7868) );
  inv01 U3059 ( .Y(n4548), .A(n7409) );
  nand02 U3060 ( .Y(n4549), .A0(n4543), .A1(n4544) );
  nand02 U3061 ( .Y(n4550), .A0(n4545), .A1(n4546) );
  nand02 U3062 ( .Y(n4541), .A0(n4547), .A1(n4548) );
  nand02 U3063 ( .Y(n4551), .A0(n4549), .A1(n4550) );
  inv01 U3064 ( .Y(n4542), .A(n4551) );
  inv01 U3065 ( .Y(n3045), .A(n4552) );
  nor02 U3066 ( .Y(n4553), .A0(n7428), .A1(n7801) );
  nor02 U3067 ( .Y(n4554), .A0(n7423), .A1(n7800) );
  nor02 U3068 ( .Y(n4555), .A0(n7409), .A1(n7799) );
  nor02 U3069 ( .Y(n4552), .A0(n4555), .A1(n4556) );
  nor02 U3070 ( .Y(n4557), .A0(n4553), .A1(n4554) );
  inv01 U3071 ( .Y(n4556), .A(n4557) );
  nand02 U3072 ( .Y(n3002), .A0(n4558), .A1(n4559) );
  inv01 U3073 ( .Y(n4560), .A(n7909) );
  inv01 U3074 ( .Y(n4561), .A(n7427) );
  inv01 U3075 ( .Y(n4562), .A(n7908) );
  inv01 U3076 ( .Y(n4563), .A(n7424) );
  inv01 U3077 ( .Y(n4564), .A(n7907) );
  inv01 U3078 ( .Y(n4565), .A(n7408) );
  nand02 U3079 ( .Y(n4566), .A0(n4560), .A1(n4561) );
  nand02 U3080 ( .Y(n4567), .A0(n4562), .A1(n4563) );
  nand02 U3081 ( .Y(n4558), .A0(n4564), .A1(n4565) );
  nand02 U3082 ( .Y(n4568), .A0(n4566), .A1(n4567) );
  inv01 U3083 ( .Y(n4559), .A(n4568) );
  inv01 U3084 ( .Y(n3011), .A(n4569) );
  nor02 U3085 ( .Y(n4570), .A0(n7427), .A1(n7724) );
  nor02 U3086 ( .Y(n4571), .A0(n7424), .A1(n7887) );
  nor02 U3087 ( .Y(n4572), .A0(n7408), .A1(n7886) );
  nor02 U3088 ( .Y(n4569), .A0(n4572), .A1(n4573) );
  nor02 U3089 ( .Y(n4574), .A0(n4570), .A1(n4571) );
  inv01 U3090 ( .Y(n4573), .A(n4574) );
  nand02 U3091 ( .Y(n3004), .A0(n4575), .A1(n4576) );
  inv01 U3092 ( .Y(n4577), .A(n7731) );
  inv01 U3093 ( .Y(n4578), .A(n7427) );
  inv01 U3094 ( .Y(n4579), .A(n7903) );
  inv01 U3095 ( .Y(n4580), .A(n7425) );
  inv01 U3096 ( .Y(n4581), .A(n7902) );
  inv01 U3097 ( .Y(n4582), .A(n7407) );
  nand02 U3098 ( .Y(n4583), .A0(n4577), .A1(n4578) );
  nand02 U3099 ( .Y(n4584), .A0(n4579), .A1(n4580) );
  nand02 U3100 ( .Y(n4575), .A0(n4581), .A1(n4582) );
  nand02 U3101 ( .Y(n4585), .A0(n4583), .A1(n4584) );
  inv01 U3102 ( .Y(n4576), .A(n4585) );
  nand02 U3103 ( .Y(n3016), .A0(n4586), .A1(n4587) );
  inv01 U3104 ( .Y(n4588), .A(n7767) );
  inv01 U3105 ( .Y(n4589), .A(n7428) );
  inv01 U3106 ( .Y(n4590), .A(n7873) );
  inv01 U3107 ( .Y(n4591), .A(n7425) );
  inv01 U3108 ( .Y(n4592), .A(n7872) );
  inv01 U3109 ( .Y(n4593), .A(n7407) );
  nand02 U3110 ( .Y(n4594), .A0(n4588), .A1(n4589) );
  nand02 U3111 ( .Y(n4595), .A0(n4590), .A1(n4591) );
  nand02 U3112 ( .Y(n4586), .A0(n4592), .A1(n4593) );
  nand02 U3113 ( .Y(n4596), .A0(n4594), .A1(n4595) );
  inv01 U3114 ( .Y(n4587), .A(n4596) );
  inv01 U3115 ( .Y(n3001), .A(n4597) );
  nor02 U3116 ( .Y(n4598), .A0(n7429), .A1(n7912) );
  nor02 U3117 ( .Y(n4599), .A0(n7425), .A1(n7911) );
  nor02 U3118 ( .Y(n4600), .A0(n7407), .A1(n7910) );
  nor02 U3119 ( .Y(n4597), .A0(n4600), .A1(n4601) );
  nor02 U3120 ( .Y(n4602), .A0(n4598), .A1(n4599) );
  inv01 U3121 ( .Y(n4601), .A(n4602) );
  nand02 U3122 ( .Y(n3000), .A0(n4603), .A1(n4604) );
  inv01 U3123 ( .Y(n4605), .A(n7915) );
  inv01 U3124 ( .Y(n4606), .A(n7428) );
  inv01 U3125 ( .Y(n4607), .A(n7914) );
  inv01 U3126 ( .Y(n4608), .A(n7423) );
  inv01 U3127 ( .Y(n4609), .A(n7913) );
  inv01 U3128 ( .Y(n4610), .A(n7409) );
  nand02 U3129 ( .Y(n4611), .A0(n4605), .A1(n4606) );
  nand02 U3130 ( .Y(n4612), .A0(n4607), .A1(n4608) );
  nand02 U3131 ( .Y(n4603), .A0(n4609), .A1(n4610) );
  nand02 U3132 ( .Y(n4613), .A0(n4611), .A1(n4612) );
  inv01 U3133 ( .Y(n4604), .A(n4613) );
  nand02 U3134 ( .Y(n2982), .A0(n4614), .A1(n4615) );
  inv01 U3135 ( .Y(n4616), .A(n7967) );
  inv01 U3136 ( .Y(n4617), .A(n7429) );
  inv01 U3137 ( .Y(n4618), .A(n7966) );
  inv01 U3138 ( .Y(n4619), .A(n7423) );
  inv01 U3139 ( .Y(n4620), .A(n7965) );
  inv01 U3140 ( .Y(n4621), .A(n7409) );
  nand02 U3141 ( .Y(n4622), .A0(n4616), .A1(n4617) );
  nand02 U3142 ( .Y(n4623), .A0(n4618), .A1(n4619) );
  nand02 U3143 ( .Y(n4614), .A0(n4620), .A1(n4621) );
  nand02 U3144 ( .Y(n4624), .A0(n4622), .A1(n4623) );
  inv01 U3145 ( .Y(n4615), .A(n4624) );
  inv01 U3146 ( .Y(n3033), .A(n4625) );
  nor02 U3147 ( .Y(n4626), .A0(n7427), .A1(n7752) );
  nor02 U3148 ( .Y(n4627), .A0(n7423), .A1(n7830) );
  nor02 U3149 ( .Y(n4628), .A0(n7409), .A1(n7829) );
  nor02 U3150 ( .Y(n4625), .A0(n4628), .A1(n4629) );
  nor02 U3151 ( .Y(n4630), .A0(n4626), .A1(n4627) );
  inv01 U3152 ( .Y(n4629), .A(n4630) );
  nand02 U3153 ( .Y(n3044), .A0(n4631), .A1(n4632) );
  inv01 U3154 ( .Y(n4633), .A(n7738) );
  inv01 U3155 ( .Y(n4634), .A(n7429) );
  inv01 U3156 ( .Y(n4635), .A(n7803) );
  inv01 U3157 ( .Y(n4636), .A(n7424) );
  inv01 U3158 ( .Y(n4637), .A(n7802) );
  inv01 U3159 ( .Y(n4638), .A(n7408) );
  nand02 U3160 ( .Y(n4639), .A0(n4633), .A1(n4634) );
  nand02 U3161 ( .Y(n4640), .A0(n4635), .A1(n4636) );
  nand02 U3162 ( .Y(n4631), .A0(n4637), .A1(n4638) );
  nand02 U3163 ( .Y(n4641), .A0(n4639), .A1(n4640) );
  inv01 U3164 ( .Y(n4632), .A(n4641) );
  nand02 U3165 ( .Y(n3029), .A0(n4642), .A1(n4643) );
  inv01 U3166 ( .Y(n4644), .A(n7756) );
  inv01 U3167 ( .Y(n4645), .A(n7428) );
  inv01 U3168 ( .Y(n4646), .A(n7841) );
  inv01 U3169 ( .Y(n4647), .A(n7424) );
  inv01 U3170 ( .Y(n4648), .A(n7840) );
  inv01 U3171 ( .Y(n4649), .A(n7408) );
  nand02 U3172 ( .Y(n4650), .A0(n4644), .A1(n4645) );
  nand02 U3173 ( .Y(n4651), .A0(n4646), .A1(n4647) );
  nand02 U3174 ( .Y(n4642), .A0(n4648), .A1(n4649) );
  nand02 U3175 ( .Y(n4652), .A0(n4650), .A1(n4651) );
  inv01 U3176 ( .Y(n4643), .A(n4652) );
  inv01 U3177 ( .Y(n3032), .A(n4653) );
  nor02 U3178 ( .Y(n4654), .A0(n7427), .A1(n7833) );
  nor02 U3179 ( .Y(n4655), .A0(n7424), .A1(n7832) );
  nor02 U3180 ( .Y(n4656), .A0(n7408), .A1(n7831) );
  nor02 U3181 ( .Y(n4653), .A0(n4656), .A1(n4657) );
  nor02 U3182 ( .Y(n4658), .A0(n4654), .A1(n4655) );
  inv01 U3183 ( .Y(n4657), .A(n4658) );
  nand02 U3184 ( .Y(n2995), .A0(n4659), .A1(n4660) );
  inv01 U3185 ( .Y(n4661), .A(n7928) );
  inv01 U3186 ( .Y(n4662), .A(n7427) );
  inv01 U3187 ( .Y(n4663), .A(n7927) );
  inv01 U3188 ( .Y(n4664), .A(n7425) );
  inv01 U3189 ( .Y(n4665), .A(n7926) );
  inv01 U3190 ( .Y(n4666), .A(n7407) );
  nand02 U3191 ( .Y(n4667), .A0(n4661), .A1(n4662) );
  nand02 U3192 ( .Y(n4668), .A0(n4663), .A1(n4664) );
  nand02 U3193 ( .Y(n4659), .A0(n4665), .A1(n4666) );
  nand02 U3194 ( .Y(n4669), .A0(n4667), .A1(n4668) );
  inv01 U3195 ( .Y(n4660), .A(n4669) );
  nand02 U3196 ( .Y(n2971), .A0(n4670), .A1(n4671) );
  inv01 U3197 ( .Y(n4672), .A(n8000) );
  inv01 U3198 ( .Y(n4673), .A(n7428) );
  inv01 U3199 ( .Y(n4674), .A(n7999) );
  inv01 U3200 ( .Y(n4675), .A(n7425) );
  inv01 U3201 ( .Y(n4676), .A(n7998) );
  inv01 U3202 ( .Y(n4677), .A(n7407) );
  nand02 U3203 ( .Y(n4678), .A0(n4672), .A1(n4673) );
  nand02 U3204 ( .Y(n4679), .A0(n4674), .A1(n4675) );
  nand02 U3205 ( .Y(n4670), .A0(n4676), .A1(n4677) );
  nand02 U3206 ( .Y(n4680), .A0(n4678), .A1(n4679) );
  inv01 U3207 ( .Y(n4671), .A(n4680) );
  inv01 U3208 ( .Y(n3034), .A(n4681) );
  nor02 U3209 ( .Y(n4682), .A0(n7427), .A1(n7753) );
  nor02 U3210 ( .Y(n4683), .A0(n7425), .A1(n7828) );
  nor02 U3211 ( .Y(n4684), .A0(n7407), .A1(n7827) );
  nor02 U3212 ( .Y(n4681), .A0(n4684), .A1(n4685) );
  nor02 U3213 ( .Y(n4686), .A0(n4682), .A1(n4683) );
  inv01 U3214 ( .Y(n4685), .A(n4686) );
  nand02 U3215 ( .Y(n2990), .A0(n4687), .A1(n4688) );
  inv01 U3216 ( .Y(n4689), .A(n7943) );
  inv01 U3217 ( .Y(n4690), .A(n7428) );
  inv01 U3218 ( .Y(n4691), .A(n7942) );
  inv01 U3219 ( .Y(n4692), .A(n7424) );
  inv01 U3220 ( .Y(n4693), .A(n7941) );
  inv01 U3221 ( .Y(n4694), .A(n7408) );
  nand02 U3222 ( .Y(n4695), .A0(n4689), .A1(n4690) );
  nand02 U3223 ( .Y(n4696), .A0(n4691), .A1(n4692) );
  nand02 U3224 ( .Y(n4687), .A0(n4693), .A1(n4694) );
  nand02 U3225 ( .Y(n4697), .A0(n4695), .A1(n4696) );
  inv01 U3226 ( .Y(n4688), .A(n4697) );
  inv01 U3227 ( .Y(n2999), .A(n4698) );
  nor02 U3228 ( .Y(n4699), .A0(n7427), .A1(n7736) );
  nor02 U3229 ( .Y(n4700), .A0(n7424), .A1(n7917) );
  nor02 U3230 ( .Y(n4701), .A0(n7408), .A1(n7916) );
  nor02 U3231 ( .Y(n4698), .A0(n4701), .A1(n4702) );
  nor02 U3232 ( .Y(n4703), .A0(n4699), .A1(n4700) );
  inv01 U3233 ( .Y(n4702), .A(n4703) );
  nand02 U3234 ( .Y(n3042), .A0(n4704), .A1(n4705) );
  inv01 U3235 ( .Y(n4706), .A(n7809) );
  inv01 U3236 ( .Y(n4707), .A(n7429) );
  inv01 U3237 ( .Y(n4708), .A(n7808) );
  inv01 U3238 ( .Y(n4709), .A(n7423) );
  inv01 U3239 ( .Y(n4710), .A(n7807) );
  inv01 U3240 ( .Y(n4711), .A(n7409) );
  nand02 U3241 ( .Y(n4712), .A0(n4706), .A1(n4707) );
  nand02 U3242 ( .Y(n4713), .A0(n4708), .A1(n4709) );
  nand02 U3243 ( .Y(n4704), .A0(n4710), .A1(n4711) );
  nand02 U3244 ( .Y(n4714), .A0(n4712), .A1(n4713) );
  inv01 U3245 ( .Y(n4705), .A(n4714) );
  nand02 U3246 ( .Y(n2979), .A0(n4715), .A1(n4716) );
  inv01 U3247 ( .Y(n4717), .A(n7976) );
  inv01 U3248 ( .Y(n4718), .A(n7429) );
  inv01 U3249 ( .Y(n4719), .A(n7975) );
  inv01 U3250 ( .Y(n4720), .A(n7423) );
  inv01 U3251 ( .Y(n4721), .A(n7974) );
  inv01 U3252 ( .Y(n4722), .A(n7409) );
  nand02 U3253 ( .Y(n4723), .A0(n4717), .A1(n4718) );
  nand02 U3254 ( .Y(n4724), .A0(n4719), .A1(n4720) );
  nand02 U3255 ( .Y(n4715), .A0(n4721), .A1(n4722) );
  nand02 U3256 ( .Y(n4725), .A0(n4723), .A1(n4724) );
  inv01 U3257 ( .Y(n4716), .A(n4725) );
  inv01 U3258 ( .Y(n3021), .A(n4726) );
  nor02 U3259 ( .Y(n4727), .A0(n7428), .A1(n7762) );
  nor02 U3260 ( .Y(n4728), .A0(n7423), .A1(n7861) );
  nor02 U3261 ( .Y(n4729), .A0(n7409), .A1(n7860) );
  nor02 U3262 ( .Y(n4726), .A0(n4729), .A1(n4730) );
  nor02 U3263 ( .Y(n4731), .A0(n4727), .A1(n4728) );
  inv01 U3264 ( .Y(n4730), .A(n4731) );
  nand02 U3265 ( .Y(n3013), .A0(n4732), .A1(n4733) );
  inv01 U3266 ( .Y(n4734), .A(n7882) );
  inv01 U3267 ( .Y(n4735), .A(n7428) );
  inv01 U3268 ( .Y(n4736), .A(n7881) );
  inv01 U3269 ( .Y(n4737), .A(n7425) );
  inv01 U3270 ( .Y(n4738), .A(n7880) );
  inv01 U3271 ( .Y(n4739), .A(n7407) );
  nand02 U3272 ( .Y(n4740), .A0(n4734), .A1(n4735) );
  nand02 U3273 ( .Y(n4741), .A0(n4736), .A1(n4737) );
  nand02 U3274 ( .Y(n4732), .A0(n4738), .A1(n4739) );
  nand02 U3275 ( .Y(n4742), .A0(n4740), .A1(n4741) );
  inv01 U3276 ( .Y(n4733), .A(n4742) );
  nand02 U3277 ( .Y(n3022), .A0(n4743), .A1(n4744) );
  inv01 U3278 ( .Y(n4745), .A(n7763) );
  inv01 U3279 ( .Y(n4746), .A(n7429) );
  inv01 U3280 ( .Y(n4747), .A(n7859) );
  inv01 U3281 ( .Y(n4748), .A(n7425) );
  inv01 U3282 ( .Y(n4749), .A(n7858) );
  inv01 U3283 ( .Y(n4750), .A(n7407) );
  nand02 U3284 ( .Y(n4751), .A0(n4745), .A1(n4746) );
  nand02 U3285 ( .Y(n4752), .A0(n4747), .A1(n4748) );
  nand02 U3286 ( .Y(n4743), .A0(n4749), .A1(n4750) );
  nand02 U3287 ( .Y(n4753), .A0(n4751), .A1(n4752) );
  inv01 U3288 ( .Y(n4744), .A(n4753) );
  inv01 U3289 ( .Y(n2998), .A(n4754) );
  nor02 U3290 ( .Y(n4755), .A0(n7429), .A1(n7737) );
  nor02 U3291 ( .Y(n4756), .A0(n7425), .A1(n7919) );
  nor02 U3292 ( .Y(n4757), .A0(n7407), .A1(n7918) );
  nor02 U3293 ( .Y(n4754), .A0(n4757), .A1(n4758) );
  nor02 U3294 ( .Y(n4759), .A0(n4755), .A1(n4756) );
  inv01 U3295 ( .Y(n4758), .A(n4759) );
  nand02 U3296 ( .Y(n3005), .A0(n4760), .A1(n4761) );
  inv01 U3297 ( .Y(n4762), .A(n7732) );
  inv01 U3298 ( .Y(n4763), .A(n7427) );
  inv01 U3299 ( .Y(n4764), .A(n7901) );
  inv01 U3300 ( .Y(n4765), .A(n7424) );
  inv01 U3301 ( .Y(n4766), .A(n7900) );
  inv01 U3302 ( .Y(n4767), .A(n7408) );
  nand02 U3303 ( .Y(n4768), .A0(n4762), .A1(n4763) );
  nand02 U3304 ( .Y(n4769), .A0(n4764), .A1(n4765) );
  nand02 U3305 ( .Y(n4760), .A0(n4766), .A1(n4767) );
  nand02 U3306 ( .Y(n4770), .A0(n4768), .A1(n4769) );
  inv01 U3307 ( .Y(n4761), .A(n4770) );
  nand02 U3308 ( .Y(n3008), .A0(n4771), .A1(n4772) );
  inv01 U3309 ( .Y(n4773), .A(n7894) );
  inv01 U3310 ( .Y(n4774), .A(n7428) );
  inv01 U3311 ( .Y(n4775), .A(n7893) );
  inv01 U3312 ( .Y(n4776), .A(n7424) );
  inv01 U3313 ( .Y(n4777), .A(n7892) );
  inv01 U3314 ( .Y(n4778), .A(n7408) );
  nand02 U3315 ( .Y(n4779), .A0(n4773), .A1(n4774) );
  nand02 U3316 ( .Y(n4780), .A0(n4775), .A1(n4776) );
  nand02 U3317 ( .Y(n4771), .A0(n4777), .A1(n4778) );
  nand02 U3318 ( .Y(n4781), .A0(n4779), .A1(n4780) );
  inv01 U3319 ( .Y(n4772), .A(n4781) );
  inv01 U3320 ( .Y(n2981), .A(n4782) );
  nor02 U3321 ( .Y(n4783), .A0(n7428), .A1(n7970) );
  nor02 U3322 ( .Y(n4784), .A0(n7424), .A1(n7969) );
  nor02 U3323 ( .Y(n4785), .A0(n7408), .A1(n7968) );
  nor02 U3324 ( .Y(n4782), .A0(n4785), .A1(n4786) );
  nor02 U3325 ( .Y(n4787), .A0(n4783), .A1(n4784) );
  inv01 U3326 ( .Y(n4786), .A(n4787) );
  nand02 U3327 ( .Y(n3039), .A0(n4788), .A1(n4789) );
  inv01 U3328 ( .Y(n4790), .A(n7743) );
  inv01 U3329 ( .Y(n4791), .A(n7428) );
  inv01 U3330 ( .Y(n4792), .A(n7815) );
  inv01 U3331 ( .Y(n4793), .A(n7423) );
  inv01 U3332 ( .Y(n4794), .A(n7814) );
  inv01 U3333 ( .Y(n4795), .A(n7409) );
  nand02 U3334 ( .Y(n4796), .A0(n4790), .A1(n4791) );
  nand02 U3335 ( .Y(n4797), .A0(n4792), .A1(n4793) );
  nand02 U3336 ( .Y(n4788), .A0(n4794), .A1(n4795) );
  nand02 U3337 ( .Y(n4798), .A0(n4796), .A1(n4797) );
  inv01 U3338 ( .Y(n4789), .A(n4798) );
  nand02 U3339 ( .Y(n2973), .A0(n4799), .A1(n4800) );
  inv01 U3340 ( .Y(n4801), .A(n7994) );
  inv01 U3341 ( .Y(n4802), .A(n7429) );
  inv01 U3342 ( .Y(n4803), .A(n7993) );
  inv01 U3343 ( .Y(n4804), .A(n7423) );
  inv01 U3344 ( .Y(n4805), .A(n7992) );
  inv01 U3345 ( .Y(n4806), .A(n7409) );
  nand02 U3346 ( .Y(n4807), .A0(n4801), .A1(n4802) );
  nand02 U3347 ( .Y(n4808), .A0(n4803), .A1(n4804) );
  nand02 U3348 ( .Y(n4799), .A0(n4805), .A1(n4806) );
  nand02 U3349 ( .Y(n4809), .A0(n4807), .A1(n4808) );
  inv01 U3350 ( .Y(n4800), .A(n4809) );
  inv01 U3351 ( .Y(n3027), .A(n4810) );
  nor02 U3352 ( .Y(n4811), .A0(n7429), .A1(n7846) );
  nor02 U3353 ( .Y(n4812), .A0(n7423), .A1(n7845) );
  nor02 U3354 ( .Y(n4813), .A0(n7409), .A1(n7844) );
  nor02 U3355 ( .Y(n4810), .A0(n4813), .A1(n4814) );
  nor02 U3356 ( .Y(n4815), .A0(n4811), .A1(n4812) );
  inv01 U3357 ( .Y(n4814), .A(n4815) );
  nand02 U3358 ( .Y(n2992), .A0(n4816), .A1(n4817) );
  inv01 U3359 ( .Y(n4818), .A(n7937) );
  inv01 U3360 ( .Y(n4819), .A(n7427) );
  inv01 U3361 ( .Y(n4820), .A(n7936) );
  inv01 U3362 ( .Y(n4821), .A(n7425) );
  inv01 U3363 ( .Y(n4822), .A(n7935) );
  inv01 U3364 ( .Y(n4823), .A(n7407) );
  nand02 U3365 ( .Y(n4824), .A0(n4818), .A1(n4819) );
  nand02 U3366 ( .Y(n4825), .A0(n4820), .A1(n4821) );
  nand02 U3367 ( .Y(n4816), .A0(n4822), .A1(n4823) );
  nand02 U3368 ( .Y(n4826), .A0(n4824), .A1(n4825) );
  inv01 U3369 ( .Y(n4817), .A(n4826) );
  inv01 U3370 ( .Y(n3031), .A(n4827) );
  nor02 U3371 ( .Y(n4828), .A0(n7428), .A1(n7836) );
  nor02 U3372 ( .Y(n4829), .A0(n7425), .A1(n7835) );
  nor02 U3373 ( .Y(n4830), .A0(n7407), .A1(n7834) );
  nor02 U3374 ( .Y(n4827), .A0(n4830), .A1(n4831) );
  nor02 U3375 ( .Y(n4832), .A0(n4828), .A1(n4829) );
  inv01 U3376 ( .Y(n4831), .A(n4832) );
  nand02 U3377 ( .Y(n3047), .A0(n4833), .A1(n4834) );
  inv01 U3378 ( .Y(n4835), .A(n7758) );
  inv01 U3379 ( .Y(n4836), .A(n7429) );
  inv01 U3380 ( .Y(n4837), .A(n7795) );
  inv01 U3381 ( .Y(n4838), .A(n7424) );
  inv01 U3382 ( .Y(n4839), .A(n7794) );
  inv01 U3383 ( .Y(n4840), .A(n7408) );
  nand02 U3384 ( .Y(n4841), .A0(n4835), .A1(n4836) );
  nand02 U3385 ( .Y(n4842), .A0(n4837), .A1(n4838) );
  nand02 U3386 ( .Y(n4833), .A0(n4839), .A1(n4840) );
  nand02 U3387 ( .Y(n4843), .A0(n4841), .A1(n4842) );
  inv01 U3388 ( .Y(n4834), .A(n4843) );
  inv01 U3389 ( .Y(n3041), .A(n4844) );
  nor02 U3390 ( .Y(n4845), .A0(n7427), .A1(n7742) );
  nor02 U3391 ( .Y(n4846), .A0(n7424), .A1(n7811) );
  nor02 U3392 ( .Y(n4847), .A0(n7408), .A1(n7810) );
  nor02 U3393 ( .Y(n4844), .A0(n4847), .A1(n4848) );
  nor02 U3394 ( .Y(n4849), .A0(n4845), .A1(n4846) );
  inv01 U3395 ( .Y(n4848), .A(n4849) );
  inv01 U3396 ( .Y(n2986), .A(n4850) );
  nor02 U3397 ( .Y(n4851), .A0(n7427), .A1(n7955) );
  nor02 U3398 ( .Y(n4852), .A0(n7425), .A1(n7954) );
  nor02 U3399 ( .Y(n4853), .A0(n7407), .A1(n7953) );
  nor02 U3400 ( .Y(n4850), .A0(n4853), .A1(n4854) );
  nor02 U3401 ( .Y(n4855), .A0(n4851), .A1(n4852) );
  inv01 U3402 ( .Y(n4854), .A(n4855) );
  nand02 U3403 ( .Y(n2994), .A0(n4856), .A1(n4857) );
  inv01 U3404 ( .Y(n4858), .A(n7931) );
  inv01 U3405 ( .Y(n4859), .A(n7429) );
  inv01 U3406 ( .Y(n4860), .A(n7930) );
  inv01 U3407 ( .Y(n4861), .A(n7423) );
  inv01 U3408 ( .Y(n4862), .A(n7929) );
  inv01 U3409 ( .Y(n4863), .A(n7409) );
  nand02 U3410 ( .Y(n4864), .A0(n4858), .A1(n4859) );
  nand02 U3411 ( .Y(n4865), .A0(n4860), .A1(n4861) );
  nand02 U3412 ( .Y(n4856), .A0(n4862), .A1(n4863) );
  nand02 U3413 ( .Y(n4866), .A0(n4864), .A1(n4865) );
  inv01 U3414 ( .Y(n4857), .A(n4866) );
  inv01 U3415 ( .Y(n2985), .A(n4867) );
  nor02 U3416 ( .Y(n4868), .A0(n7429), .A1(n7958) );
  nor02 U3417 ( .Y(n4869), .A0(n7423), .A1(n7957) );
  nor02 U3418 ( .Y(n4870), .A0(n7409), .A1(n7956) );
  nor02 U3419 ( .Y(n4867), .A0(n4870), .A1(n4871) );
  nor02 U3420 ( .Y(n4872), .A0(n4868), .A1(n4869) );
  inv01 U3421 ( .Y(n4871), .A(n4872) );
  nand02 U3422 ( .Y(n3014), .A0(n4873), .A1(n4874) );
  inv01 U3423 ( .Y(n4875), .A(n7879) );
  inv01 U3424 ( .Y(n4876), .A(n7427) );
  inv01 U3425 ( .Y(n4877), .A(n7878) );
  inv01 U3426 ( .Y(n4878), .A(n7424) );
  inv01 U3427 ( .Y(n4879), .A(n7877) );
  inv01 U3428 ( .Y(n4880), .A(n7408) );
  nand02 U3429 ( .Y(n4881), .A0(n4875), .A1(n4876) );
  nand02 U3430 ( .Y(n4882), .A0(n4877), .A1(n4878) );
  nand02 U3431 ( .Y(n4873), .A0(n4879), .A1(n4880) );
  nand02 U3432 ( .Y(n4883), .A0(n4881), .A1(n4882) );
  inv01 U3433 ( .Y(n4874), .A(n4883) );
  nand02 U3434 ( .Y(n3023), .A0(n4884), .A1(n4885) );
  inv01 U3435 ( .Y(n4886), .A(n7761) );
  inv01 U3436 ( .Y(n4887), .A(n7427) );
  inv01 U3437 ( .Y(n4888), .A(n7857) );
  inv01 U3438 ( .Y(n4889), .A(n7424) );
  inv01 U3439 ( .Y(n4890), .A(n7856) );
  inv01 U3440 ( .Y(n4891), .A(n7408) );
  nand02 U3441 ( .Y(n4892), .A0(n4886), .A1(n4887) );
  nand02 U3442 ( .Y(n4893), .A0(n4888), .A1(n4889) );
  nand02 U3443 ( .Y(n4884), .A0(n4890), .A1(n4891) );
  nand02 U3444 ( .Y(n4894), .A0(n4892), .A1(n4893) );
  inv01 U3445 ( .Y(n4885), .A(n4894) );
  inv01 U3446 ( .Y(n2975), .A(n4895) );
  nor02 U3447 ( .Y(n4896), .A0(n7428), .A1(n7988) );
  nor02 U3448 ( .Y(n4897), .A0(n7424), .A1(n7987) );
  nor02 U3449 ( .Y(n4898), .A0(n7408), .A1(n7986) );
  nor02 U3450 ( .Y(n4895), .A0(n4898), .A1(n4899) );
  nor02 U3451 ( .Y(n4900), .A0(n4896), .A1(n4897) );
  inv01 U3452 ( .Y(n4899), .A(n4900) );
  nand02 U3453 ( .Y(n3019), .A0(n4901), .A1(n4902) );
  inv01 U3454 ( .Y(n4903), .A(n7867) );
  inv01 U3455 ( .Y(n4904), .A(n7429) );
  inv01 U3456 ( .Y(n4905), .A(n7866) );
  inv01 U3457 ( .Y(n4906), .A(n7425) );
  inv01 U3458 ( .Y(n4907), .A(n7865) );
  inv01 U3459 ( .Y(n4908), .A(n7407) );
  nand02 U3460 ( .Y(n4909), .A0(n4903), .A1(n4904) );
  nand02 U3461 ( .Y(n4910), .A0(n4905), .A1(n4906) );
  nand02 U3462 ( .Y(n4901), .A0(n4907), .A1(n4908) );
  nand02 U3463 ( .Y(n4911), .A0(n4909), .A1(n4910) );
  inv01 U3464 ( .Y(n4902), .A(n4911) );
  nand02 U3465 ( .Y(n3040), .A0(n4912), .A1(n4913) );
  inv01 U3466 ( .Y(n4914), .A(n7744) );
  inv01 U3467 ( .Y(n4915), .A(n7429) );
  inv01 U3468 ( .Y(n4916), .A(n7813) );
  inv01 U3469 ( .Y(n4917), .A(n7425) );
  inv01 U3470 ( .Y(n4918), .A(n7812) );
  inv01 U3471 ( .Y(n4919), .A(n7407) );
  nand02 U3472 ( .Y(n4920), .A0(n4914), .A1(n4915) );
  nand02 U3473 ( .Y(n4921), .A0(n4916), .A1(n4917) );
  nand02 U3474 ( .Y(n4912), .A0(n4918), .A1(n4919) );
  nand02 U3475 ( .Y(n4922), .A0(n4920), .A1(n4921) );
  inv01 U3476 ( .Y(n4913), .A(n4922) );
  inv01 U3477 ( .Y(n3028), .A(n4923) );
  nor02 U3478 ( .Y(n4924), .A0(n7428), .A1(n7757) );
  nor02 U3479 ( .Y(n4925), .A0(n7425), .A1(n7843) );
  nor02 U3480 ( .Y(n4926), .A0(n7407), .A1(n7842) );
  nor02 U3481 ( .Y(n4923), .A0(n4926), .A1(n4927) );
  nor02 U3482 ( .Y(n4928), .A0(n4924), .A1(n4925) );
  inv01 U3483 ( .Y(n4927), .A(n4928) );
  nand02 U3484 ( .Y(n3003), .A0(n4929), .A1(n4930) );
  inv01 U3485 ( .Y(n4931), .A(n7906) );
  inv01 U3486 ( .Y(n4932), .A(n7427) );
  inv01 U3487 ( .Y(n4933), .A(n7905) );
  inv01 U3488 ( .Y(n4934), .A(n7423) );
  inv01 U3489 ( .Y(n4935), .A(n7904) );
  inv01 U3490 ( .Y(n4936), .A(n7409) );
  nand02 U3491 ( .Y(n4937), .A0(n4931), .A1(n4932) );
  nand02 U3492 ( .Y(n4938), .A0(n4933), .A1(n4934) );
  nand02 U3493 ( .Y(n4929), .A0(n4935), .A1(n4936) );
  nand02 U3494 ( .Y(n4939), .A0(n4937), .A1(n4938) );
  inv01 U3495 ( .Y(n4930), .A(n4939) );
  nand02 U3496 ( .Y(n2997), .A0(n4940), .A1(n4941) );
  inv01 U3497 ( .Y(n4942), .A(n7922) );
  inv01 U3498 ( .Y(n4943), .A(n7428) );
  inv01 U3499 ( .Y(n4944), .A(n7921) );
  inv01 U3500 ( .Y(n4945), .A(n7423) );
  inv01 U3501 ( .Y(n4946), .A(n7920) );
  inv01 U3502 ( .Y(n4947), .A(n7409) );
  nand02 U3503 ( .Y(n4948), .A0(n4942), .A1(n4943) );
  nand02 U3504 ( .Y(n4949), .A0(n4944), .A1(n4945) );
  nand02 U3505 ( .Y(n4940), .A0(n4946), .A1(n4947) );
  nand02 U3506 ( .Y(n4950), .A0(n4948), .A1(n4949) );
  inv01 U3507 ( .Y(n4941), .A(n4950) );
  inv01 U3508 ( .Y(n3009), .A(n4951) );
  nor02 U3509 ( .Y(n4952), .A0(n7427), .A1(n7725) );
  nor02 U3510 ( .Y(n4953), .A0(n7423), .A1(n7891) );
  nor02 U3511 ( .Y(n4954), .A0(n7409), .A1(n7890) );
  nor02 U3512 ( .Y(n4951), .A0(n4954), .A1(n4955) );
  nor02 U3513 ( .Y(n4956), .A0(n4952), .A1(n4953) );
  inv01 U3514 ( .Y(n4955), .A(n4956) );
  inv02 U3515 ( .Y(n6835), .A(n6834) );
  inv02 U3516 ( .Y(n6855), .A(n6854) );
  inv02 U3517 ( .Y(n6875), .A(n6874) );
  inv02 U3518 ( .Y(n6893), .A(n6892) );
  inv02 U3519 ( .Y(n6879), .A(n6878) );
  inv02 U3520 ( .Y(n6849), .A(n6848) );
  inv02 U3521 ( .Y(n6873), .A(n6872) );
  inv02 U3522 ( .Y(n6843), .A(n6842) );
  inv02 U3523 ( .Y(n6887), .A(n6886) );
  inv02 U3524 ( .Y(n6891), .A(n6890) );
  inv02 U3525 ( .Y(n6831), .A(n6830) );
  inv02 U3526 ( .Y(n6845), .A(n6844) );
  inv02 U3527 ( .Y(n6847), .A(n6846) );
  inv02 U3528 ( .Y(n6883), .A(n6882) );
  inv02 U3529 ( .Y(n6869), .A(n6868) );
  inv02 U3530 ( .Y(n6837), .A(n6836) );
  inv02 U3531 ( .Y(n6881), .A(n6880) );
  inv02 U3532 ( .Y(n6851), .A(n6850) );
  inv02 U3533 ( .Y(n6877), .A(n6876) );
  inv02 U3534 ( .Y(n6889), .A(n6888) );
  inv02 U3535 ( .Y(n6839), .A(n6838) );
  inv02 U3536 ( .Y(n6853), .A(n6852) );
  inv02 U3537 ( .Y(n7167), .A(n7166) );
  inv02 U3538 ( .Y(n7165), .A(n7590) );
  inv02 U3539 ( .Y(n7211), .A(n7598) );
  inv02 U3540 ( .Y(n6885), .A(n6884) );
  inv02 U3541 ( .Y(n6833), .A(n6832) );
  inv02 U3542 ( .Y(n7208), .A(n7607) );
  inv02 U3543 ( .Y(n7205), .A(n7613) );
  inv02 U3544 ( .Y(n7200), .A(n7612) );
  inv02 U3545 ( .Y(n6841), .A(n6840) );
  inv02 U3546 ( .Y(n7206), .A(n7616) );
  inv02 U3547 ( .Y(n7201), .A(n7620) );
  inv02 U3548 ( .Y(n6871), .A(n6870) );
  inv02 U3549 ( .Y(n7204), .A(n7623) );
  inv02 U3550 ( .Y(n7187), .A(n7625) );
  inv02 U3551 ( .Y(n7207), .A(n7629) );
  inv02 U3552 ( .Y(n7210), .A(n7632) );
  buf02 U3553 ( .Y(n7203), .A(r0_11_) );
  inv02 U3554 ( .Y(n7209), .A(n7644) );
  inv02 U3555 ( .Y(n7213), .A(n7654) );
  inv02 U3556 ( .Y(n7214), .A(n7656) );
  inv02 U3557 ( .Y(n7202), .A(n7647) );
  inv02 U3558 ( .Y(n7186), .A(n7646) );
  inv02 U3559 ( .Y(n7212), .A(n7649) );
  inv02 U3560 ( .Y(n7125), .A(n7124) );
  inv02 U3561 ( .Y(n7123), .A(n7642) );
  inv02 U3562 ( .Y(n7121), .A(n7120) );
  inv02 U3563 ( .Y(result407_50_), .A(n7022) );
  inv02 U3564 ( .Y(s_op2_49_), .A(n6998) );
  inv02 U3565 ( .Y(s_op2_46_), .A(n7058) );
  inv02 U3566 ( .Y(s_op2_43_), .A(n6980) );
  inv02 U3567 ( .Y(s_op2_42_), .A(n6974) );
  inv02 U3568 ( .Y(s_op2_23_), .A(n7064) );
  inv02 U3569 ( .Y(s_op2_21_), .A(n7070) );
  inv04 U3570 ( .Y(n7164), .A(n7652) );
  inv01 U3571 ( .Y(n2907), .A(n4957) );
  nor02 U3572 ( .Y(n4958), .A0(n7433), .A1(n2763) );
  nor02 U3573 ( .Y(n4959), .A0(n7889), .A1(n7412) );
  nor02 U3574 ( .Y(n4960), .A0(n7888), .A1(n7417) );
  nor02 U3575 ( .Y(n4957), .A0(n4960), .A1(n4961) );
  nor02 U3576 ( .Y(n4962), .A0(n4958), .A1(n4959) );
  inv01 U3577 ( .Y(n4961), .A(n4962) );
  inv01 U3578 ( .Y(n2876), .A(n4963) );
  nor02 U3579 ( .Y(n4964), .A0(n7616), .A1(n7432) );
  nor02 U3580 ( .Y(n4965), .A0(n7975), .A1(n7413) );
  nor02 U3581 ( .Y(n4966), .A0(n7974), .A1(n7415) );
  nor02 U3582 ( .Y(n4963), .A0(n4966), .A1(n4967) );
  nor02 U3583 ( .Y(n4968), .A0(n4964), .A1(n4965) );
  inv01 U3584 ( .Y(n4967), .A(n4968) );
  inv01 U3585 ( .Y(n2868), .A(n4969) );
  nor02 U3586 ( .Y(n4970), .A0(n7578), .A1(n7433) );
  nor02 U3587 ( .Y(n4971), .A0(n7999), .A1(n7412) );
  nor02 U3588 ( .Y(n4972), .A0(n7998), .A1(n7417) );
  nor02 U3589 ( .Y(n4969), .A0(n4972), .A1(n4973) );
  nor02 U3590 ( .Y(n4974), .A0(n4970), .A1(n4971) );
  inv01 U3591 ( .Y(n4973), .A(n4974) );
  inv01 U3592 ( .Y(n2927), .A(n4975) );
  nor02 U3593 ( .Y(n4976), .A0(n7432), .A1(n2741) );
  nor02 U3594 ( .Y(n4977), .A0(n7838), .A1(n7413) );
  nor02 U3595 ( .Y(n4978), .A0(n7837), .A1(n7415) );
  nor02 U3596 ( .Y(n4975), .A0(n4978), .A1(n4979) );
  nor02 U3597 ( .Y(n4980), .A0(n4976), .A1(n4977) );
  inv01 U3598 ( .Y(n4979), .A(n4980) );
  inv01 U3599 ( .Y(n2899), .A(n4981) );
  nor02 U3600 ( .Y(n4982), .A0(n7431), .A1(n2772) );
  nor02 U3601 ( .Y(n4983), .A0(n7908), .A1(n7411) );
  nor02 U3602 ( .Y(n4984), .A0(n7907), .A1(n7416) );
  nor02 U3603 ( .Y(n4981), .A0(n4984), .A1(n4985) );
  nor02 U3604 ( .Y(n4986), .A0(n4982), .A1(n4983) );
  inv01 U3605 ( .Y(n4985), .A(n4986) );
  inv01 U3606 ( .Y(n2928), .A(n4987) );
  nor02 U3607 ( .Y(n4988), .A0(n7432), .A1(n2740) );
  nor02 U3608 ( .Y(n4989), .A0(n7835), .A1(n7412) );
  nor02 U3609 ( .Y(n4990), .A0(n7834), .A1(n7417) );
  nor02 U3610 ( .Y(n4987), .A0(n4990), .A1(n4991) );
  nor02 U3611 ( .Y(n4992), .A0(n4988), .A1(n4989) );
  inv01 U3612 ( .Y(n4991), .A(n4992) );
  inv01 U3613 ( .Y(n2878), .A(n4993) );
  nor02 U3614 ( .Y(n4994), .A0(n7623), .A1(n7432) );
  nor02 U3615 ( .Y(n4995), .A0(n7969), .A1(n7411) );
  nor02 U3616 ( .Y(n4996), .A0(n7968), .A1(n7416) );
  nor02 U3617 ( .Y(n4993), .A0(n4996), .A1(n4997) );
  nor02 U3618 ( .Y(n4998), .A0(n4994), .A1(n4995) );
  inv01 U3619 ( .Y(n4997), .A(n4998) );
  inv01 U3620 ( .Y(n2902), .A(n4999) );
  nor02 U3621 ( .Y(n5000), .A0(n7431), .A1(n2769) );
  nor02 U3622 ( .Y(n5001), .A0(n7901), .A1(n7411) );
  nor02 U3623 ( .Y(n5002), .A0(n7900), .A1(n7416) );
  nor02 U3624 ( .Y(n4999), .A0(n5002), .A1(n5003) );
  nor02 U3625 ( .Y(n5004), .A0(n5000), .A1(n5001) );
  inv01 U3626 ( .Y(n5003), .A(n5004) );
  inv01 U3627 ( .Y(n2922), .A(n5005) );
  nor02 U3628 ( .Y(n5006), .A0(n7431), .A1(n2747) );
  nor02 U3629 ( .Y(n5007), .A0(n7851), .A1(n7412) );
  nor02 U3630 ( .Y(n5008), .A0(n7850), .A1(n7417) );
  nor02 U3631 ( .Y(n5005), .A0(n5008), .A1(n5009) );
  nor02 U3632 ( .Y(n5010), .A0(n5006), .A1(n5007) );
  inv01 U3633 ( .Y(n5009), .A(n5010) );
  inv01 U3634 ( .Y(n2888), .A(n5011) );
  nor02 U3635 ( .Y(n5012), .A0(n7649), .A1(n7433) );
  nor02 U3636 ( .Y(n5013), .A0(n7939), .A1(n7413) );
  nor02 U3637 ( .Y(n5014), .A0(n7938), .A1(n7415) );
  nor02 U3638 ( .Y(n5011), .A0(n5014), .A1(n5015) );
  nor02 U3639 ( .Y(n5016), .A0(n5012), .A1(n5013) );
  inv01 U3640 ( .Y(n5015), .A(n5016) );
  inv01 U3641 ( .Y(n2915), .A(n5017) );
  nor02 U3642 ( .Y(n5018), .A0(n7433), .A1(n2755) );
  nor02 U3643 ( .Y(n5019), .A0(n7869), .A1(n7413) );
  nor02 U3644 ( .Y(n5020), .A0(n7868), .A1(n7415) );
  nor02 U3645 ( .Y(n5017), .A0(n5020), .A1(n5021) );
  nor02 U3646 ( .Y(n5022), .A0(n5018), .A1(n5019) );
  inv01 U3647 ( .Y(n5021), .A(n5022) );
  inv01 U3648 ( .Y(n2894), .A(n5023) );
  nor02 U3649 ( .Y(n5024), .A0(n7433), .A1(n2778) );
  nor02 U3650 ( .Y(n5025), .A0(n7921), .A1(n7413) );
  nor02 U3651 ( .Y(n5026), .A0(n7920), .A1(n7415) );
  nor02 U3652 ( .Y(n5023), .A0(n5026), .A1(n5027) );
  nor02 U3653 ( .Y(n5028), .A0(n5024), .A1(n5025) );
  inv01 U3654 ( .Y(n5027), .A(n5028) );
  inv01 U3655 ( .Y(n2920), .A(n5029) );
  nor02 U3656 ( .Y(n5030), .A0(n7431), .A1(n2749) );
  nor02 U3657 ( .Y(n5031), .A0(n7857), .A1(n7411) );
  nor02 U3658 ( .Y(n5032), .A0(n7856), .A1(n7416) );
  nor02 U3659 ( .Y(n5029), .A0(n5032), .A1(n5033) );
  nor02 U3660 ( .Y(n5034), .A0(n5030), .A1(n5031) );
  inv01 U3661 ( .Y(n5033), .A(n5034) );
  inv01 U3662 ( .Y(n2929), .A(n5035) );
  nor02 U3663 ( .Y(n5036), .A0(n7433), .A1(n2739) );
  nor02 U3664 ( .Y(n5037), .A0(n7832), .A1(n7411) );
  nor02 U3665 ( .Y(n5038), .A0(n7831), .A1(n7416) );
  nor02 U3666 ( .Y(n5035), .A0(n5038), .A1(n5039) );
  nor02 U3667 ( .Y(n5040), .A0(n5036), .A1(n5037) );
  inv01 U3668 ( .Y(n5039), .A(n5040) );
  inv01 U3669 ( .Y(n2914), .A(n5041) );
  nor02 U3670 ( .Y(n5042), .A0(n7433), .A1(n2756) );
  nor02 U3671 ( .Y(n5043), .A0(n7871), .A1(n7411) );
  nor02 U3672 ( .Y(n5044), .A0(n7870), .A1(n7416) );
  nor02 U3673 ( .Y(n5041), .A0(n5044), .A1(n5045) );
  nor02 U3674 ( .Y(n5046), .A0(n5042), .A1(n5043) );
  inv01 U3675 ( .Y(n5045), .A(n5046) );
  inv01 U3676 ( .Y(n2903), .A(n5047) );
  nor02 U3677 ( .Y(n5048), .A0(n7433), .A1(n2768) );
  nor02 U3678 ( .Y(n5049), .A0(n7899), .A1(n7413) );
  nor02 U3679 ( .Y(n5050), .A0(n7898), .A1(n7415) );
  nor02 U3680 ( .Y(n5047), .A0(n5050), .A1(n5051) );
  nor02 U3681 ( .Y(n5052), .A0(n5048), .A1(n5049) );
  inv01 U3682 ( .Y(n5051), .A(n5052) );
  inv01 U3683 ( .Y(n2881), .A(n5053) );
  nor02 U3684 ( .Y(n5054), .A0(n7632), .A1(n7431) );
  nor02 U3685 ( .Y(n5055), .A0(n7960), .A1(n7411) );
  nor02 U3686 ( .Y(n5056), .A0(n7959), .A1(n7416) );
  nor02 U3687 ( .Y(n5053), .A0(n5056), .A1(n5057) );
  nor02 U3688 ( .Y(n5058), .A0(n5054), .A1(n5055) );
  inv01 U3689 ( .Y(n5057), .A(n5058) );
  inv01 U3690 ( .Y(n2912), .A(n5059) );
  nor02 U3691 ( .Y(n5060), .A0(n7432), .A1(n2758) );
  nor02 U3692 ( .Y(n5061), .A0(n7875), .A1(n7413) );
  nor02 U3693 ( .Y(n5062), .A0(n7874), .A1(n7415) );
  nor02 U3694 ( .Y(n5059), .A0(n5062), .A1(n5063) );
  nor02 U3695 ( .Y(n5064), .A0(n5060), .A1(n5061) );
  inv01 U3696 ( .Y(n5063), .A(n5064) );
  inv01 U3697 ( .Y(n2895), .A(n5065) );
  nor02 U3698 ( .Y(n5066), .A0(n7433), .A1(n2777) );
  nor02 U3699 ( .Y(n5067), .A0(n7919), .A1(n7412) );
  nor02 U3700 ( .Y(n5068), .A0(n7918), .A1(n7417) );
  nor02 U3701 ( .Y(n5065), .A0(n5068), .A1(n5069) );
  nor02 U3702 ( .Y(n5070), .A0(n5066), .A1(n5067) );
  inv01 U3703 ( .Y(n5069), .A(n5070) );
  inv01 U3704 ( .Y(n2913), .A(n5071) );
  nor02 U3705 ( .Y(n5072), .A0(n7433), .A1(n2757) );
  nor02 U3706 ( .Y(n5073), .A0(n7873), .A1(n7412) );
  nor02 U3707 ( .Y(n5074), .A0(n7872), .A1(n7417) );
  nor02 U3708 ( .Y(n5071), .A0(n5074), .A1(n5075) );
  nor02 U3709 ( .Y(n5076), .A0(n5072), .A1(n5073) );
  inv01 U3710 ( .Y(n5075), .A(n5076) );
  inv01 U3711 ( .Y(n2909), .A(n5077) );
  nor02 U3712 ( .Y(n5078), .A0(n7431), .A1(n2761) );
  nor02 U3713 ( .Y(n5079), .A0(n7884), .A1(n7413) );
  nor02 U3714 ( .Y(n5080), .A0(n7883), .A1(n7415) );
  nor02 U3715 ( .Y(n5077), .A0(n5080), .A1(n5081) );
  nor02 U3716 ( .Y(n5082), .A0(n5078), .A1(n5079) );
  inv01 U3717 ( .Y(n5081), .A(n5082) );
  inv01 U3718 ( .Y(n2923), .A(n5083) );
  nor02 U3719 ( .Y(n5084), .A0(n7431), .A1(n2746) );
  nor02 U3720 ( .Y(n5085), .A0(n7848), .A1(n7411) );
  nor02 U3721 ( .Y(n5086), .A0(n7847), .A1(n7416) );
  nor02 U3722 ( .Y(n5083), .A0(n5086), .A1(n5087) );
  nor02 U3723 ( .Y(n5088), .A0(n5084), .A1(n5085) );
  inv01 U3724 ( .Y(n5087), .A(n5088) );
  inv01 U3725 ( .Y(n2886), .A(n5089) );
  nor02 U3726 ( .Y(n5090), .A0(n7647), .A1(n7431) );
  nor02 U3727 ( .Y(n5091), .A0(n7945), .A1(n7412) );
  nor02 U3728 ( .Y(n5092), .A0(n7944), .A1(n7417) );
  nor02 U3729 ( .Y(n5089), .A0(n5092), .A1(n5093) );
  nor02 U3730 ( .Y(n5094), .A0(n5090), .A1(n5091) );
  inv01 U3731 ( .Y(n5093), .A(n5094) );
  inv01 U3732 ( .Y(n2935), .A(n5095) );
  nor02 U3733 ( .Y(n5096), .A0(n7432), .A1(n2733) );
  nor02 U3734 ( .Y(n5097), .A0(n7817), .A1(n7411) );
  nor02 U3735 ( .Y(n5098), .A0(n7816), .A1(n7416) );
  nor02 U3736 ( .Y(n5095), .A0(n5098), .A1(n5099) );
  nor02 U3737 ( .Y(n5100), .A0(n5096), .A1(n5097) );
  inv01 U3738 ( .Y(n5099), .A(n5100) );
  inv01 U3739 ( .Y(n2939), .A(n5101) );
  nor02 U3740 ( .Y(n5102), .A0(n7433), .A1(n2780) );
  nor02 U3741 ( .Y(n5103), .A0(n7808), .A1(n7413) );
  nor02 U3742 ( .Y(n5104), .A0(n7807), .A1(n7415) );
  nor02 U3743 ( .Y(n5101), .A0(n5104), .A1(n5105) );
  nor02 U3744 ( .Y(n5106), .A0(n5102), .A1(n5103) );
  inv01 U3745 ( .Y(n5105), .A(n5106) );
  inv01 U3746 ( .Y(n2883), .A(n5107) );
  nor02 U3747 ( .Y(n5108), .A0(n7644), .A1(n7431) );
  nor02 U3748 ( .Y(n5109), .A0(n7954), .A1(n7412) );
  nor02 U3749 ( .Y(n5110), .A0(n7953), .A1(n7417) );
  nor02 U3750 ( .Y(n5107), .A0(n5110), .A1(n5111) );
  nor02 U3751 ( .Y(n5112), .A0(n5108), .A1(n5109) );
  inv01 U3752 ( .Y(n5111), .A(n5112) );
  inv01 U3753 ( .Y(n2916), .A(n5113) );
  nor02 U3754 ( .Y(n5114), .A0(n7433), .A1(n2753) );
  nor02 U3755 ( .Y(n5115), .A0(n7866), .A1(n7412) );
  nor02 U3756 ( .Y(n5116), .A0(n7865), .A1(n7417) );
  nor02 U3757 ( .Y(n5113), .A0(n5116), .A1(n5117) );
  nor02 U3758 ( .Y(n5118), .A0(n5114), .A1(n5115) );
  inv01 U3759 ( .Y(n5117), .A(n5118) );
  inv01 U3760 ( .Y(n2921), .A(n5119) );
  nor02 U3761 ( .Y(n5120), .A0(n7432), .A1(n2748) );
  nor02 U3762 ( .Y(n5121), .A0(n7854), .A1(n7413) );
  nor02 U3763 ( .Y(n5122), .A0(n7853), .A1(n7415) );
  nor02 U3764 ( .Y(n5119), .A0(n5122), .A1(n5123) );
  nor02 U3765 ( .Y(n5124), .A0(n5120), .A1(n5121) );
  inv01 U3766 ( .Y(n5123), .A(n5124) );
  inv01 U3767 ( .Y(n2931), .A(n5125) );
  nor02 U3768 ( .Y(n5126), .A0(n7433), .A1(n2737) );
  nor02 U3769 ( .Y(n5127), .A0(n7828), .A1(n7412) );
  nor02 U3770 ( .Y(n5128), .A0(n7827), .A1(n7417) );
  nor02 U3771 ( .Y(n5125), .A0(n5128), .A1(n5129) );
  nor02 U3772 ( .Y(n5130), .A0(n5126), .A1(n5127) );
  inv01 U3773 ( .Y(n5129), .A(n5130) );
  inv01 U3774 ( .Y(n2872), .A(n5131) );
  nor02 U3775 ( .Y(n5132), .A0(n7598), .A1(n7433) );
  nor02 U3776 ( .Y(n5133), .A0(n7987), .A1(n7411) );
  nor02 U3777 ( .Y(n5134), .A0(n7986), .A1(n7416) );
  nor02 U3778 ( .Y(n5131), .A0(n5134), .A1(n5135) );
  nor02 U3779 ( .Y(n5136), .A0(n5132), .A1(n5133) );
  inv01 U3780 ( .Y(n5135), .A(n5136) );
  inv01 U3781 ( .Y(n2869), .A(n5137) );
  nor02 U3782 ( .Y(n5138), .A0(n7582), .A1(n7432) );
  nor02 U3783 ( .Y(n5139), .A0(n7996), .A1(n7411) );
  nor02 U3784 ( .Y(n5140), .A0(n7995), .A1(n7416) );
  nor02 U3785 ( .Y(n5137), .A0(n5140), .A1(n5141) );
  nor02 U3786 ( .Y(n5142), .A0(n5138), .A1(n5139) );
  inv01 U3787 ( .Y(n5141), .A(n5142) );
  inv01 U3788 ( .Y(n2917), .A(n5143) );
  nor02 U3789 ( .Y(n5144), .A0(n7433), .A1(n2752) );
  nor02 U3790 ( .Y(n5145), .A0(n7863), .A1(n7411) );
  nor02 U3791 ( .Y(n5146), .A0(n7862), .A1(n7416) );
  nor02 U3792 ( .Y(n5143), .A0(n5146), .A1(n5147) );
  nor02 U3793 ( .Y(n5148), .A0(n5144), .A1(n5145) );
  inv01 U3794 ( .Y(n5147), .A(n5148) );
  inv01 U3795 ( .Y(n2889), .A(n5149) );
  nor02 U3796 ( .Y(n5150), .A0(n7660), .A1(n7432) );
  nor02 U3797 ( .Y(n5151), .A0(n7936), .A1(n7412) );
  nor02 U3798 ( .Y(n5152), .A0(n7935), .A1(n7417) );
  nor02 U3799 ( .Y(n5149), .A0(n5152), .A1(n5153) );
  nor02 U3800 ( .Y(n5154), .A0(n5150), .A1(n5151) );
  inv01 U3801 ( .Y(n5153), .A(n5154) );
  inv01 U3802 ( .Y(n2879), .A(n5155) );
  nor02 U3803 ( .Y(n5156), .A0(n7625), .A1(n7431) );
  nor02 U3804 ( .Y(n5157), .A0(n7966), .A1(n7413) );
  nor02 U3805 ( .Y(n5158), .A0(n7965), .A1(n7415) );
  nor02 U3806 ( .Y(n5155), .A0(n5158), .A1(n5159) );
  nor02 U3807 ( .Y(n5160), .A0(n5156), .A1(n5157) );
  inv01 U3808 ( .Y(n5159), .A(n5160) );
  inv01 U3809 ( .Y(n2919), .A(n5161) );
  nor02 U3810 ( .Y(n5162), .A0(n7433), .A1(n2750) );
  nor02 U3811 ( .Y(n5163), .A0(n7859), .A1(n7412) );
  nor02 U3812 ( .Y(n5164), .A0(n7858), .A1(n7417) );
  nor02 U3813 ( .Y(n5161), .A0(n5164), .A1(n5165) );
  nor02 U3814 ( .Y(n5166), .A0(n5162), .A1(n5163) );
  inv01 U3815 ( .Y(n5165), .A(n5166) );
  inv01 U3816 ( .Y(n2871), .A(n5167) );
  nor02 U3817 ( .Y(n5168), .A0(n7590), .A1(n7431) );
  nor02 U3818 ( .Y(n5169), .A0(n7990), .A1(n7412) );
  nor02 U3819 ( .Y(n5170), .A0(n7989), .A1(n7417) );
  nor02 U3820 ( .Y(n5167), .A0(n5170), .A1(n5171) );
  nor02 U3821 ( .Y(n5172), .A0(n5168), .A1(n5169) );
  inv01 U3822 ( .Y(n5171), .A(n5172) );
  inv01 U3823 ( .Y(n2941), .A(n5173) );
  nor02 U3824 ( .Y(n5174), .A0(n7432), .A1(n2776) );
  nor02 U3825 ( .Y(n5175), .A0(n7803), .A1(n7411) );
  nor02 U3826 ( .Y(n5176), .A0(n7802), .A1(n7416) );
  nor02 U3827 ( .Y(n5173), .A0(n5176), .A1(n5177) );
  nor02 U3828 ( .Y(n5178), .A0(n5174), .A1(n5175) );
  inv01 U3829 ( .Y(n5177), .A(n5178) );
  inv01 U3830 ( .Y(n2900), .A(n5179) );
  nor02 U3831 ( .Y(n5180), .A0(n7431), .A1(n2771) );
  nor02 U3832 ( .Y(n5181), .A0(n7905), .A1(n7413) );
  nor02 U3833 ( .Y(n5182), .A0(n7904), .A1(n7415) );
  nor02 U3834 ( .Y(n5179), .A0(n5182), .A1(n5183) );
  nor02 U3835 ( .Y(n5184), .A0(n5180), .A1(n5181) );
  inv01 U3836 ( .Y(n5183), .A(n5184) );
  inv01 U3837 ( .Y(n2906), .A(n5185) );
  nor02 U3838 ( .Y(n5186), .A0(n7431), .A1(n2764) );
  nor02 U3839 ( .Y(n5187), .A0(n7891), .A1(n7413) );
  nor02 U3840 ( .Y(n5188), .A0(n7890), .A1(n7415) );
  nor02 U3841 ( .Y(n5185), .A0(n5188), .A1(n5189) );
  nor02 U3842 ( .Y(n5190), .A0(n5186), .A1(n5187) );
  inv01 U3843 ( .Y(n5189), .A(n5190) );
  inv01 U3844 ( .Y(n2877), .A(n5191) );
  nor02 U3845 ( .Y(n5192), .A0(n7620), .A1(n7431) );
  nor02 U3846 ( .Y(n5193), .A0(n7972), .A1(n7412) );
  nor02 U3847 ( .Y(n5194), .A0(n7971), .A1(n7417) );
  nor02 U3848 ( .Y(n5191), .A0(n5194), .A1(n5195) );
  nor02 U3849 ( .Y(n5196), .A0(n5192), .A1(n5193) );
  inv01 U3850 ( .Y(n5195), .A(n5196) );
  inv01 U3851 ( .Y(n2898), .A(n5197) );
  nor02 U3852 ( .Y(n5198), .A0(n7433), .A1(n2773) );
  nor02 U3853 ( .Y(n5199), .A0(n7911), .A1(n7412) );
  nor02 U3854 ( .Y(n5200), .A0(n7910), .A1(n7417) );
  nor02 U3855 ( .Y(n5197), .A0(n5200), .A1(n5201) );
  nor02 U3856 ( .Y(n5202), .A0(n5198), .A1(n5199) );
  inv01 U3857 ( .Y(n5201), .A(n5202) );
  inv01 U3858 ( .Y(n2932), .A(n5203) );
  nor02 U3859 ( .Y(n5204), .A0(n7433), .A1(n2736) );
  nor02 U3860 ( .Y(n5205), .A0(n7826), .A1(n7411) );
  nor02 U3861 ( .Y(n5206), .A0(n7825), .A1(n7416) );
  nor02 U3862 ( .Y(n5203), .A0(n5206), .A1(n5207) );
  nor02 U3863 ( .Y(n5208), .A0(n5204), .A1(n5205) );
  inv01 U3864 ( .Y(n5207), .A(n5208) );
  inv01 U3865 ( .Y(n2936), .A(n5209) );
  nor02 U3866 ( .Y(n5210), .A0(n7433), .A1(n2783) );
  nor02 U3867 ( .Y(n5211), .A0(n7815), .A1(n7413) );
  nor02 U3868 ( .Y(n5212), .A0(n7814), .A1(n7415) );
  nor02 U3869 ( .Y(n5209), .A0(n5212), .A1(n5213) );
  nor02 U3870 ( .Y(n5214), .A0(n5210), .A1(n5211) );
  inv01 U3871 ( .Y(n5213), .A(n5214) );
  inv01 U3872 ( .Y(n2908), .A(n5215) );
  nor02 U3873 ( .Y(n5216), .A0(n7431), .A1(n2762) );
  nor02 U3874 ( .Y(n5217), .A0(n7887), .A1(n7411) );
  nor02 U3875 ( .Y(n5218), .A0(n7886), .A1(n7416) );
  nor02 U3876 ( .Y(n5215), .A0(n5218), .A1(n5219) );
  nor02 U3877 ( .Y(n5220), .A0(n5216), .A1(n5217) );
  inv01 U3878 ( .Y(n5219), .A(n5220) );
  inv01 U3879 ( .Y(n2873), .A(n5221) );
  nor02 U3880 ( .Y(n5222), .A0(n7607), .A1(n7431) );
  nor02 U3881 ( .Y(n5223), .A0(n7984), .A1(n7413) );
  nor02 U3882 ( .Y(n5224), .A0(n7983), .A1(n7415) );
  nor02 U3883 ( .Y(n5221), .A0(n5224), .A1(n5225) );
  nor02 U3884 ( .Y(n5226), .A0(n5222), .A1(n5223) );
  inv01 U3885 ( .Y(n5225), .A(n5226) );
  inv01 U3886 ( .Y(n2891), .A(n5227) );
  nor02 U3887 ( .Y(n5228), .A0(n7641), .A1(n7433) );
  nor02 U3888 ( .Y(n5229), .A0(n7930), .A1(n7413) );
  nor02 U3889 ( .Y(n5230), .A0(n7929), .A1(n7415) );
  nor02 U3890 ( .Y(n5227), .A0(n5230), .A1(n5231) );
  nor02 U3891 ( .Y(n5232), .A0(n5228), .A1(n5229) );
  inv01 U3892 ( .Y(n5231), .A(n5232) );
  inv01 U3893 ( .Y(n2926), .A(n5233) );
  nor02 U3894 ( .Y(n5234), .A0(n7432), .A1(n2742) );
  nor02 U3895 ( .Y(n5235), .A0(n7841), .A1(n7411) );
  nor02 U3896 ( .Y(n5236), .A0(n7840), .A1(n7416) );
  nor02 U3897 ( .Y(n5233), .A0(n5236), .A1(n5237) );
  nor02 U3898 ( .Y(n5238), .A0(n5234), .A1(n5235) );
  inv01 U3899 ( .Y(n5237), .A(n5238) );
  inv01 U3900 ( .Y(n2938), .A(n5239) );
  nor02 U3901 ( .Y(n5240), .A0(n7431), .A1(n2781) );
  nor02 U3902 ( .Y(n5241), .A0(n7811), .A1(n7411) );
  nor02 U3903 ( .Y(n5242), .A0(n7810), .A1(n7416) );
  nor02 U3904 ( .Y(n5239), .A0(n5242), .A1(n5243) );
  nor02 U3905 ( .Y(n5244), .A0(n5240), .A1(n5241) );
  inv01 U3906 ( .Y(n5243), .A(n5244) );
  inv01 U3907 ( .Y(n2870), .A(n5245) );
  nor02 U3908 ( .Y(n5246), .A0(n7591), .A1(n7433) );
  nor02 U3909 ( .Y(n5247), .A0(n7993), .A1(n7413) );
  nor02 U3910 ( .Y(n5248), .A0(n7992), .A1(n7415) );
  nor02 U3911 ( .Y(n5245), .A0(n5248), .A1(n5249) );
  nor02 U3912 ( .Y(n5250), .A0(n5246), .A1(n5247) );
  inv01 U3913 ( .Y(n5249), .A(n5250) );
  inv01 U3914 ( .Y(n2875), .A(n5251) );
  nor02 U3915 ( .Y(n5252), .A0(n7612), .A1(n7432) );
  nor02 U3916 ( .Y(n5253), .A0(n7978), .A1(n7411) );
  nor02 U3917 ( .Y(n5254), .A0(n7977), .A1(n7416) );
  nor02 U3918 ( .Y(n5251), .A0(n5254), .A1(n5255) );
  nor02 U3919 ( .Y(n5256), .A0(n5252), .A1(n5253) );
  inv01 U3920 ( .Y(n5255), .A(n5256) );
  inv01 U3921 ( .Y(n2934), .A(n5257) );
  nor02 U3922 ( .Y(n5258), .A0(n7433), .A1(n2734) );
  nor02 U3923 ( .Y(n5259), .A0(n7820), .A1(n7412) );
  nor02 U3924 ( .Y(n5260), .A0(n7819), .A1(n7417) );
  nor02 U3925 ( .Y(n5257), .A0(n5260), .A1(n5261) );
  nor02 U3926 ( .Y(n5262), .A0(n5258), .A1(n5259) );
  inv01 U3927 ( .Y(n5261), .A(n5262) );
  inv01 U3928 ( .Y(n2897), .A(n5263) );
  nor02 U3929 ( .Y(n5264), .A0(n7432), .A1(n2774) );
  nor02 U3930 ( .Y(n5265), .A0(n7914), .A1(n7413) );
  nor02 U3931 ( .Y(n5266), .A0(n7913), .A1(n7415) );
  nor02 U3932 ( .Y(n5263), .A0(n5266), .A1(n5267) );
  nor02 U3933 ( .Y(n5268), .A0(n5264), .A1(n5265) );
  inv01 U3934 ( .Y(n5267), .A(n5268) );
  inv01 U3935 ( .Y(n2943), .A(n5269) );
  nor02 U3936 ( .Y(n5270), .A0(n7432), .A1(n2754) );
  nor02 U3937 ( .Y(n5271), .A0(n7797), .A1(n7412) );
  nor02 U3938 ( .Y(n5272), .A0(n7796), .A1(n7417) );
  nor02 U3939 ( .Y(n5269), .A0(n5272), .A1(n5273) );
  nor02 U3940 ( .Y(n5274), .A0(n5270), .A1(n5271) );
  inv01 U3941 ( .Y(n5273), .A(n5274) );
  inv01 U3942 ( .Y(n2882), .A(n5275) );
  nor02 U3943 ( .Y(n5276), .A0(n7636), .A1(n7431) );
  nor02 U3944 ( .Y(n5277), .A0(n7957), .A1(n7413) );
  nor02 U3945 ( .Y(n5278), .A0(n7956), .A1(n7415) );
  nor02 U3946 ( .Y(n5275), .A0(n5278), .A1(n5279) );
  nor02 U3947 ( .Y(n5280), .A0(n5276), .A1(n5277) );
  inv01 U3948 ( .Y(n5279), .A(n5280) );
  inv01 U3949 ( .Y(n2925), .A(n5281) );
  nor02 U3950 ( .Y(n5282), .A0(n7432), .A1(n2744) );
  nor02 U3951 ( .Y(n5283), .A0(n7843), .A1(n7412) );
  nor02 U3952 ( .Y(n5284), .A0(n7842), .A1(n7417) );
  nor02 U3953 ( .Y(n5281), .A0(n5284), .A1(n5285) );
  nor02 U3954 ( .Y(n5286), .A0(n5282), .A1(n5283) );
  inv01 U3955 ( .Y(n5285), .A(n5286) );
  inv01 U3956 ( .Y(n2940), .A(n5287) );
  nor02 U3957 ( .Y(n5288), .A0(n7432), .A1(n2779) );
  nor02 U3958 ( .Y(n5289), .A0(n7805), .A1(n7412) );
  nor02 U3959 ( .Y(n5290), .A0(n7804), .A1(n7417) );
  nor02 U3960 ( .Y(n5287), .A0(n5290), .A1(n5291) );
  nor02 U3961 ( .Y(n5292), .A0(n5288), .A1(n5289) );
  inv01 U3962 ( .Y(n5291), .A(n5292) );
  inv01 U3963 ( .Y(n2911), .A(n5293) );
  nor02 U3964 ( .Y(n5294), .A0(n7432), .A1(n2759) );
  nor02 U3965 ( .Y(n5295), .A0(n7878), .A1(n7411) );
  nor02 U3966 ( .Y(n5296), .A0(n7877), .A1(n7416) );
  nor02 U3967 ( .Y(n5293), .A0(n5296), .A1(n5297) );
  nor02 U3968 ( .Y(n5298), .A0(n5294), .A1(n5295) );
  inv01 U3969 ( .Y(n5297), .A(n5298) );
  inv01 U3970 ( .Y(n2924), .A(n5299) );
  nor02 U3971 ( .Y(n5300), .A0(n7431), .A1(n2745) );
  nor02 U3972 ( .Y(n5301), .A0(n7845), .A1(n7413) );
  nor02 U3973 ( .Y(n5302), .A0(n7844), .A1(n7415) );
  nor02 U3974 ( .Y(n5299), .A0(n5302), .A1(n5303) );
  nor02 U3975 ( .Y(n5304), .A0(n5300), .A1(n5301) );
  inv01 U3976 ( .Y(n5303), .A(n5304) );
  inv01 U3977 ( .Y(n2896), .A(n5305) );
  nor02 U3978 ( .Y(n5306), .A0(n7431), .A1(n2775) );
  nor02 U3979 ( .Y(n5307), .A0(n7917), .A1(n7411) );
  nor02 U3980 ( .Y(n5308), .A0(n7916), .A1(n7416) );
  nor02 U3981 ( .Y(n5305), .A0(n5308), .A1(n5309) );
  nor02 U3982 ( .Y(n5310), .A0(n5306), .A1(n5307) );
  inv01 U3983 ( .Y(n5309), .A(n5310) );
  inv01 U3984 ( .Y(n2942), .A(n5311) );
  nor02 U3985 ( .Y(n5312), .A0(n7431), .A1(n2765) );
  nor02 U3986 ( .Y(n5313), .A0(n7800), .A1(n7413) );
  nor02 U3987 ( .Y(n5314), .A0(n7799), .A1(n7415) );
  nor02 U3988 ( .Y(n5311), .A0(n5314), .A1(n5315) );
  nor02 U3989 ( .Y(n5316), .A0(n5312), .A1(n5313) );
  inv01 U3990 ( .Y(n5315), .A(n5316) );
  inv01 U3991 ( .Y(n2890), .A(n5317) );
  nor02 U3992 ( .Y(n5318), .A0(n7642), .A1(n7432) );
  nor02 U3993 ( .Y(n5319), .A0(n7933), .A1(n7411) );
  nor02 U3994 ( .Y(n5320), .A0(n7932), .A1(n7416) );
  nor02 U3995 ( .Y(n5317), .A0(n5320), .A1(n5321) );
  nor02 U3996 ( .Y(n5322), .A0(n5318), .A1(n5319) );
  inv01 U3997 ( .Y(n5321), .A(n5322) );
  inv01 U3998 ( .Y(n2887), .A(n5323) );
  nor02 U3999 ( .Y(n5324), .A0(n7646), .A1(n7432) );
  nor02 U4000 ( .Y(n5325), .A0(n7942), .A1(n7411) );
  nor02 U4001 ( .Y(n5326), .A0(n7941), .A1(n7416) );
  nor02 U4002 ( .Y(n5323), .A0(n5326), .A1(n5327) );
  nor02 U4003 ( .Y(n5328), .A0(n5324), .A1(n5325) );
  inv01 U4004 ( .Y(n5327), .A(n5328) );
  inv01 U4005 ( .Y(n2933), .A(n5329) );
  nor02 U4006 ( .Y(n5330), .A0(n7431), .A1(n2735) );
  nor02 U4007 ( .Y(n5331), .A0(n7823), .A1(n7413) );
  nor02 U4008 ( .Y(n5332), .A0(n7822), .A1(n7415) );
  nor02 U4009 ( .Y(n5329), .A0(n5332), .A1(n5333) );
  nor02 U4010 ( .Y(n5334), .A0(n5330), .A1(n5331) );
  inv01 U4011 ( .Y(n5333), .A(n5334) );
  inv01 U4012 ( .Y(n2930), .A(n5335) );
  nor02 U4013 ( .Y(n5336), .A0(n7432), .A1(n2738) );
  nor02 U4014 ( .Y(n5337), .A0(n7830), .A1(n7413) );
  nor02 U4015 ( .Y(n5338), .A0(n7829), .A1(n7415) );
  nor02 U4016 ( .Y(n5335), .A0(n5338), .A1(n5339) );
  nor02 U4017 ( .Y(n5340), .A0(n5336), .A1(n5337) );
  inv01 U4018 ( .Y(n5339), .A(n5340) );
  inv01 U4019 ( .Y(n2901), .A(n5341) );
  nor02 U4020 ( .Y(n5342), .A0(n7431), .A1(n2770) );
  nor02 U4021 ( .Y(n5343), .A0(n7903), .A1(n7412) );
  nor02 U4022 ( .Y(n5344), .A0(n7902), .A1(n7417) );
  nor02 U4023 ( .Y(n5341), .A0(n5344), .A1(n5345) );
  nor02 U4024 ( .Y(n5346), .A0(n5342), .A1(n5343) );
  inv01 U4025 ( .Y(n5345), .A(n5346) );
  inv01 U4026 ( .Y(n2937), .A(n5347) );
  nor02 U4027 ( .Y(n5348), .A0(n7431), .A1(n2782) );
  nor02 U4028 ( .Y(n5349), .A0(n7813), .A1(n7412) );
  nor02 U4029 ( .Y(n5350), .A0(n7812), .A1(n7417) );
  nor02 U4030 ( .Y(n5347), .A0(n5350), .A1(n5351) );
  nor02 U4031 ( .Y(n5352), .A0(n5348), .A1(n5349) );
  inv01 U4032 ( .Y(n5351), .A(n5352) );
  inv01 U4033 ( .Y(n2905), .A(n5353) );
  nor02 U4034 ( .Y(n5354), .A0(n7433), .A1(n2766) );
  nor02 U4035 ( .Y(n5355), .A0(n7893), .A1(n7411) );
  nor02 U4036 ( .Y(n5356), .A0(n7892), .A1(n7416) );
  nor02 U4037 ( .Y(n5353), .A0(n5356), .A1(n5357) );
  nor02 U4038 ( .Y(n5358), .A0(n5354), .A1(n5355) );
  inv01 U4039 ( .Y(n5357), .A(n5358) );
  inv01 U4040 ( .Y(n2884), .A(n5359) );
  nor02 U4041 ( .Y(n5360), .A0(n7654), .A1(n7433) );
  nor02 U4042 ( .Y(n5361), .A0(n7951), .A1(n7411) );
  nor02 U4043 ( .Y(n5362), .A0(n7950), .A1(n7416) );
  nor02 U4044 ( .Y(n5359), .A0(n5362), .A1(n5363) );
  nor02 U4045 ( .Y(n5364), .A0(n5360), .A1(n5361) );
  inv01 U4046 ( .Y(n5363), .A(n5364) );
  inv01 U4047 ( .Y(n2874), .A(n5365) );
  nor02 U4048 ( .Y(n5366), .A0(n7613), .A1(n7432) );
  nor02 U4049 ( .Y(n5367), .A0(n7981), .A1(n7412) );
  nor02 U4050 ( .Y(n5368), .A0(n7980), .A1(n7417) );
  nor02 U4051 ( .Y(n5365), .A0(n5368), .A1(n5369) );
  nor02 U4052 ( .Y(n5370), .A0(n5366), .A1(n5367) );
  inv01 U4053 ( .Y(n5369), .A(n5370) );
  inv01 U4054 ( .Y(n2910), .A(n5371) );
  nor02 U4055 ( .Y(n5372), .A0(n7432), .A1(n2760) );
  nor02 U4056 ( .Y(n5373), .A0(n7881), .A1(n7412) );
  nor02 U4057 ( .Y(n5374), .A0(n7880), .A1(n7417) );
  nor02 U4058 ( .Y(n5371), .A0(n5374), .A1(n5375) );
  nor02 U4059 ( .Y(n5376), .A0(n5372), .A1(n5373) );
  inv01 U4060 ( .Y(n5375), .A(n5376) );
  inv01 U4061 ( .Y(n2904), .A(n5377) );
  nor02 U4062 ( .Y(n5378), .A0(n7431), .A1(n2767) );
  nor02 U4063 ( .Y(n5379), .A0(n7896), .A1(n7412) );
  nor02 U4064 ( .Y(n5380), .A0(n7895), .A1(n7417) );
  nor02 U4065 ( .Y(n5377), .A0(n5380), .A1(n5381) );
  nor02 U4066 ( .Y(n5382), .A0(n5378), .A1(n5379) );
  inv01 U4067 ( .Y(n5381), .A(n5382) );
  inv01 U4068 ( .Y(n2918), .A(n5383) );
  nor02 U4069 ( .Y(n5384), .A0(n7432), .A1(n2751) );
  nor02 U4070 ( .Y(n5385), .A0(n7861), .A1(n7413) );
  nor02 U4071 ( .Y(n5386), .A0(n7860), .A1(n7415) );
  nor02 U4072 ( .Y(n5383), .A0(n5386), .A1(n5387) );
  nor02 U4073 ( .Y(n5388), .A0(n5384), .A1(n5385) );
  inv01 U4074 ( .Y(n5387), .A(n5388) );
  inv01 U4075 ( .Y(n2892), .A(n5389) );
  nor02 U4076 ( .Y(n5390), .A0(n7652), .A1(n7431) );
  nor02 U4077 ( .Y(n5391), .A0(n7927), .A1(n7412) );
  nor02 U4078 ( .Y(n5392), .A0(n7926), .A1(n7417) );
  nor02 U4079 ( .Y(n5389), .A0(n5392), .A1(n5393) );
  nor02 U4080 ( .Y(n5394), .A0(n5390), .A1(n5391) );
  inv01 U4081 ( .Y(n5393), .A(n5394) );
  inv01 U4082 ( .Y(n2885), .A(n5395) );
  nor02 U4083 ( .Y(n5396), .A0(n7656), .A1(n7433) );
  nor02 U4084 ( .Y(n5397), .A0(n7948), .A1(n7413) );
  nor02 U4085 ( .Y(n5398), .A0(n7947), .A1(n7415) );
  nor02 U4086 ( .Y(n5395), .A0(n5398), .A1(n5399) );
  nor02 U4087 ( .Y(n5400), .A0(n5396), .A1(n5397) );
  inv01 U4088 ( .Y(n5399), .A(n5400) );
  inv01 U4089 ( .Y(n2880), .A(n5401) );
  nor02 U4090 ( .Y(n5402), .A0(n7629), .A1(n7432) );
  nor02 U4091 ( .Y(n5403), .A0(n7963), .A1(n7412) );
  nor02 U4092 ( .Y(n5404), .A0(n7962), .A1(n7417) );
  nor02 U4093 ( .Y(n5401), .A0(n5404), .A1(n5405) );
  nor02 U4094 ( .Y(n5406), .A0(n5402), .A1(n5403) );
  inv01 U4095 ( .Y(n5405), .A(n5406) );
  inv01 U4096 ( .Y(n2944), .A(n5407) );
  nor02 U4097 ( .Y(n5408), .A0(n7432), .A1(n2743) );
  nor02 U4098 ( .Y(n5409), .A0(n7795), .A1(n7411) );
  nor02 U4099 ( .Y(n5410), .A0(n7794), .A1(n7416) );
  nor02 U4100 ( .Y(n5407), .A0(n5410), .A1(n5411) );
  nor02 U4101 ( .Y(n5412), .A0(n5408), .A1(n5409) );
  inv01 U4102 ( .Y(n5411), .A(n5412) );
  inv01 U4103 ( .Y(n2893), .A(n5413) );
  nor02 U4104 ( .Y(n5414), .A0(n7658), .A1(n7433) );
  nor02 U4105 ( .Y(n5415), .A0(n7924), .A1(n7411) );
  nor02 U4106 ( .Y(n5416), .A0(n7923), .A1(n7416) );
  nor02 U4107 ( .Y(n5413), .A0(n5416), .A1(n5417) );
  nor02 U4108 ( .Y(n5418), .A0(n5414), .A1(n5415) );
  inv01 U4109 ( .Y(n5417), .A(n5418) );
  inv01 U4110 ( .Y(n2945), .A(n5419) );
  nor02 U4111 ( .Y(n5420), .A0(n7432), .A1(n2732) );
  nor02 U4112 ( .Y(n5421), .A0(n7792), .A1(n7413) );
  nor02 U4113 ( .Y(n5422), .A0(n7790), .A1(n7415) );
  nor02 U4114 ( .Y(n5419), .A0(n5422), .A1(n5423) );
  nor02 U4115 ( .Y(n5424), .A0(n5420), .A1(n5421) );
  inv01 U4116 ( .Y(n5423), .A(n5424) );
  inv01 U4117 ( .Y(n7462), .A(n5425) );
  nor02 U4118 ( .Y(n5426), .A0(n7395), .A1(n7465) );
  nor02 U4119 ( .Y(n5427), .A0(n7403), .A1(n7464) );
  inv01 U4120 ( .Y(n5428), .A(n7466) );
  nor02 U4121 ( .Y(n5425), .A0(n5428), .A1(n5429) );
  nor02 U4122 ( .Y(n5430), .A0(n5426), .A1(n5427) );
  inv01 U4123 ( .Y(n5429), .A(n5430) );
  inv01 U4124 ( .Y(n7449), .A(n5431) );
  nor02 U4125 ( .Y(n5432), .A0(n7393), .A1(n7455) );
  nor02 U4126 ( .Y(n5433), .A0(n7403), .A1(n7453) );
  inv01 U4127 ( .Y(n5434), .A(n7456) );
  nor02 U4128 ( .Y(n5431), .A0(n5434), .A1(n5435) );
  nor02 U4129 ( .Y(n5436), .A0(n5432), .A1(n5433) );
  inv01 U4130 ( .Y(n5435), .A(n5436) );
  inv01 U4131 ( .Y(n7472), .A(n5437) );
  nor02 U4132 ( .Y(n5438), .A0(n7394), .A1(n7464) );
  nor02 U4133 ( .Y(n5439), .A0(n7403), .A1(n7474) );
  inv01 U4134 ( .Y(n5440), .A(n7475) );
  nor02 U4135 ( .Y(n5437), .A0(n5440), .A1(n5441) );
  nor02 U4136 ( .Y(n5442), .A0(n5438), .A1(n5439) );
  inv01 U4137 ( .Y(n5441), .A(n5442) );
  buf04 U4138 ( .Y(n7395), .A(n7392) );
  buf04 U4139 ( .Y(n7394), .A(n7391) );
  inv01 U4140 ( .Y(n7667), .A(n5443) );
  nor02 U4141 ( .Y(n5444), .A0(n7394), .A1(n7453) );
  nor02 U4142 ( .Y(n5445), .A0(n7404), .A1(n7465) );
  inv01 U4143 ( .Y(n5446), .A(n3838) );
  nor02 U4144 ( .Y(n5443), .A0(n5446), .A1(n5447) );
  nor02 U4145 ( .Y(n5448), .A0(n5444), .A1(n5445) );
  inv01 U4146 ( .Y(n5447), .A(n5448) );
  inv01 U4147 ( .Y(n7441), .A(n5449) );
  nor02 U4148 ( .Y(n5450), .A0(n7663), .A1(n5451) );
  nor02 U4149 ( .Y(n5452), .A0(n7663), .A1(n5453) );
  nor02 U4150 ( .Y(n5454), .A0(n7663), .A1(n5455) );
  nor02 U4151 ( .Y(n5456), .A0(n7663), .A1(n5457) );
  nor02 U4152 ( .Y(n5458), .A0(r0_0_), .A1(n5459) );
  nor02 U4153 ( .Y(n5460), .A0(r0_0_), .A1(n5461) );
  nor02 U4154 ( .Y(n5462), .A0(r0_0_), .A1(n5463) );
  nor02 U4155 ( .Y(n5464), .A0(r0_0_), .A1(n5465) );
  nor02 U4156 ( .Y(n5449), .A0(n5466), .A1(n5467) );
  nor02 U4157 ( .Y(n5468), .A0(r0_2_), .A1(r0_1_) );
  inv01 U4158 ( .Y(n5451), .A(n5468) );
  nor02 U4159 ( .Y(n5469), .A0(n7400), .A1(r0_1_) );
  inv01 U4160 ( .Y(n5453), .A(n5469) );
  nor02 U4161 ( .Y(n5470), .A0(r0_2_), .A1(n7401) );
  inv01 U4162 ( .Y(n5455), .A(n5470) );
  nor02 U4163 ( .Y(n5471), .A0(n7400), .A1(n7401) );
  inv01 U4164 ( .Y(n5457), .A(n5471) );
  nor02 U4165 ( .Y(n5472), .A0(r0_2_), .A1(r0_1_) );
  inv01 U4166 ( .Y(n5459), .A(n5472) );
  nor02 U4167 ( .Y(n5473), .A0(n7400), .A1(r0_1_) );
  inv01 U4168 ( .Y(n5461), .A(n5473) );
  nor02 U4169 ( .Y(n5474), .A0(r0_2_), .A1(n7401) );
  inv01 U4170 ( .Y(n5463), .A(n5474) );
  nor02 U4171 ( .Y(n5475), .A0(n7400), .A1(n7401) );
  inv01 U4172 ( .Y(n5465), .A(n5475) );
  nor02 U4173 ( .Y(n5476), .A0(n5450), .A1(n5452) );
  inv01 U4174 ( .Y(n5477), .A(n5476) );
  nor02 U4175 ( .Y(n5478), .A0(n5454), .A1(n5456) );
  inv01 U4176 ( .Y(n5479), .A(n5478) );
  nor02 U4177 ( .Y(n5480), .A0(n5477), .A1(n5479) );
  inv01 U4178 ( .Y(n5466), .A(n5480) );
  nor02 U4179 ( .Y(n5481), .A0(n5458), .A1(n5460) );
  inv01 U4180 ( .Y(n5482), .A(n5481) );
  nor02 U4181 ( .Y(n5483), .A0(n5462), .A1(n5464) );
  inv01 U4182 ( .Y(n5484), .A(n5483) );
  nor02 U4183 ( .Y(n5485), .A0(n5482), .A1(n5484) );
  inv01 U4184 ( .Y(n5467), .A(n5485) );
  inv02 U4185 ( .Y(n7663), .A(n7454) );
  buf04 U4186 ( .Y(n5486), .A(n7484) );
  inv01 U4187 ( .Y(n7484), .A(n7446) );
  nand02 U4188 ( .Y(n7540), .A0(n5487), .A1(n5488) );
  inv02 U4189 ( .Y(n5489), .A(n7500) );
  inv02 U4190 ( .Y(n5490), .A(n7476) );
  inv02 U4191 ( .Y(n5491), .A(n7521) );
  inv02 U4192 ( .Y(n5492), .A(n7368) );
  inv02 U4193 ( .Y(n5493), .A(n7369) );
  inv02 U4194 ( .Y(n5494), .A(n7370) );
  nand02 U4195 ( .Y(n5495), .A0(n5491), .A1(n5496) );
  nand02 U4196 ( .Y(n5497), .A0(n5492), .A1(n5498) );
  nand02 U4197 ( .Y(n5499), .A0(n5493), .A1(n5500) );
  nand02 U4198 ( .Y(n5501), .A0(n5493), .A1(n5502) );
  nand02 U4199 ( .Y(n5503), .A0(n5494), .A1(n5504) );
  nand02 U4200 ( .Y(n5505), .A0(n5494), .A1(n5506) );
  nand02 U4201 ( .Y(n5507), .A0(n5494), .A1(n5508) );
  nand02 U4202 ( .Y(n5509), .A0(n5494), .A1(n5510) );
  nand02 U4203 ( .Y(n5511), .A0(n5489), .A1(n5490) );
  inv01 U4204 ( .Y(n5496), .A(n5511) );
  nand02 U4205 ( .Y(n5512), .A0(n5489), .A1(n5490) );
  inv01 U4206 ( .Y(n5498), .A(n5512) );
  nand02 U4207 ( .Y(n5513), .A0(n5489), .A1(n5491) );
  inv01 U4208 ( .Y(n5500), .A(n5513) );
  nand02 U4209 ( .Y(n5514), .A0(n5489), .A1(n5492) );
  inv01 U4210 ( .Y(n5502), .A(n5514) );
  nand02 U4211 ( .Y(n5515), .A0(n5490), .A1(n5491) );
  inv01 U4212 ( .Y(n5504), .A(n5515) );
  nand02 U4213 ( .Y(n5516), .A0(n5490), .A1(n5492) );
  inv01 U4214 ( .Y(n5506), .A(n5516) );
  nand02 U4215 ( .Y(n5517), .A0(n5491), .A1(n5493) );
  inv01 U4216 ( .Y(n5508), .A(n5517) );
  nand02 U4217 ( .Y(n5518), .A0(n5492), .A1(n5493) );
  inv01 U4218 ( .Y(n5510), .A(n5518) );
  nand02 U4219 ( .Y(n5519), .A0(n5495), .A1(n5497) );
  inv01 U4220 ( .Y(n5520), .A(n5519) );
  nand02 U4221 ( .Y(n5521), .A0(n5499), .A1(n5501) );
  inv01 U4222 ( .Y(n5522), .A(n5521) );
  nand02 U4223 ( .Y(n5523), .A0(n5520), .A1(n5522) );
  inv01 U4224 ( .Y(n5487), .A(n5523) );
  nand02 U4225 ( .Y(n5524), .A0(n5503), .A1(n5505) );
  inv01 U4226 ( .Y(n5525), .A(n5524) );
  nand02 U4227 ( .Y(n5526), .A0(n5507), .A1(n5509) );
  inv01 U4228 ( .Y(n5527), .A(n5526) );
  nand02 U4229 ( .Y(n5528), .A0(n5525), .A1(n5527) );
  inv01 U4230 ( .Y(n5488), .A(n5528) );
  nand02 U4231 ( .Y(n7533), .A0(n5529), .A1(n5530) );
  inv02 U4232 ( .Y(n5531), .A(n7494) );
  inv02 U4233 ( .Y(n5532), .A(n7516) );
  inv02 U4234 ( .Y(n5533), .A(n7368) );
  inv02 U4235 ( .Y(n5534), .A(n7369) );
  inv02 U4236 ( .Y(n5535), .A(n7370) );
  nand02 U4237 ( .Y(n5536), .A0(n5532), .A1(n5537) );
  nand02 U4238 ( .Y(n5538), .A0(n5533), .A1(n5539) );
  nand02 U4239 ( .Y(n5540), .A0(n5534), .A1(n5541) );
  nand02 U4240 ( .Y(n5542), .A0(n5534), .A1(n5543) );
  nand02 U4241 ( .Y(n5544), .A0(n5535), .A1(n5545) );
  nand02 U4242 ( .Y(n5546), .A0(n5535), .A1(n5547) );
  nand02 U4243 ( .Y(n5548), .A0(n5535), .A1(n5549) );
  nand02 U4244 ( .Y(n5550), .A0(n5535), .A1(n5551) );
  nand02 U4245 ( .Y(n5552), .A0(n5531), .A1(n7459) );
  inv01 U4246 ( .Y(n5537), .A(n5552) );
  nand02 U4247 ( .Y(n5553), .A0(n5531), .A1(n5658) );
  inv01 U4248 ( .Y(n5539), .A(n5553) );
  nand02 U4249 ( .Y(n5554), .A0(n5531), .A1(n5532) );
  inv01 U4250 ( .Y(n5541), .A(n5554) );
  nand02 U4251 ( .Y(n5555), .A0(n5531), .A1(n5533) );
  inv01 U4252 ( .Y(n5543), .A(n5555) );
  nand02 U4253 ( .Y(n5556), .A0(n5658), .A1(n5532) );
  inv01 U4254 ( .Y(n5545), .A(n5556) );
  nand02 U4255 ( .Y(n5557), .A0(n5658), .A1(n5533) );
  inv01 U4256 ( .Y(n5547), .A(n5557) );
  nand02 U4257 ( .Y(n5558), .A0(n5532), .A1(n5534) );
  inv01 U4258 ( .Y(n5549), .A(n5558) );
  nand02 U4259 ( .Y(n5559), .A0(n5533), .A1(n5534) );
  inv01 U4260 ( .Y(n5551), .A(n5559) );
  nand02 U4261 ( .Y(n5560), .A0(n5536), .A1(n5538) );
  inv01 U4262 ( .Y(n5561), .A(n5560) );
  nand02 U4263 ( .Y(n5562), .A0(n5540), .A1(n5542) );
  inv01 U4264 ( .Y(n5563), .A(n5562) );
  nand02 U4265 ( .Y(n5564), .A0(n5561), .A1(n5563) );
  inv01 U4266 ( .Y(n5529), .A(n5564) );
  nand02 U4267 ( .Y(n5565), .A0(n5544), .A1(n5546) );
  inv01 U4268 ( .Y(n5566), .A(n5565) );
  nand02 U4269 ( .Y(n5567), .A0(n5548), .A1(n5550) );
  inv01 U4270 ( .Y(n5568), .A(n5567) );
  nand02 U4271 ( .Y(n5569), .A0(n5566), .A1(n5568) );
  inv01 U4272 ( .Y(n5530), .A(n5569) );
  nand02 U4273 ( .Y(n7523), .A0(n5570), .A1(n5571) );
  inv02 U4274 ( .Y(n5572), .A(n7481) );
  inv02 U4275 ( .Y(n5573), .A(n7458) );
  inv02 U4276 ( .Y(n5574), .A(n7506) );
  inv02 U4277 ( .Y(n5575), .A(n7368) );
  inv02 U4278 ( .Y(n5576), .A(n7369) );
  inv02 U4279 ( .Y(n5577), .A(n7370) );
  nand02 U4280 ( .Y(n5578), .A0(n5574), .A1(n5579) );
  nand02 U4281 ( .Y(n5580), .A0(n5575), .A1(n5581) );
  nand02 U4282 ( .Y(n5582), .A0(n5576), .A1(n5583) );
  nand02 U4283 ( .Y(n5584), .A0(n5576), .A1(n5585) );
  nand02 U4284 ( .Y(n5586), .A0(n5577), .A1(n5587) );
  nand02 U4285 ( .Y(n5588), .A0(n5577), .A1(n5589) );
  nand02 U4286 ( .Y(n5590), .A0(n5577), .A1(n5591) );
  nand02 U4287 ( .Y(n5592), .A0(n5577), .A1(n5593) );
  nand02 U4288 ( .Y(n5594), .A0(n5572), .A1(n5573) );
  inv01 U4289 ( .Y(n5579), .A(n5594) );
  nand02 U4290 ( .Y(n5595), .A0(n5572), .A1(n5573) );
  inv01 U4291 ( .Y(n5581), .A(n5595) );
  nand02 U4292 ( .Y(n5596), .A0(n5572), .A1(n5574) );
  inv01 U4293 ( .Y(n5583), .A(n5596) );
  nand02 U4294 ( .Y(n5597), .A0(n5572), .A1(n5575) );
  inv01 U4295 ( .Y(n5585), .A(n5597) );
  nand02 U4296 ( .Y(n5598), .A0(n5573), .A1(n5574) );
  inv01 U4297 ( .Y(n5587), .A(n5598) );
  nand02 U4298 ( .Y(n5599), .A0(n5573), .A1(n5575) );
  inv01 U4299 ( .Y(n5589), .A(n5599) );
  nand02 U4300 ( .Y(n5600), .A0(n5574), .A1(n5576) );
  inv01 U4301 ( .Y(n5591), .A(n5600) );
  nand02 U4302 ( .Y(n5601), .A0(n5575), .A1(n5576) );
  inv01 U4303 ( .Y(n5593), .A(n5601) );
  nand02 U4304 ( .Y(n5602), .A0(n5578), .A1(n5580) );
  inv01 U4305 ( .Y(n5603), .A(n5602) );
  nand02 U4306 ( .Y(n5604), .A0(n5582), .A1(n5584) );
  inv01 U4307 ( .Y(n5605), .A(n5604) );
  nand02 U4308 ( .Y(n5606), .A0(n5603), .A1(n5605) );
  inv01 U4309 ( .Y(n5570), .A(n5606) );
  nand02 U4310 ( .Y(n5607), .A0(n5586), .A1(n5588) );
  inv01 U4311 ( .Y(n5608), .A(n5607) );
  nand02 U4312 ( .Y(n5609), .A0(n5590), .A1(n5592) );
  inv01 U4313 ( .Y(n5610), .A(n5609) );
  nand02 U4314 ( .Y(n5611), .A0(n5608), .A1(n5610) );
  inv01 U4315 ( .Y(n5571), .A(n5611) );
  nand02 U4316 ( .Y(n7470), .A0(n5612), .A1(n5613) );
  inv02 U4317 ( .Y(n5614), .A(n7473) );
  inv02 U4318 ( .Y(n5615), .A(n7472) );
  inv02 U4319 ( .Y(n5616), .A(n7471) );
  inv02 U4320 ( .Y(n5617), .A(n7368) );
  inv02 U4321 ( .Y(n5618), .A(n7369) );
  inv02 U4322 ( .Y(n5619), .A(n7370) );
  nand02 U4323 ( .Y(n5620), .A0(n5616), .A1(n5621) );
  nand02 U4324 ( .Y(n5622), .A0(n5617), .A1(n5623) );
  nand02 U4325 ( .Y(n5624), .A0(n5618), .A1(n5625) );
  nand02 U4326 ( .Y(n5626), .A0(n5618), .A1(n5627) );
  nand02 U4327 ( .Y(n5628), .A0(n5619), .A1(n5629) );
  nand02 U4328 ( .Y(n5630), .A0(n5619), .A1(n5631) );
  nand02 U4329 ( .Y(n5632), .A0(n5619), .A1(n5633) );
  nand02 U4330 ( .Y(n5634), .A0(n5619), .A1(n5635) );
  nand02 U4331 ( .Y(n5636), .A0(n5614), .A1(n5615) );
  inv01 U4332 ( .Y(n5621), .A(n5636) );
  nand02 U4333 ( .Y(n5637), .A0(n5614), .A1(n5615) );
  inv01 U4334 ( .Y(n5623), .A(n5637) );
  nand02 U4335 ( .Y(n5638), .A0(n5614), .A1(n5616) );
  inv01 U4336 ( .Y(n5625), .A(n5638) );
  nand02 U4337 ( .Y(n5639), .A0(n5614), .A1(n5617) );
  inv01 U4338 ( .Y(n5627), .A(n5639) );
  nand02 U4339 ( .Y(n5640), .A0(n5615), .A1(n5616) );
  inv01 U4340 ( .Y(n5629), .A(n5640) );
  nand02 U4341 ( .Y(n5641), .A0(n5615), .A1(n5617) );
  inv01 U4342 ( .Y(n5631), .A(n5641) );
  nand02 U4343 ( .Y(n5642), .A0(n5616), .A1(n5618) );
  inv01 U4344 ( .Y(n5633), .A(n5642) );
  nand02 U4345 ( .Y(n5643), .A0(n5617), .A1(n5618) );
  inv01 U4346 ( .Y(n5635), .A(n5643) );
  nand02 U4347 ( .Y(n5644), .A0(n5620), .A1(n5622) );
  inv01 U4348 ( .Y(n5645), .A(n5644) );
  nand02 U4349 ( .Y(n5646), .A0(n5624), .A1(n5626) );
  inv01 U4350 ( .Y(n5647), .A(n5646) );
  nand02 U4351 ( .Y(n5648), .A0(n5645), .A1(n5647) );
  inv01 U4352 ( .Y(n5612), .A(n5648) );
  nand02 U4353 ( .Y(n5649), .A0(n5628), .A1(n5630) );
  inv01 U4354 ( .Y(n5650), .A(n5649) );
  nand02 U4355 ( .Y(n5651), .A0(n5632), .A1(n5634) );
  inv01 U4356 ( .Y(n5652), .A(n5651) );
  nand02 U4357 ( .Y(n5653), .A0(n5650), .A1(n5652) );
  inv01 U4358 ( .Y(n5613), .A(n5653) );
  inv02 U4359 ( .Y(n7473), .A(n6589) );
  nand02 U4360 ( .Y(n7491), .A0(n5654), .A1(n5655) );
  inv02 U4361 ( .Y(n5656), .A(n7461) );
  inv02 U4362 ( .Y(n5657), .A(n7463) );
  inv02 U4363 ( .Y(n5658), .A(n7467) );
  inv02 U4364 ( .Y(n5659), .A(n7368) );
  inv02 U4365 ( .Y(n5660), .A(n7369) );
  inv02 U4366 ( .Y(n5661), .A(n7370) );
  nand02 U4367 ( .Y(n5662), .A0(n5658), .A1(n5663) );
  nand02 U4368 ( .Y(n5664), .A0(n5659), .A1(n5665) );
  nand02 U4369 ( .Y(n5666), .A0(n5660), .A1(n5667) );
  nand02 U4370 ( .Y(n5668), .A0(n5660), .A1(n5669) );
  nand02 U4371 ( .Y(n5670), .A0(n5661), .A1(n5671) );
  nand02 U4372 ( .Y(n5672), .A0(n5661), .A1(n5673) );
  nand02 U4373 ( .Y(n5674), .A0(n5661), .A1(n5675) );
  nand02 U4374 ( .Y(n5676), .A0(n5661), .A1(n5677) );
  nand02 U4375 ( .Y(n5678), .A0(n5656), .A1(n5657) );
  inv01 U4376 ( .Y(n5663), .A(n5678) );
  nand02 U4377 ( .Y(n5679), .A0(n5656), .A1(n5657) );
  inv01 U4378 ( .Y(n5665), .A(n5679) );
  nand02 U4379 ( .Y(n5680), .A0(n5656), .A1(n5658) );
  inv01 U4380 ( .Y(n5667), .A(n5680) );
  nand02 U4381 ( .Y(n5681), .A0(n5656), .A1(n5659) );
  inv01 U4382 ( .Y(n5669), .A(n5681) );
  nand02 U4383 ( .Y(n5682), .A0(n5657), .A1(n5658) );
  inv01 U4384 ( .Y(n5671), .A(n5682) );
  nand02 U4385 ( .Y(n5683), .A0(n5657), .A1(n5659) );
  inv01 U4386 ( .Y(n5673), .A(n5683) );
  nand02 U4387 ( .Y(n5684), .A0(n5658), .A1(n5660) );
  inv01 U4388 ( .Y(n5675), .A(n5684) );
  nand02 U4389 ( .Y(n5685), .A0(n5659), .A1(n5660) );
  inv01 U4390 ( .Y(n5677), .A(n5685) );
  nand02 U4391 ( .Y(n5686), .A0(n5662), .A1(n5664) );
  inv01 U4392 ( .Y(n5687), .A(n5686) );
  nand02 U4393 ( .Y(n5688), .A0(n5666), .A1(n5668) );
  inv01 U4394 ( .Y(n5689), .A(n5688) );
  nand02 U4395 ( .Y(n5690), .A0(n5687), .A1(n5689) );
  inv01 U4396 ( .Y(n5654), .A(n5690) );
  nand02 U4397 ( .Y(n5691), .A0(n5670), .A1(n5672) );
  inv01 U4398 ( .Y(n5692), .A(n5691) );
  nand02 U4399 ( .Y(n5693), .A0(n5674), .A1(n5676) );
  inv01 U4400 ( .Y(n5694), .A(n5693) );
  nand02 U4401 ( .Y(n5695), .A0(n5692), .A1(n5694) );
  inv01 U4402 ( .Y(n5655), .A(n5695) );
  inv02 U4403 ( .Y(n7463), .A(n6601) );
  nand02 U4404 ( .Y(n7666), .A0(n5696), .A1(n5697) );
  inv02 U4405 ( .Y(n5698), .A(n7488) );
  inv02 U4406 ( .Y(n5699), .A(n7667) );
  inv02 U4407 ( .Y(n5700), .A(n7510) );
  inv02 U4408 ( .Y(n5701), .A(n7527) );
  inv02 U4409 ( .Y(n5702), .A(n7369) );
  inv02 U4410 ( .Y(n5703), .A(n7370) );
  nand02 U4411 ( .Y(n5704), .A0(n5700), .A1(n5705) );
  nand02 U4412 ( .Y(n5706), .A0(n5701), .A1(n5707) );
  nand02 U4413 ( .Y(n5708), .A0(n5702), .A1(n5709) );
  nand02 U4414 ( .Y(n5710), .A0(n5702), .A1(n5711) );
  nand02 U4415 ( .Y(n5712), .A0(n5703), .A1(n5713) );
  nand02 U4416 ( .Y(n5714), .A0(n5703), .A1(n5715) );
  nand02 U4417 ( .Y(n5716), .A0(n5703), .A1(n5717) );
  nand02 U4418 ( .Y(n5718), .A0(n5703), .A1(n5719) );
  nand02 U4419 ( .Y(n5720), .A0(n5698), .A1(n5699) );
  inv01 U4420 ( .Y(n5705), .A(n5720) );
  nand02 U4421 ( .Y(n5721), .A0(n5698), .A1(n5699) );
  inv01 U4422 ( .Y(n5707), .A(n5721) );
  nand02 U4423 ( .Y(n5722), .A0(n5698), .A1(n5700) );
  inv01 U4424 ( .Y(n5709), .A(n5722) );
  nand02 U4425 ( .Y(n5723), .A0(n5698), .A1(n5701) );
  inv01 U4426 ( .Y(n5711), .A(n5723) );
  nand02 U4427 ( .Y(n5724), .A0(n5699), .A1(n5700) );
  inv01 U4428 ( .Y(n5713), .A(n5724) );
  nand02 U4429 ( .Y(n5725), .A0(n5699), .A1(n5701) );
  inv01 U4430 ( .Y(n5715), .A(n5725) );
  nand02 U4431 ( .Y(n5726), .A0(n5700), .A1(n5702) );
  inv01 U4432 ( .Y(n5717), .A(n5726) );
  nand02 U4433 ( .Y(n5727), .A0(n5701), .A1(n5702) );
  inv01 U4434 ( .Y(n5719), .A(n5727) );
  nand02 U4435 ( .Y(n5728), .A0(n5704), .A1(n5706) );
  inv01 U4436 ( .Y(n5729), .A(n5728) );
  nand02 U4437 ( .Y(n5730), .A0(n5708), .A1(n5710) );
  inv01 U4438 ( .Y(n5731), .A(n5730) );
  nand02 U4439 ( .Y(n5732), .A0(n5729), .A1(n5731) );
  inv01 U4440 ( .Y(n5696), .A(n5732) );
  nand02 U4441 ( .Y(n5733), .A0(n5712), .A1(n5714) );
  inv01 U4442 ( .Y(n5734), .A(n5733) );
  nand02 U4443 ( .Y(n5735), .A0(n5716), .A1(n5718) );
  inv01 U4444 ( .Y(n5736), .A(n5735) );
  nand02 U4445 ( .Y(n5737), .A0(n5734), .A1(n5736) );
  inv01 U4446 ( .Y(n5697), .A(n5737) );
  nand02 U4447 ( .Y(n7508), .A0(n5738), .A1(n5739) );
  inv02 U4448 ( .Y(n5740), .A(n7510) );
  inv02 U4449 ( .Y(n5741), .A(n7509) );
  inv02 U4450 ( .Y(n5742), .A(n7486) );
  inv02 U4451 ( .Y(n5743), .A(n7369) );
  inv02 U4452 ( .Y(n5744), .A(n7380) );
  inv02 U4453 ( .Y(n5745), .A(n7370) );
  nand02 U4454 ( .Y(n5746), .A0(n5742), .A1(n5747) );
  nand02 U4455 ( .Y(n5748), .A0(n5743), .A1(n5749) );
  nand02 U4456 ( .Y(n5750), .A0(n5744), .A1(n5751) );
  nand02 U4457 ( .Y(n5752), .A0(n5744), .A1(n5753) );
  nand02 U4458 ( .Y(n5754), .A0(n5745), .A1(n5755) );
  nand02 U4459 ( .Y(n5756), .A0(n5745), .A1(n5757) );
  nand02 U4460 ( .Y(n5758), .A0(n5745), .A1(n5759) );
  nand02 U4461 ( .Y(n5760), .A0(n5745), .A1(n5761) );
  nand02 U4462 ( .Y(n5762), .A0(n5740), .A1(n5741) );
  inv01 U4463 ( .Y(n5747), .A(n5762) );
  nand02 U4464 ( .Y(n5763), .A0(n5740), .A1(n5741) );
  inv01 U4465 ( .Y(n5749), .A(n5763) );
  nand02 U4466 ( .Y(n5764), .A0(n5740), .A1(n5742) );
  inv01 U4467 ( .Y(n5751), .A(n5764) );
  nand02 U4468 ( .Y(n5765), .A0(n5740), .A1(n5743) );
  inv01 U4469 ( .Y(n5753), .A(n5765) );
  nand02 U4470 ( .Y(n5766), .A0(n5741), .A1(n5742) );
  inv01 U4471 ( .Y(n5755), .A(n5766) );
  nand02 U4472 ( .Y(n5767), .A0(n5741), .A1(n5743) );
  inv01 U4473 ( .Y(n5757), .A(n5767) );
  nand02 U4474 ( .Y(n5768), .A0(n5742), .A1(n5744) );
  inv01 U4475 ( .Y(n5759), .A(n5768) );
  nand02 U4476 ( .Y(n5769), .A0(n5743), .A1(n5744) );
  inv01 U4477 ( .Y(n5761), .A(n5769) );
  nand02 U4478 ( .Y(n5770), .A0(n5746), .A1(n5748) );
  inv01 U4479 ( .Y(n5771), .A(n5770) );
  nand02 U4480 ( .Y(n5772), .A0(n5750), .A1(n5752) );
  inv01 U4481 ( .Y(n5773), .A(n5772) );
  nand02 U4482 ( .Y(n5774), .A0(n5771), .A1(n5773) );
  inv01 U4483 ( .Y(n5738), .A(n5774) );
  nand02 U4484 ( .Y(n5775), .A0(n5754), .A1(n5756) );
  inv01 U4485 ( .Y(n5776), .A(n5775) );
  nand02 U4486 ( .Y(n5777), .A0(n5758), .A1(n5760) );
  inv01 U4487 ( .Y(n5778), .A(n5777) );
  nand02 U4488 ( .Y(n5779), .A0(n5776), .A1(n5778) );
  inv01 U4489 ( .Y(n5739), .A(n5779) );
  inv01 U4490 ( .Y(n7485), .A(n5780) );
  nor02 U4491 ( .Y(n5781), .A0(n7488), .A1(n5782) );
  nor02 U4492 ( .Y(n5783), .A0(n7488), .A1(n5784) );
  nor02 U4493 ( .Y(n5785), .A0(n7488), .A1(n5786) );
  nor02 U4494 ( .Y(n5787), .A0(n7488), .A1(n5788) );
  nor02 U4495 ( .Y(n5789), .A0(n7369), .A1(n5790) );
  nor02 U4496 ( .Y(n5791), .A0(n7369), .A1(n5792) );
  nor02 U4497 ( .Y(n5793), .A0(n7369), .A1(n5794) );
  nor02 U4498 ( .Y(n5795), .A0(n7369), .A1(n5796) );
  nor02 U4499 ( .Y(n5780), .A0(n5797), .A1(n5798) );
  nor02 U4500 ( .Y(n5799), .A0(n7486), .A1(n7487) );
  inv01 U4501 ( .Y(n5782), .A(n5799) );
  nor02 U4502 ( .Y(n5800), .A0(n7370), .A1(n7487) );
  inv01 U4503 ( .Y(n5784), .A(n5800) );
  nor02 U4504 ( .Y(n5801), .A0(n7486), .A1(n7377) );
  inv01 U4505 ( .Y(n5786), .A(n5801) );
  nor02 U4506 ( .Y(n5802), .A0(n7370), .A1(n7377) );
  inv01 U4507 ( .Y(n5788), .A(n5802) );
  nor02 U4508 ( .Y(n5803), .A0(n7486), .A1(n7487) );
  inv01 U4509 ( .Y(n5790), .A(n5803) );
  nor02 U4510 ( .Y(n5804), .A0(n7370), .A1(n7487) );
  inv01 U4511 ( .Y(n5792), .A(n5804) );
  nor02 U4512 ( .Y(n5805), .A0(n7486), .A1(n7377) );
  inv01 U4513 ( .Y(n5794), .A(n5805) );
  nor02 U4514 ( .Y(n5806), .A0(n7370), .A1(n7377) );
  inv01 U4515 ( .Y(n5796), .A(n5806) );
  nor02 U4516 ( .Y(n5807), .A0(n5781), .A1(n5783) );
  inv01 U4517 ( .Y(n5808), .A(n5807) );
  nor02 U4518 ( .Y(n5809), .A0(n5785), .A1(n5787) );
  inv01 U4519 ( .Y(n5810), .A(n5809) );
  nor02 U4520 ( .Y(n5811), .A0(n5808), .A1(n5810) );
  inv01 U4521 ( .Y(n5797), .A(n5811) );
  nor02 U4522 ( .Y(n5812), .A0(n5789), .A1(n5791) );
  inv01 U4523 ( .Y(n5813), .A(n5812) );
  nor02 U4524 ( .Y(n5814), .A0(n5793), .A1(n5795) );
  inv01 U4525 ( .Y(n5815), .A(n5814) );
  nor02 U4526 ( .Y(n5816), .A0(n5813), .A1(n5815) );
  inv01 U4527 ( .Y(n5798), .A(n5816) );
  inv04 U4528 ( .Y(n7377), .A(n7376) );
  inv02 U4529 ( .Y(n7487), .A(n6494) );
  inv02 U4530 ( .Y(n7488), .A(n6583) );
  nand02 U4531 ( .Y(n7460), .A0(n5817), .A1(n5818) );
  inv02 U4532 ( .Y(n5819), .A(n7463) );
  inv02 U4533 ( .Y(n5820), .A(n7462) );
  inv02 U4534 ( .Y(n5821), .A(n7461) );
  inv02 U4535 ( .Y(n5822), .A(n7368) );
  inv02 U4536 ( .Y(n5823), .A(n7369) );
  inv02 U4537 ( .Y(n5824), .A(n7370) );
  nand02 U4538 ( .Y(n5825), .A0(n5821), .A1(n5826) );
  nand02 U4539 ( .Y(n5827), .A0(n5822), .A1(n5828) );
  nand02 U4540 ( .Y(n5829), .A0(n5823), .A1(n5830) );
  nand02 U4541 ( .Y(n5831), .A0(n5823), .A1(n5832) );
  nand02 U4542 ( .Y(n5833), .A0(n5824), .A1(n5834) );
  nand02 U4543 ( .Y(n5835), .A0(n5824), .A1(n5836) );
  nand02 U4544 ( .Y(n5837), .A0(n5824), .A1(n5838) );
  nand02 U4545 ( .Y(n5839), .A0(n5824), .A1(n5840) );
  nand02 U4546 ( .Y(n5841), .A0(n5819), .A1(n5820) );
  inv01 U4547 ( .Y(n5826), .A(n5841) );
  nand02 U4548 ( .Y(n5842), .A0(n5819), .A1(n5820) );
  inv01 U4549 ( .Y(n5828), .A(n5842) );
  nand02 U4550 ( .Y(n5843), .A0(n5819), .A1(n5821) );
  inv01 U4551 ( .Y(n5830), .A(n5843) );
  nand02 U4552 ( .Y(n5844), .A0(n5819), .A1(n5822) );
  inv01 U4553 ( .Y(n5832), .A(n5844) );
  nand02 U4554 ( .Y(n5845), .A0(n5820), .A1(n5821) );
  inv01 U4555 ( .Y(n5834), .A(n5845) );
  nand02 U4556 ( .Y(n5846), .A0(n5820), .A1(n5822) );
  inv01 U4557 ( .Y(n5836), .A(n5846) );
  nand02 U4558 ( .Y(n5847), .A0(n5821), .A1(n5823) );
  inv01 U4559 ( .Y(n5838), .A(n5847) );
  nand02 U4560 ( .Y(n5848), .A0(n5822), .A1(n5823) );
  inv01 U4561 ( .Y(n5840), .A(n5848) );
  nand02 U4562 ( .Y(n5849), .A0(n5825), .A1(n5827) );
  inv01 U4563 ( .Y(n5850), .A(n5849) );
  nand02 U4564 ( .Y(n5851), .A0(n5829), .A1(n5831) );
  inv01 U4565 ( .Y(n5852), .A(n5851) );
  nand02 U4566 ( .Y(n5853), .A0(n5850), .A1(n5852) );
  inv01 U4567 ( .Y(n5817), .A(n5853) );
  nand02 U4568 ( .Y(n5854), .A0(n5833), .A1(n5835) );
  inv01 U4569 ( .Y(n5855), .A(n5854) );
  nand02 U4570 ( .Y(n5856), .A0(n5837), .A1(n5839) );
  inv01 U4571 ( .Y(n5857), .A(n5856) );
  nand02 U4572 ( .Y(n5858), .A0(n5855), .A1(n5857) );
  inv01 U4573 ( .Y(n5818), .A(n5858) );
  nand02 U4574 ( .Y(n7503), .A0(n5859), .A1(n5860) );
  inv02 U4575 ( .Y(n5861), .A(n7458) );
  inv02 U4576 ( .Y(n5862), .A(n7447) );
  inv02 U4577 ( .Y(n5863), .A(n7481) );
  inv02 U4578 ( .Y(n5864), .A(n7368) );
  inv02 U4579 ( .Y(n5865), .A(n7369) );
  inv02 U4580 ( .Y(n5866), .A(n7370) );
  nand02 U4581 ( .Y(n5867), .A0(n5863), .A1(n5868) );
  nand02 U4582 ( .Y(n5869), .A0(n5864), .A1(n5870) );
  nand02 U4583 ( .Y(n5871), .A0(n5865), .A1(n5872) );
  nand02 U4584 ( .Y(n5873), .A0(n5865), .A1(n5874) );
  nand02 U4585 ( .Y(n5875), .A0(n5866), .A1(n5876) );
  nand02 U4586 ( .Y(n5877), .A0(n5866), .A1(n5878) );
  nand02 U4587 ( .Y(n5879), .A0(n5866), .A1(n5880) );
  nand02 U4588 ( .Y(n5881), .A0(n5866), .A1(n5882) );
  nand02 U4589 ( .Y(n5883), .A0(n5861), .A1(n5862) );
  inv01 U4590 ( .Y(n5868), .A(n5883) );
  nand02 U4591 ( .Y(n5884), .A0(n5861), .A1(n5862) );
  inv01 U4592 ( .Y(n5870), .A(n5884) );
  nand02 U4593 ( .Y(n5885), .A0(n5861), .A1(n5863) );
  inv01 U4594 ( .Y(n5872), .A(n5885) );
  nand02 U4595 ( .Y(n5886), .A0(n5861), .A1(n5864) );
  inv01 U4596 ( .Y(n5874), .A(n5886) );
  nand02 U4597 ( .Y(n5887), .A0(n5862), .A1(n5863) );
  inv01 U4598 ( .Y(n5876), .A(n5887) );
  nand02 U4599 ( .Y(n5888), .A0(n5862), .A1(n5864) );
  inv01 U4600 ( .Y(n5878), .A(n5888) );
  nand02 U4601 ( .Y(n5889), .A0(n5863), .A1(n5865) );
  inv01 U4602 ( .Y(n5880), .A(n5889) );
  nand02 U4603 ( .Y(n5890), .A0(n5864), .A1(n5865) );
  inv01 U4604 ( .Y(n5882), .A(n5890) );
  nand02 U4605 ( .Y(n5891), .A0(n5867), .A1(n5869) );
  inv01 U4606 ( .Y(n5892), .A(n5891) );
  nand02 U4607 ( .Y(n5893), .A0(n5871), .A1(n5873) );
  inv01 U4608 ( .Y(n5894), .A(n5893) );
  nand02 U4609 ( .Y(n5895), .A0(n5892), .A1(n5894) );
  inv01 U4610 ( .Y(n5859), .A(n5895) );
  nand02 U4611 ( .Y(n5896), .A0(n5875), .A1(n5877) );
  inv01 U4612 ( .Y(n5897), .A(n5896) );
  nand02 U4613 ( .Y(n5898), .A0(n5879), .A1(n5881) );
  inv01 U4614 ( .Y(n5899), .A(n5898) );
  nand02 U4615 ( .Y(n5900), .A0(n5897), .A1(n5899) );
  inv01 U4616 ( .Y(n5860), .A(n5900) );
  nand02 U4617 ( .Y(n7445), .A0(n5901), .A1(n5902) );
  inv02 U4618 ( .Y(n5903), .A(n7451) );
  inv02 U4619 ( .Y(n5904), .A(n7449) );
  inv02 U4620 ( .Y(n5905), .A(n7447) );
  inv02 U4621 ( .Y(n5906), .A(n7368) );
  inv02 U4622 ( .Y(n5907), .A(n7369) );
  inv02 U4623 ( .Y(n5908), .A(n7370) );
  nand02 U4624 ( .Y(n5909), .A0(n5905), .A1(n5910) );
  nand02 U4625 ( .Y(n5911), .A0(n5906), .A1(n5912) );
  nand02 U4626 ( .Y(n5913), .A0(n5907), .A1(n5914) );
  nand02 U4627 ( .Y(n5915), .A0(n5907), .A1(n5916) );
  nand02 U4628 ( .Y(n5917), .A0(n5908), .A1(n5918) );
  nand02 U4629 ( .Y(n5919), .A0(n5908), .A1(n5920) );
  nand02 U4630 ( .Y(n5921), .A0(n5908), .A1(n5922) );
  nand02 U4631 ( .Y(n5923), .A0(n5908), .A1(n5924) );
  nand02 U4632 ( .Y(n5925), .A0(n5903), .A1(n5904) );
  inv01 U4633 ( .Y(n5910), .A(n5925) );
  nand02 U4634 ( .Y(n5926), .A0(n5903), .A1(n5904) );
  inv01 U4635 ( .Y(n5912), .A(n5926) );
  nand02 U4636 ( .Y(n5927), .A0(n5903), .A1(n5905) );
  inv01 U4637 ( .Y(n5914), .A(n5927) );
  nand02 U4638 ( .Y(n5928), .A0(n5903), .A1(n5906) );
  inv01 U4639 ( .Y(n5916), .A(n5928) );
  nand02 U4640 ( .Y(n5929), .A0(n5904), .A1(n5905) );
  inv01 U4641 ( .Y(n5918), .A(n5929) );
  nand02 U4642 ( .Y(n5930), .A0(n5904), .A1(n5906) );
  inv01 U4643 ( .Y(n5920), .A(n5930) );
  nand02 U4644 ( .Y(n5931), .A0(n5905), .A1(n5907) );
  inv01 U4645 ( .Y(n5922), .A(n5931) );
  nand02 U4646 ( .Y(n5932), .A0(n5906), .A1(n5907) );
  inv01 U4647 ( .Y(n5924), .A(n5932) );
  nand02 U4648 ( .Y(n5933), .A0(n5909), .A1(n5911) );
  inv01 U4649 ( .Y(n5934), .A(n5933) );
  nand02 U4650 ( .Y(n5935), .A0(n5913), .A1(n5915) );
  inv01 U4651 ( .Y(n5936), .A(n5935) );
  nand02 U4652 ( .Y(n5937), .A0(n5934), .A1(n5936) );
  inv01 U4653 ( .Y(n5901), .A(n5937) );
  nand02 U4654 ( .Y(n5938), .A0(n5917), .A1(n5919) );
  inv01 U4655 ( .Y(n5939), .A(n5938) );
  nand02 U4656 ( .Y(n5940), .A0(n5921), .A1(n5923) );
  inv01 U4657 ( .Y(n5941), .A(n5940) );
  nand02 U4658 ( .Y(n5942), .A0(n5939), .A1(n5941) );
  inv01 U4659 ( .Y(n5902), .A(n5942) );
  inv01 U4660 ( .Y(n7513), .A(n5943) );
  nor02 U4661 ( .Y(n5944), .A0(n7467), .A1(n5945) );
  nor02 U4662 ( .Y(n5946), .A0(n7467), .A1(n5947) );
  nor02 U4663 ( .Y(n5948), .A0(n7467), .A1(n5949) );
  nor02 U4664 ( .Y(n5950), .A0(n7467), .A1(n5951) );
  nor02 U4665 ( .Y(n5952), .A0(n7370), .A1(n5953) );
  nor02 U4666 ( .Y(n5954), .A0(n7370), .A1(n5955) );
  nor02 U4667 ( .Y(n5956), .A0(n7370), .A1(n5957) );
  nor02 U4668 ( .Y(n5958), .A0(n7370), .A1(n5959) );
  nor02 U4669 ( .Y(n5943), .A0(n5960), .A1(n5961) );
  nor02 U4670 ( .Y(n5962), .A0(n7494), .A1(n7461) );
  inv01 U4671 ( .Y(n5945), .A(n5962) );
  nor02 U4672 ( .Y(n5963), .A0(n7368), .A1(n7461) );
  inv01 U4673 ( .Y(n5947), .A(n5963) );
  nor02 U4674 ( .Y(n5964), .A0(n7494), .A1(n7369) );
  inv01 U4675 ( .Y(n5949), .A(n5964) );
  nor02 U4676 ( .Y(n5965), .A0(n7368), .A1(n7369) );
  inv01 U4677 ( .Y(n5951), .A(n5965) );
  nor02 U4678 ( .Y(n5966), .A0(n7494), .A1(n7461) );
  inv01 U4679 ( .Y(n5953), .A(n5966) );
  nor02 U4680 ( .Y(n5967), .A0(n7368), .A1(n7461) );
  inv01 U4681 ( .Y(n5955), .A(n5967) );
  nor02 U4682 ( .Y(n5968), .A0(n7494), .A1(n7369) );
  inv01 U4683 ( .Y(n5957), .A(n5968) );
  nor02 U4684 ( .Y(n5969), .A0(n7368), .A1(n7369) );
  inv01 U4685 ( .Y(n5959), .A(n5969) );
  nor02 U4686 ( .Y(n5970), .A0(n5944), .A1(n5946) );
  inv01 U4687 ( .Y(n5971), .A(n5970) );
  nor02 U4688 ( .Y(n5972), .A0(n5948), .A1(n5950) );
  inv01 U4689 ( .Y(n5973), .A(n5972) );
  nor02 U4690 ( .Y(n5974), .A0(n5971), .A1(n5973) );
  inv01 U4691 ( .Y(n5960), .A(n5974) );
  nor02 U4692 ( .Y(n5975), .A0(n5952), .A1(n5954) );
  inv01 U4693 ( .Y(n5976), .A(n5975) );
  nor02 U4694 ( .Y(n5977), .A0(n5956), .A1(n5958) );
  inv01 U4695 ( .Y(n5978), .A(n5977) );
  nor02 U4696 ( .Y(n5979), .A0(n5976), .A1(n5978) );
  inv01 U4697 ( .Y(n5961), .A(n5979) );
  inv02 U4698 ( .Y(n7451), .A(n6595) );
  inv08 U4699 ( .Y(n7368), .A(n5486) );
  nand02 U4700 ( .Y(n7479), .A0(n5980), .A1(n5981) );
  inv02 U4701 ( .Y(n5982), .A(n7447) );
  inv02 U4702 ( .Y(n5983), .A(n7451) );
  inv02 U4703 ( .Y(n5984), .A(n7458) );
  inv02 U4704 ( .Y(n5985), .A(n7368) );
  inv02 U4705 ( .Y(n5986), .A(n7369) );
  inv02 U4706 ( .Y(n5987), .A(n7370) );
  nand02 U4707 ( .Y(n5988), .A0(n5984), .A1(n5989) );
  nand02 U4708 ( .Y(n5990), .A0(n5985), .A1(n5991) );
  nand02 U4709 ( .Y(n5992), .A0(n5986), .A1(n5993) );
  nand02 U4710 ( .Y(n5994), .A0(n5986), .A1(n5995) );
  nand02 U4711 ( .Y(n5996), .A0(n5987), .A1(n5997) );
  nand02 U4712 ( .Y(n5998), .A0(n5987), .A1(n5999) );
  nand02 U4713 ( .Y(n6000), .A0(n5987), .A1(n6001) );
  nand02 U4714 ( .Y(n6002), .A0(n5987), .A1(n6003) );
  nand02 U4715 ( .Y(n6004), .A0(n5982), .A1(n5983) );
  inv01 U4716 ( .Y(n5989), .A(n6004) );
  nand02 U4717 ( .Y(n6005), .A0(n5982), .A1(n5983) );
  inv01 U4718 ( .Y(n5991), .A(n6005) );
  nand02 U4719 ( .Y(n6006), .A0(n5982), .A1(n5984) );
  inv01 U4720 ( .Y(n5993), .A(n6006) );
  nand02 U4721 ( .Y(n6007), .A0(n5982), .A1(n5985) );
  inv01 U4722 ( .Y(n5995), .A(n6007) );
  nand02 U4723 ( .Y(n6008), .A0(n5983), .A1(n5984) );
  inv01 U4724 ( .Y(n5997), .A(n6008) );
  nand02 U4725 ( .Y(n6009), .A0(n5983), .A1(n5985) );
  inv01 U4726 ( .Y(n5999), .A(n6009) );
  nand02 U4727 ( .Y(n6010), .A0(n5984), .A1(n5986) );
  inv01 U4728 ( .Y(n6001), .A(n6010) );
  nand02 U4729 ( .Y(n6011), .A0(n5985), .A1(n5986) );
  inv01 U4730 ( .Y(n6003), .A(n6011) );
  nand02 U4731 ( .Y(n6012), .A0(n5988), .A1(n5990) );
  inv01 U4732 ( .Y(n6013), .A(n6012) );
  nand02 U4733 ( .Y(n6014), .A0(n5992), .A1(n5994) );
  inv01 U4734 ( .Y(n6015), .A(n6014) );
  nand02 U4735 ( .Y(n6016), .A0(n6013), .A1(n6015) );
  inv01 U4736 ( .Y(n5980), .A(n6016) );
  nand02 U4737 ( .Y(n6017), .A0(n5996), .A1(n5998) );
  inv01 U4738 ( .Y(n6018), .A(n6017) );
  nand02 U4739 ( .Y(n6019), .A0(n6000), .A1(n6002) );
  inv01 U4740 ( .Y(n6020), .A(n6019) );
  nand02 U4741 ( .Y(n6021), .A0(n6018), .A1(n6020) );
  inv01 U4742 ( .Y(n5981), .A(n6021) );
  nand02 U4743 ( .Y(n7519), .A0(n6022), .A1(n6023) );
  inv02 U4744 ( .Y(n6024), .A(n7476) );
  inv02 U4745 ( .Y(n6025), .A(n7471) );
  inv02 U4746 ( .Y(n6026), .A(n7500) );
  inv02 U4747 ( .Y(n6027), .A(n7368) );
  inv02 U4748 ( .Y(n6028), .A(n7369) );
  inv02 U4749 ( .Y(n6029), .A(n7370) );
  nand02 U4750 ( .Y(n6030), .A0(n6026), .A1(n6031) );
  nand02 U4751 ( .Y(n6032), .A0(n6027), .A1(n6033) );
  nand02 U4752 ( .Y(n6034), .A0(n6028), .A1(n6035) );
  nand02 U4753 ( .Y(n6036), .A0(n6028), .A1(n6037) );
  nand02 U4754 ( .Y(n6038), .A0(n6029), .A1(n6039) );
  nand02 U4755 ( .Y(n6040), .A0(n6029), .A1(n6041) );
  nand02 U4756 ( .Y(n6042), .A0(n6029), .A1(n6043) );
  nand02 U4757 ( .Y(n6044), .A0(n6029), .A1(n6045) );
  nand02 U4758 ( .Y(n6046), .A0(n6024), .A1(n6025) );
  inv01 U4759 ( .Y(n6031), .A(n6046) );
  nand02 U4760 ( .Y(n6047), .A0(n6024), .A1(n6025) );
  inv01 U4761 ( .Y(n6033), .A(n6047) );
  nand02 U4762 ( .Y(n6048), .A0(n6024), .A1(n6026) );
  inv01 U4763 ( .Y(n6035), .A(n6048) );
  nand02 U4764 ( .Y(n6049), .A0(n6024), .A1(n6027) );
  inv01 U4765 ( .Y(n6037), .A(n6049) );
  nand02 U4766 ( .Y(n6050), .A0(n6025), .A1(n6026) );
  inv01 U4767 ( .Y(n6039), .A(n6050) );
  nand02 U4768 ( .Y(n6051), .A0(n6025), .A1(n6027) );
  inv01 U4769 ( .Y(n6041), .A(n6051) );
  nand02 U4770 ( .Y(n6052), .A0(n6026), .A1(n6028) );
  inv01 U4771 ( .Y(n6043), .A(n6052) );
  nand02 U4772 ( .Y(n6053), .A0(n6027), .A1(n6028) );
  inv01 U4773 ( .Y(n6045), .A(n6053) );
  nand02 U4774 ( .Y(n6054), .A0(n6030), .A1(n6032) );
  inv01 U4775 ( .Y(n6055), .A(n6054) );
  nand02 U4776 ( .Y(n6056), .A0(n6034), .A1(n6036) );
  inv01 U4777 ( .Y(n6057), .A(n6056) );
  nand02 U4778 ( .Y(n6058), .A0(n6055), .A1(n6057) );
  inv01 U4779 ( .Y(n6022), .A(n6058) );
  nand02 U4780 ( .Y(n6059), .A0(n6038), .A1(n6040) );
  inv01 U4781 ( .Y(n6060), .A(n6059) );
  nand02 U4782 ( .Y(n6061), .A0(n6042), .A1(n6044) );
  inv01 U4783 ( .Y(n6062), .A(n6061) );
  nand02 U4784 ( .Y(n6063), .A0(n6060), .A1(n6062) );
  inv01 U4785 ( .Y(n6023), .A(n6063) );
  nand02 U4786 ( .Y(n7497), .A0(n6064), .A1(n6065) );
  inv02 U4787 ( .Y(n6066), .A(n7471) );
  inv02 U4788 ( .Y(n6067), .A(n7473) );
  inv02 U4789 ( .Y(n6068), .A(n7476) );
  inv02 U4790 ( .Y(n6069), .A(n7368) );
  inv02 U4791 ( .Y(n6070), .A(n7369) );
  inv02 U4792 ( .Y(n6071), .A(n7370) );
  nand02 U4793 ( .Y(n6072), .A0(n6068), .A1(n6073) );
  nand02 U4794 ( .Y(n6074), .A0(n6069), .A1(n6075) );
  nand02 U4795 ( .Y(n6076), .A0(n6070), .A1(n6077) );
  nand02 U4796 ( .Y(n6078), .A0(n6070), .A1(n6079) );
  nand02 U4797 ( .Y(n6080), .A0(n6071), .A1(n6081) );
  nand02 U4798 ( .Y(n6082), .A0(n6071), .A1(n6083) );
  nand02 U4799 ( .Y(n6084), .A0(n6071), .A1(n6085) );
  nand02 U4800 ( .Y(n6086), .A0(n6071), .A1(n6087) );
  nand02 U4801 ( .Y(n6088), .A0(n6066), .A1(n6067) );
  inv01 U4802 ( .Y(n6073), .A(n6088) );
  nand02 U4803 ( .Y(n6089), .A0(n6066), .A1(n6067) );
  inv01 U4804 ( .Y(n6075), .A(n6089) );
  nand02 U4805 ( .Y(n6090), .A0(n6066), .A1(n6068) );
  inv01 U4806 ( .Y(n6077), .A(n6090) );
  nand02 U4807 ( .Y(n6091), .A0(n6066), .A1(n6069) );
  inv01 U4808 ( .Y(n6079), .A(n6091) );
  nand02 U4809 ( .Y(n6092), .A0(n6067), .A1(n6068) );
  inv01 U4810 ( .Y(n6081), .A(n6092) );
  nand02 U4811 ( .Y(n6093), .A0(n6067), .A1(n6069) );
  inv01 U4812 ( .Y(n6083), .A(n6093) );
  nand02 U4813 ( .Y(n6094), .A0(n6068), .A1(n6070) );
  inv01 U4814 ( .Y(n6085), .A(n6094) );
  nand02 U4815 ( .Y(n6095), .A0(n6069), .A1(n6070) );
  inv01 U4816 ( .Y(n6087), .A(n6095) );
  nand02 U4817 ( .Y(n6096), .A0(n6072), .A1(n6074) );
  inv01 U4818 ( .Y(n6097), .A(n6096) );
  nand02 U4819 ( .Y(n6098), .A0(n6076), .A1(n6078) );
  inv01 U4820 ( .Y(n6099), .A(n6098) );
  nand02 U4821 ( .Y(n6100), .A0(n6097), .A1(n6099) );
  inv01 U4822 ( .Y(n6064), .A(n6100) );
  nand02 U4823 ( .Y(n6101), .A0(n6080), .A1(n6082) );
  inv01 U4824 ( .Y(n6102), .A(n6101) );
  nand02 U4825 ( .Y(n6103), .A0(n6084), .A1(n6086) );
  inv01 U4826 ( .Y(n6104), .A(n6103) );
  nand02 U4827 ( .Y(n6105), .A0(n6102), .A1(n6104) );
  inv01 U4828 ( .Y(n6065), .A(n6105) );
  buf08 U4829 ( .Y(n6106), .A(n7422) );
  inv04 U4830 ( .Y(n7422), .A(n7791) );
  buf12 U4831 ( .Y(n6107), .A(n7410) );
  inv02 U4832 ( .Y(n7410), .A(n8003) );
  nor02 U4833 ( .Y(n6108), .A0(n7639), .A1(n7380) );
  inv02 U4834 ( .Y(n7639), .A(n7375) );
  or04 U4835 ( .Y(n6109), .A0(n7696), .A1(n7697), .A2(n7698), .A3(n7699) );
  inv02 U4836 ( .Y(n6110), .A(n6109) );
  or04 U4837 ( .Y(n6111), .A0(n7714), .A1(n7715), .A2(n7716), .A3(n7717) );
  inv02 U4838 ( .Y(n6112), .A(n6111) );
  inv02 U4839 ( .Y(n7745), .A(n6113) );
  inv01 U4840 ( .Y(n6114), .A(n3331) );
  inv01 U4841 ( .Y(n6115), .A(n7765) );
  inv01 U4842 ( .Y(n6116), .A(n3111) );
  inv02 U4843 ( .Y(n6117), .A(n7764) );
  nand02 U4844 ( .Y(n6113), .A0(n6118), .A1(n6119) );
  nand02 U4845 ( .Y(n6120), .A0(n6114), .A1(n6115) );
  inv01 U4846 ( .Y(n6118), .A(n6120) );
  nand02 U4847 ( .Y(n6121), .A0(n6116), .A1(n6117) );
  inv01 U4848 ( .Y(n6119), .A(n6121) );
  inv02 U4849 ( .Y(n7718), .A(n6122) );
  inv01 U4850 ( .Y(n6123), .A(n3089) );
  inv01 U4851 ( .Y(n6124), .A(n7741) );
  inv01 U4852 ( .Y(n6125), .A(n7740) );
  inv02 U4853 ( .Y(n6126), .A(n7739) );
  nand02 U4854 ( .Y(n6122), .A0(n6127), .A1(n6128) );
  nand02 U4855 ( .Y(n6129), .A0(n6123), .A1(n6124) );
  inv01 U4856 ( .Y(n6127), .A(n6129) );
  nand02 U4857 ( .Y(n6130), .A0(n6125), .A1(n6126) );
  inv01 U4858 ( .Y(n6128), .A(n6130) );
  inv02 U4859 ( .Y(n6132), .A(n6131) );
  nor02 U4860 ( .Y(n7682), .A0(n6133), .A1(n6134) );
  nor02 U4861 ( .Y(n6135), .A0(n7692), .A1(n7693) );
  inv01 U4862 ( .Y(n6133), .A(n6135) );
  nor02 U4863 ( .Y(n6136), .A0(n7694), .A1(n7695) );
  inv01 U4864 ( .Y(n6134), .A(n6136) );
  nor02 U4865 ( .Y(n7700), .A0(n6137), .A1(n6138) );
  nor02 U4866 ( .Y(n6139), .A0(n7710), .A1(n7711) );
  inv01 U4867 ( .Y(n6137), .A(n6139) );
  nor02 U4868 ( .Y(n6140), .A0(n7712), .A1(n7713) );
  inv01 U4869 ( .Y(n6138), .A(n6140) );
  or04 U4870 ( .Y(n6141), .A0(n7706), .A1(n7707), .A2(n7708), .A3(n7709) );
  inv01 U4871 ( .Y(n6142), .A(n6141) );
  or04 U4872 ( .Y(n6143), .A0(n7688), .A1(n7689), .A2(n7690), .A3(n7691) );
  inv01 U4873 ( .Y(n6144), .A(n6143) );
  inv02 U4874 ( .Y(n7758), .A(r1_2_1_) );
  inv04 U4875 ( .Y(n7719), .A(n6145) );
  inv01 U4876 ( .Y(n6146), .A(n3121) );
  inv01 U4877 ( .Y(n6147), .A(n7735) );
  inv01 U4878 ( .Y(n6148), .A(n7734) );
  inv01 U4879 ( .Y(n6149), .A(n7733) );
  nand02 U4880 ( .Y(n6145), .A0(n6150), .A1(n6151) );
  nand02 U4881 ( .Y(n6152), .A0(n6146), .A1(n6147) );
  inv02 U4882 ( .Y(n6150), .A(n6152) );
  nand02 U4883 ( .Y(n6153), .A0(n6148), .A1(n6149) );
  inv02 U4884 ( .Y(n6151), .A(n6153) );
  inv04 U4885 ( .Y(n7746), .A(n6154) );
  inv01 U4886 ( .Y(n6155), .A(n3113) );
  inv01 U4887 ( .Y(n6156), .A(n3109) );
  inv01 U4888 ( .Y(n6157), .A(n7760) );
  inv01 U4889 ( .Y(n6158), .A(n7759) );
  nand02 U4890 ( .Y(n6154), .A0(n6159), .A1(n6160) );
  nand02 U4891 ( .Y(n6161), .A0(n6155), .A1(n6156) );
  inv02 U4892 ( .Y(n6159), .A(n6161) );
  nand02 U4893 ( .Y(n6162), .A0(n6157), .A1(n6158) );
  inv02 U4894 ( .Y(n6160), .A(n6162) );
  inv02 U4895 ( .Y(n6164), .A(n6163) );
  inv02 U4896 ( .Y(n6166), .A(n6165) );
  inv02 U4897 ( .Y(n6168), .A(n6167) );
  inv02 U4898 ( .Y(n6170), .A(n6169) );
  inv02 U4899 ( .Y(n6172), .A(n6171) );
  inv02 U4900 ( .Y(n6174), .A(n6173) );
  inv02 U4901 ( .Y(n6176), .A(n6175) );
  inv02 U4902 ( .Y(n6178), .A(n6177) );
  inv02 U4903 ( .Y(n6180), .A(n6179) );
  inv02 U4904 ( .Y(n6182), .A(n6181) );
  inv02 U4905 ( .Y(n6184), .A(n6183) );
  inv04 U4906 ( .Y(n7747), .A(n6185) );
  inv01 U4907 ( .Y(n6186), .A(n3117) );
  inv01 U4908 ( .Y(n6187), .A(n7755) );
  inv01 U4909 ( .Y(n6188), .A(n3333) );
  inv02 U4910 ( .Y(n6189), .A(n7754) );
  nand02 U4911 ( .Y(n6185), .A0(n6190), .A1(n6191) );
  nand02 U4912 ( .Y(n6192), .A0(n6186), .A1(n6187) );
  inv02 U4913 ( .Y(n6190), .A(n6192) );
  nand02 U4914 ( .Y(n6193), .A0(n6188), .A1(n6189) );
  inv02 U4915 ( .Y(n6191), .A(n6193) );
  inv01 U4916 ( .Y(n7720), .A(n6194) );
  inv01 U4917 ( .Y(n6195), .A(n7729) );
  inv01 U4918 ( .Y(n6196), .A(n7728) );
  inv01 U4919 ( .Y(n6197), .A(n3107) );
  inv01 U4920 ( .Y(n6198), .A(n7727) );
  nand02 U4921 ( .Y(n6194), .A0(n6199), .A1(n6200) );
  nand02 U4922 ( .Y(n6201), .A0(n6195), .A1(n6196) );
  inv01 U4923 ( .Y(n6199), .A(n6201) );
  nand02 U4924 ( .Y(n6202), .A0(n6197), .A1(n6198) );
  inv01 U4925 ( .Y(n6200), .A(n6202) );
  buf04 U4926 ( .Y(n6203), .A(n8002) );
  inv02 U4927 ( .Y(n7640), .A(n7384) );
  buf04 U4928 ( .Y(n6204), .A(n7381) );
  nor02 U4929 ( .Y(n7683), .A0(n6205), .A1(n6206) );
  nor02 U4930 ( .Y(n6207), .A0(n7684), .A1(n7685) );
  inv02 U4931 ( .Y(n6205), .A(n6207) );
  nor02 U4932 ( .Y(n6208), .A0(n7686), .A1(n7687) );
  inv01 U4933 ( .Y(n6206), .A(n6208) );
  nor02 U4934 ( .Y(n7701), .A0(n6209), .A1(n6210) );
  nor02 U4935 ( .Y(n6211), .A0(n7702), .A1(n7703) );
  inv02 U4936 ( .Y(n6209), .A(n6211) );
  nor02 U4937 ( .Y(n6212), .A0(n7704), .A1(n7705) );
  inv01 U4938 ( .Y(n6210), .A(n6212) );
  inv01 U4939 ( .Y(n7721), .A(n6213) );
  inv01 U4940 ( .Y(n6214), .A(n3119) );
  inv01 U4941 ( .Y(n6215), .A(n3115) );
  inv01 U4942 ( .Y(n6216), .A(n7723) );
  inv01 U4943 ( .Y(n6217), .A(n7722) );
  nand02 U4944 ( .Y(n6213), .A0(n6218), .A1(n6219) );
  nand02 U4945 ( .Y(n6220), .A0(n6214), .A1(n6215) );
  inv01 U4946 ( .Y(n6218), .A(n6220) );
  nand02 U4947 ( .Y(n6221), .A0(n6216), .A1(n6217) );
  inv01 U4948 ( .Y(n6219), .A(n6221) );
  inv04 U4949 ( .Y(n7748), .A(n6222) );
  inv01 U4950 ( .Y(n6223), .A(n3101) );
  inv01 U4951 ( .Y(n6224), .A(n3099) );
  inv01 U4952 ( .Y(n6225), .A(n7750) );
  inv01 U4953 ( .Y(n6226), .A(n7749) );
  nand02 U4954 ( .Y(n6222), .A0(n6227), .A1(n6228) );
  nand02 U4955 ( .Y(n6229), .A0(n6223), .A1(n6224) );
  inv02 U4956 ( .Y(n6227), .A(n6229) );
  nand02 U4957 ( .Y(n6230), .A0(n6225), .A1(n6226) );
  inv02 U4958 ( .Y(n6228), .A(n6230) );
  inv02 U4959 ( .Y(n6232), .A(n6231) );
  inv02 U4960 ( .Y(n6234), .A(n6233) );
  inv02 U4961 ( .Y(n6236), .A(n6235) );
  inv02 U4962 ( .Y(n6238), .A(n6237) );
  inv02 U4963 ( .Y(n6240), .A(n6239) );
  inv02 U4964 ( .Y(n6242), .A(n6241) );
  inv02 U4965 ( .Y(n6244), .A(n6243) );
  inv02 U4966 ( .Y(n6246), .A(n6245) );
  inv02 U4967 ( .Y(n6248), .A(n6247) );
  inv02 U4968 ( .Y(n6250), .A(n6249) );
  inv02 U4969 ( .Y(n6252), .A(n6251) );
  inv02 U4970 ( .Y(n7737), .A(r1_2_50_) );
  inv02 U4971 ( .Y(n7768), .A(r1_2_31_) );
  inv02 U4972 ( .Y(n7724), .A(r1_2_37_) );
  inv02 U4973 ( .Y(n7736), .A(r1_2_49_) );
  inv02 U4974 ( .Y(n7742), .A(r1_2_7_) );
  inv02 U4975 ( .Y(n7762), .A(r1_2_27_) );
  inv02 U4976 ( .Y(n7761), .A(r1_2_25_) );
  inv02 U4977 ( .Y(n7725), .A(r1_2_39_) );
  inv02 U4978 ( .Y(n7752), .A(r1_2_15_) );
  inv02 U4979 ( .Y(n7732), .A(r1_2_43_) );
  inv02 U4980 ( .Y(n7751), .A(r1_2_13_) );
  inv02 U4981 ( .Y(n7756), .A(r1_2_19_) );
  inv02 U4982 ( .Y(n7767), .A(r1_2_32_) );
  inv02 U4983 ( .Y(n7731), .A(r1_2_44_) );
  inv02 U4984 ( .Y(n7743), .A(r1_2_9_) );
  inv02 U4985 ( .Y(n7757), .A(r1_2_20_) );
  inv02 U4986 ( .Y(n7730), .A(r1_2_42_) );
  inv02 U4987 ( .Y(n7766), .A(r1_2_30_) );
  inv02 U4988 ( .Y(n7726), .A(r1_2_38_) );
  inv02 U4989 ( .Y(n7753), .A(r1_2_14_) );
  inv02 U4990 ( .Y(n7744), .A(r1_2_8_) );
  inv02 U4991 ( .Y(n7763), .A(r1_2_26_) );
  inv02 U4992 ( .Y(n7738), .A(r1_2_4_) );
  buf02 U4993 ( .Y(n6253), .A(s_rad_i_8_) );
  buf02 U4994 ( .Y(n6256), .A(s_rad_i_8_) );
  buf02 U4995 ( .Y(n6254), .A(s_rad_i_8_) );
  buf02 U4996 ( .Y(n6255), .A(s_rad_i_8_) );
  buf02 U4997 ( .Y(n6257), .A(s_rad_i_12_) );
  buf02 U4998 ( .Y(n6260), .A(s_rad_i_12_) );
  buf02 U4999 ( .Y(n6258), .A(s_rad_i_12_) );
  buf02 U5000 ( .Y(n6259), .A(s_rad_i_12_) );
  buf02 U5001 ( .Y(n6261), .A(s_rad_i_24_) );
  buf02 U5002 ( .Y(n6264), .A(s_rad_i_24_) );
  buf02 U5003 ( .Y(n6262), .A(s_rad_i_24_) );
  buf02 U5004 ( .Y(n6263), .A(s_rad_i_24_) );
  buf02 U5005 ( .Y(n6265), .A(s_rad_i_44_) );
  buf02 U5006 ( .Y(n6267), .A(s_rad_i_44_) );
  buf02 U5007 ( .Y(n6266), .A(s_rad_i_44_) );
  buf02 U5008 ( .Y(n6268), .A(s_rad_i_9_) );
  buf02 U5009 ( .Y(n6270), .A(s_rad_i_9_) );
  buf02 U5010 ( .Y(n6269), .A(s_rad_i_9_) );
  buf02 U5011 ( .Y(n6271), .A(s_rad_i_38_) );
  buf02 U5012 ( .Y(n6273), .A(s_rad_i_38_) );
  buf02 U5013 ( .Y(n6272), .A(s_rad_i_38_) );
  buf02 U5014 ( .Y(n6274), .A(s_rad_i_50_) );
  buf02 U5015 ( .Y(n6276), .A(s_rad_i_50_) );
  buf02 U5016 ( .Y(n6275), .A(s_rad_i_50_) );
  buf02 U5017 ( .Y(n6277), .A(s_rad_i_20_) );
  buf02 U5018 ( .Y(n6279), .A(s_rad_i_20_) );
  buf02 U5019 ( .Y(n6278), .A(s_rad_i_20_) );
  buf02 U5020 ( .Y(n6280), .A(s_rad_i_32_) );
  buf02 U5021 ( .Y(n6282), .A(s_rad_i_32_) );
  buf02 U5022 ( .Y(n6281), .A(s_rad_i_32_) );
  buf02 U5023 ( .Y(n6283), .A(s_rad_i_4_) );
  buf02 U5024 ( .Y(n6285), .A(s_rad_i_4_) );
  buf02 U5025 ( .Y(n6284), .A(s_rad_i_4_) );
  buf02 U5026 ( .Y(n6286), .A(s_rad_i_14_) );
  buf02 U5027 ( .Y(n6288), .A(s_rad_i_14_) );
  buf02 U5028 ( .Y(n6287), .A(s_rad_i_14_) );
  buf02 U5029 ( .Y(n6289), .A(s_rad_i_26_) );
  buf02 U5030 ( .Y(n6291), .A(s_rad_i_26_) );
  buf02 U5031 ( .Y(n6290), .A(s_rad_i_26_) );
  buf02 U5032 ( .Y(n6292), .A(s_rad_i_42_) );
  buf02 U5033 ( .Y(n6294), .A(s_rad_i_42_) );
  buf02 U5034 ( .Y(n6293), .A(s_rad_i_42_) );
  ao221 U5035 ( .Y(n6295), .A0(n7581), .A1(n7390), .B0(n7621), .B1(n7374), 
        .C0(n7631) );
  inv01 U5036 ( .Y(n6296), .A(n6295) );
  ao221 U5037 ( .Y(n6297), .A0(n7595), .A1(n7388), .B0(n7589), .B1(n7390), 
        .C0(n7638) );
  inv01 U5038 ( .Y(n6298), .A(n6297) );
  ao221 U5039 ( .Y(n6299), .A0(n7608), .A1(n7384), .B0(n7609), .B1(n7388), 
        .C0(n7634) );
  inv01 U5040 ( .Y(n6300), .A(n6299) );
  inv02 U5041 ( .Y(n7464), .A(r0_46_) );
  inv02 U5042 ( .Y(n7453), .A(r0_48_) );
  inv02 U5043 ( .Y(n7465), .A(r0_47_) );
  nand02 U5044 ( .Y(n7502), .A0(n6301), .A1(n6302) );
  inv02 U5045 ( .Y(n6303), .A(n7580) );
  inv01 U5046 ( .Y(n6304), .A(n7388) );
  inv01 U5047 ( .Y(n6305), .A(n7390) );
  inv01 U5048 ( .Y(n6306), .A(n7525) );
  inv01 U5049 ( .Y(n6307), .A(n7549) );
  nand02 U5050 ( .Y(n6308), .A0(n6305), .A1(n6309) );
  nand02 U5051 ( .Y(n6310), .A0(n6306), .A1(n6311) );
  nand02 U5052 ( .Y(n6312), .A0(n6307), .A1(n6313) );
  nand02 U5053 ( .Y(n6314), .A0(n6307), .A1(n6315) );
  nand02 U5054 ( .Y(n6316), .A0(n6303), .A1(n6304) );
  inv01 U5055 ( .Y(n6309), .A(n6316) );
  nand02 U5056 ( .Y(n6317), .A0(n6303), .A1(n6304) );
  inv01 U5057 ( .Y(n6311), .A(n6317) );
  nand02 U5058 ( .Y(n6318), .A0(n6303), .A1(n6305) );
  inv01 U5059 ( .Y(n6313), .A(n6318) );
  nand02 U5060 ( .Y(n6319), .A0(n6303), .A1(n6306) );
  inv01 U5061 ( .Y(n6315), .A(n6319) );
  nand02 U5062 ( .Y(n6320), .A0(n6308), .A1(n6310) );
  inv01 U5063 ( .Y(n6301), .A(n6320) );
  nand02 U5064 ( .Y(n6321), .A0(n6312), .A1(n6314) );
  inv01 U5065 ( .Y(n6302), .A(n6321) );
  nand02 U5066 ( .Y(n7512), .A0(n6322), .A1(n6323) );
  inv02 U5067 ( .Y(n6324), .A(n7588) );
  inv01 U5068 ( .Y(n6325), .A(n7388) );
  inv01 U5069 ( .Y(n6326), .A(n7390) );
  inv01 U5070 ( .Y(n6327), .A(n7537) );
  inv01 U5071 ( .Y(n6328), .A(n7554) );
  nand02 U5072 ( .Y(n6329), .A0(n6326), .A1(n6330) );
  nand02 U5073 ( .Y(n6331), .A0(n6327), .A1(n6332) );
  nand02 U5074 ( .Y(n6333), .A0(n6328), .A1(n6334) );
  nand02 U5075 ( .Y(n6335), .A0(n6328), .A1(n6336) );
  nand02 U5076 ( .Y(n6337), .A0(n6324), .A1(n6325) );
  inv01 U5077 ( .Y(n6330), .A(n6337) );
  nand02 U5078 ( .Y(n6338), .A0(n6324), .A1(n6325) );
  inv01 U5079 ( .Y(n6332), .A(n6338) );
  nand02 U5080 ( .Y(n6339), .A0(n6324), .A1(n6326) );
  inv01 U5081 ( .Y(n6334), .A(n6339) );
  nand02 U5082 ( .Y(n6340), .A0(n6324), .A1(n6327) );
  inv01 U5083 ( .Y(n6336), .A(n6340) );
  nand02 U5084 ( .Y(n6341), .A0(n6329), .A1(n6331) );
  inv01 U5085 ( .Y(n6322), .A(n6341) );
  nand02 U5086 ( .Y(n6342), .A0(n6333), .A1(n6335) );
  inv01 U5087 ( .Y(n6323), .A(n6342) );
  nand02 U5088 ( .Y(n7496), .A0(n6343), .A1(n6344) );
  inv02 U5089 ( .Y(n6345), .A(n7576) );
  inv01 U5090 ( .Y(n6346), .A(n7388) );
  inv01 U5091 ( .Y(n6347), .A(n7390) );
  inv01 U5092 ( .Y(n6348), .A(n7521) );
  inv01 U5093 ( .Y(n6349), .A(n7543) );
  nand02 U5094 ( .Y(n6350), .A0(n6347), .A1(n6351) );
  nand02 U5095 ( .Y(n6352), .A0(n6348), .A1(n6353) );
  nand02 U5096 ( .Y(n6354), .A0(n6349), .A1(n6355) );
  nand02 U5097 ( .Y(n6356), .A0(n6349), .A1(n6357) );
  nand02 U5098 ( .Y(n6358), .A0(n6345), .A1(n6346) );
  inv01 U5099 ( .Y(n6351), .A(n6358) );
  nand02 U5100 ( .Y(n6359), .A0(n6345), .A1(n6346) );
  inv01 U5101 ( .Y(n6353), .A(n6359) );
  nand02 U5102 ( .Y(n6360), .A0(n6345), .A1(n6347) );
  inv01 U5103 ( .Y(n6355), .A(n6360) );
  nand02 U5104 ( .Y(n6361), .A0(n6345), .A1(n6348) );
  inv01 U5105 ( .Y(n6357), .A(n6361) );
  nand02 U5106 ( .Y(n6362), .A0(n6350), .A1(n6352) );
  inv01 U5107 ( .Y(n6343), .A(n6362) );
  nand02 U5108 ( .Y(n6363), .A0(n6354), .A1(n6356) );
  inv01 U5109 ( .Y(n6344), .A(n6363) );
  ao221 U5110 ( .Y(n6364), .A0(n7528), .A1(n7388), .B0(n7530), .B1(n7390), 
        .C0(n7669) );
  inv01 U5111 ( .Y(n6365), .A(n6364) );
  nand02 U5112 ( .Y(n7478), .A0(n6366), .A1(n6367) );
  inv02 U5113 ( .Y(n6368), .A(n7561) );
  inv01 U5114 ( .Y(n6369), .A(n7388) );
  inv01 U5115 ( .Y(n6370), .A(n7390) );
  inv01 U5116 ( .Y(n6371), .A(n7506) );
  inv01 U5117 ( .Y(n6372), .A(n7525) );
  nand02 U5118 ( .Y(n6373), .A0(n6370), .A1(n6374) );
  nand02 U5119 ( .Y(n6375), .A0(n6371), .A1(n6376) );
  nand02 U5120 ( .Y(n6377), .A0(n6372), .A1(n6378) );
  nand02 U5121 ( .Y(n6379), .A0(n6372), .A1(n6380) );
  nand02 U5122 ( .Y(n6381), .A0(n6368), .A1(n6369) );
  inv01 U5123 ( .Y(n6374), .A(n6381) );
  nand02 U5124 ( .Y(n6382), .A0(n6368), .A1(n6369) );
  inv01 U5125 ( .Y(n6376), .A(n6382) );
  nand02 U5126 ( .Y(n6383), .A0(n6368), .A1(n6370) );
  inv01 U5127 ( .Y(n6378), .A(n6383) );
  nand02 U5128 ( .Y(n6384), .A0(n6368), .A1(n6371) );
  inv01 U5129 ( .Y(n6380), .A(n6384) );
  nand02 U5130 ( .Y(n6385), .A0(n6373), .A1(n6375) );
  inv01 U5131 ( .Y(n6366), .A(n6385) );
  nand02 U5132 ( .Y(n6386), .A0(n6377), .A1(n6379) );
  inv01 U5133 ( .Y(n6367), .A(n6386) );
  nand02 U5134 ( .Y(n7469), .A0(n6387), .A1(n6388) );
  inv02 U5135 ( .Y(n6389), .A(n7557) );
  inv01 U5136 ( .Y(n6390), .A(n7388) );
  inv01 U5137 ( .Y(n6391), .A(n7390) );
  inv01 U5138 ( .Y(n6392), .A(n7500) );
  inv01 U5139 ( .Y(n6393), .A(n7521) );
  nand02 U5140 ( .Y(n6394), .A0(n6391), .A1(n6395) );
  nand02 U5141 ( .Y(n6396), .A0(n6392), .A1(n6397) );
  nand02 U5142 ( .Y(n6398), .A0(n6393), .A1(n6399) );
  nand02 U5143 ( .Y(n6400), .A0(n6393), .A1(n6401) );
  nand02 U5144 ( .Y(n6402), .A0(n6389), .A1(n6390) );
  inv01 U5145 ( .Y(n6395), .A(n6402) );
  nand02 U5146 ( .Y(n6403), .A0(n6389), .A1(n6390) );
  inv01 U5147 ( .Y(n6397), .A(n6403) );
  nand02 U5148 ( .Y(n6404), .A0(n6389), .A1(n6391) );
  inv01 U5149 ( .Y(n6399), .A(n6404) );
  nand02 U5150 ( .Y(n6405), .A0(n6389), .A1(n6392) );
  inv01 U5151 ( .Y(n6401), .A(n6405) );
  nand02 U5152 ( .Y(n6406), .A0(n6394), .A1(n6396) );
  inv01 U5153 ( .Y(n6387), .A(n6406) );
  nand02 U5154 ( .Y(n6407), .A0(n6398), .A1(n6400) );
  inv01 U5155 ( .Y(n6388), .A(n6407) );
  ao221 U5156 ( .Y(n6408), .A0(n7494), .A1(n7390), .B0(n7516), .B1(n7388), 
        .C0(n7553) );
  inv01 U5157 ( .Y(n6409), .A(n6408) );
  nand02 U5158 ( .Y(n7539), .A0(n6410), .A1(n6411) );
  inv02 U5159 ( .Y(n6412), .A(n7615) );
  inv01 U5160 ( .Y(n6413), .A(n7388) );
  inv01 U5161 ( .Y(n6414), .A(n7390) );
  inv01 U5162 ( .Y(n6415), .A(n7558) );
  inv01 U5163 ( .Y(n6416), .A(n7577) );
  nand02 U5164 ( .Y(n6417), .A0(n6414), .A1(n6418) );
  nand02 U5165 ( .Y(n6419), .A0(n6415), .A1(n6420) );
  nand02 U5166 ( .Y(n6421), .A0(n6416), .A1(n6422) );
  nand02 U5167 ( .Y(n6423), .A0(n6416), .A1(n6424) );
  nand02 U5168 ( .Y(n6425), .A0(n6412), .A1(n6413) );
  inv01 U5169 ( .Y(n6418), .A(n6425) );
  nand02 U5170 ( .Y(n6426), .A0(n6412), .A1(n6413) );
  inv01 U5171 ( .Y(n6420), .A(n6426) );
  nand02 U5172 ( .Y(n6427), .A0(n6412), .A1(n6414) );
  inv01 U5173 ( .Y(n6422), .A(n6427) );
  nand02 U5174 ( .Y(n6428), .A0(n6412), .A1(n6415) );
  inv01 U5175 ( .Y(n6424), .A(n6428) );
  nand02 U5176 ( .Y(n6429), .A0(n6417), .A1(n6419) );
  inv01 U5177 ( .Y(n6410), .A(n6429) );
  nand02 U5178 ( .Y(n6430), .A0(n6421), .A1(n6423) );
  inv01 U5179 ( .Y(n6411), .A(n6430) );
  nand02 U5180 ( .Y(n7444), .A0(n6431), .A1(n6432) );
  inv02 U5181 ( .Y(n6433), .A(n7546) );
  inv01 U5182 ( .Y(n6434), .A(n7388) );
  inv01 U5183 ( .Y(n6435), .A(n7390) );
  inv01 U5184 ( .Y(n6436), .A(n7481) );
  inv01 U5185 ( .Y(n6437), .A(n7506) );
  nand02 U5186 ( .Y(n6438), .A0(n6435), .A1(n6439) );
  nand02 U5187 ( .Y(n6440), .A0(n6436), .A1(n6441) );
  nand02 U5188 ( .Y(n6442), .A0(n6437), .A1(n6443) );
  nand02 U5189 ( .Y(n6444), .A0(n6437), .A1(n6445) );
  nand02 U5190 ( .Y(n6446), .A0(n6433), .A1(n6434) );
  inv01 U5191 ( .Y(n6439), .A(n6446) );
  nand02 U5192 ( .Y(n6447), .A0(n6433), .A1(n6434) );
  inv01 U5193 ( .Y(n6441), .A(n6447) );
  nand02 U5194 ( .Y(n6448), .A0(n6433), .A1(n6435) );
  inv01 U5195 ( .Y(n6443), .A(n6448) );
  nand02 U5196 ( .Y(n6449), .A0(n6433), .A1(n6436) );
  inv01 U5197 ( .Y(n6445), .A(n6449) );
  nand02 U5198 ( .Y(n6450), .A0(n6438), .A1(n6440) );
  inv01 U5199 ( .Y(n6431), .A(n6450) );
  nand02 U5200 ( .Y(n6451), .A0(n6442), .A1(n6444) );
  inv01 U5201 ( .Y(n6432), .A(n6451) );
  nand02 U5202 ( .Y(n7490), .A0(n6452), .A1(n6453) );
  inv02 U5203 ( .Y(n6454), .A(n7571) );
  inv01 U5204 ( .Y(n6455), .A(n7388) );
  inv01 U5205 ( .Y(n6456), .A(n7390) );
  inv01 U5206 ( .Y(n6457), .A(n7516) );
  inv01 U5207 ( .Y(n6458), .A(n7537) );
  nand02 U5208 ( .Y(n6459), .A0(n6456), .A1(n6460) );
  nand02 U5209 ( .Y(n6461), .A0(n6457), .A1(n6462) );
  nand02 U5210 ( .Y(n6463), .A0(n6458), .A1(n6464) );
  nand02 U5211 ( .Y(n6465), .A0(n6458), .A1(n6466) );
  nand02 U5212 ( .Y(n6467), .A0(n6454), .A1(n6455) );
  inv01 U5213 ( .Y(n6460), .A(n6467) );
  nand02 U5214 ( .Y(n6468), .A0(n6454), .A1(n6455) );
  inv01 U5215 ( .Y(n6462), .A(n6468) );
  nand02 U5216 ( .Y(n6469), .A0(n6454), .A1(n6456) );
  inv01 U5217 ( .Y(n6464), .A(n6469) );
  nand02 U5218 ( .Y(n6470), .A0(n6454), .A1(n6457) );
  inv01 U5219 ( .Y(n6466), .A(n6470) );
  nand02 U5220 ( .Y(n6471), .A0(n6459), .A1(n6461) );
  inv01 U5221 ( .Y(n6452), .A(n6471) );
  nand02 U5222 ( .Y(n6472), .A0(n6463), .A1(n6465) );
  inv01 U5223 ( .Y(n6453), .A(n6472) );
  nand02 U5224 ( .Y(n7518), .A0(n6473), .A1(n6474) );
  inv02 U5225 ( .Y(n6475), .A(n7596) );
  inv01 U5226 ( .Y(n6476), .A(n7388) );
  inv01 U5227 ( .Y(n6477), .A(n7390) );
  inv01 U5228 ( .Y(n6478), .A(n7543) );
  inv01 U5229 ( .Y(n6479), .A(n7558) );
  nand02 U5230 ( .Y(n6480), .A0(n6477), .A1(n6481) );
  nand02 U5231 ( .Y(n6482), .A0(n6478), .A1(n6483) );
  nand02 U5232 ( .Y(n6484), .A0(n6479), .A1(n6485) );
  nand02 U5233 ( .Y(n6486), .A0(n6479), .A1(n6487) );
  nand02 U5234 ( .Y(n6488), .A0(n6475), .A1(n6476) );
  inv01 U5235 ( .Y(n6481), .A(n6488) );
  nand02 U5236 ( .Y(n6489), .A0(n6475), .A1(n6476) );
  inv01 U5237 ( .Y(n6483), .A(n6489) );
  nand02 U5238 ( .Y(n6490), .A0(n6475), .A1(n6477) );
  inv01 U5239 ( .Y(n6485), .A(n6490) );
  nand02 U5240 ( .Y(n6491), .A0(n6475), .A1(n6478) );
  inv01 U5241 ( .Y(n6487), .A(n6491) );
  nand02 U5242 ( .Y(n6492), .A0(n6480), .A1(n6482) );
  inv01 U5243 ( .Y(n6473), .A(n6492) );
  nand02 U5244 ( .Y(n6493), .A0(n6484), .A1(n6486) );
  inv01 U5245 ( .Y(n6474), .A(n6493) );
  nor02 U5246 ( .Y(n6495), .A0(n7507), .A1(n7568) );
  nor02 U5247 ( .Y(n6496), .A0(n7566), .A1(n7567) );
  inv01 U5248 ( .Y(n6497), .A(n3329) );
  nor02 U5249 ( .Y(n6494), .A0(n6497), .A1(n6498) );
  nor02 U5250 ( .Y(n6499), .A0(n6495), .A1(n6496) );
  inv01 U5251 ( .Y(n6498), .A(n6499) );
  ao221 U5252 ( .Y(n6500), .A0(n7562), .A1(n7390), .B0(n7581), .B1(n7388), 
        .C0(n7619) );
  inv01 U5253 ( .Y(n6501), .A(n6500) );
  ao221 U5254 ( .Y(n6502), .A0(n7597), .A1(n7388), .B0(n7601), .B1(n7384), 
        .C0(n7628) );
  inv01 U5255 ( .Y(n6503), .A(n6502) );
  nand02 U5256 ( .Y(n7552), .A0(n6504), .A1(n6505) );
  inv02 U5257 ( .Y(n6506), .A(n7624) );
  inv01 U5258 ( .Y(n6507), .A(n7388) );
  inv01 U5259 ( .Y(n6508), .A(n7384) );
  inv01 U5260 ( .Y(n6509), .A(n7595) );
  inv01 U5261 ( .Y(n6510), .A(n7589) );
  nand02 U5262 ( .Y(n6511), .A0(n6508), .A1(n6512) );
  nand02 U5263 ( .Y(n6513), .A0(n6509), .A1(n6514) );
  nand02 U5264 ( .Y(n6515), .A0(n6510), .A1(n6516) );
  nand02 U5265 ( .Y(n6517), .A0(n6510), .A1(n6518) );
  nand02 U5266 ( .Y(n6519), .A0(n6506), .A1(n6507) );
  inv01 U5267 ( .Y(n6512), .A(n6519) );
  nand02 U5268 ( .Y(n6520), .A0(n6506), .A1(n6507) );
  inv01 U5269 ( .Y(n6514), .A(n6520) );
  nand02 U5270 ( .Y(n6521), .A0(n6506), .A1(n6508) );
  inv01 U5271 ( .Y(n6516), .A(n6521) );
  nand02 U5272 ( .Y(n6522), .A0(n6506), .A1(n6509) );
  inv01 U5273 ( .Y(n6518), .A(n6522) );
  nand02 U5274 ( .Y(n6523), .A0(n6511), .A1(n6513) );
  inv01 U5275 ( .Y(n6504), .A(n6523) );
  nand02 U5276 ( .Y(n6524), .A0(n6515), .A1(n6517) );
  inv01 U5277 ( .Y(n6505), .A(n6524) );
  inv01 U5278 ( .Y(n7509), .A(n6525) );
  nor02 U5279 ( .Y(n6526), .A0(n7566), .A1(n7568) );
  nor02 U5280 ( .Y(n6527), .A0(n7586), .A1(n7567) );
  inv01 U5281 ( .Y(n6528), .A(n3335) );
  nor02 U5282 ( .Y(n6525), .A0(n6528), .A1(n6529) );
  nor02 U5283 ( .Y(n6530), .A0(n6526), .A1(n6527) );
  inv01 U5284 ( .Y(n6529), .A(n6530) );
  nand02 U5285 ( .Y(n7551), .A0(n6531), .A1(n6532) );
  inv02 U5286 ( .Y(n6533), .A(n7622) );
  inv01 U5287 ( .Y(n6534), .A(n7388) );
  inv01 U5288 ( .Y(n6535), .A(n7390) );
  inv01 U5289 ( .Y(n6536), .A(n7569) );
  inv01 U5290 ( .Y(n6537), .A(n7587) );
  nand02 U5291 ( .Y(n6538), .A0(n6535), .A1(n6539) );
  nand02 U5292 ( .Y(n6540), .A0(n6536), .A1(n6541) );
  nand02 U5293 ( .Y(n6542), .A0(n6537), .A1(n6543) );
  nand02 U5294 ( .Y(n6544), .A0(n6537), .A1(n6545) );
  nand02 U5295 ( .Y(n6546), .A0(n6533), .A1(n6534) );
  inv01 U5296 ( .Y(n6539), .A(n6546) );
  nand02 U5297 ( .Y(n6547), .A0(n6533), .A1(n6534) );
  inv01 U5298 ( .Y(n6541), .A(n6547) );
  nand02 U5299 ( .Y(n6548), .A0(n6533), .A1(n6535) );
  inv01 U5300 ( .Y(n6543), .A(n6548) );
  nand02 U5301 ( .Y(n6549), .A0(n6533), .A1(n6536) );
  inv01 U5302 ( .Y(n6545), .A(n6549) );
  nand02 U5303 ( .Y(n6550), .A0(n6538), .A1(n6540) );
  inv01 U5304 ( .Y(n6531), .A(n6550) );
  nand02 U5305 ( .Y(n6551), .A0(n6542), .A1(n6544) );
  inv01 U5306 ( .Y(n6532), .A(n6551) );
  inv02 U5307 ( .Y(n7567), .A(n7388) );
  nand02 U5308 ( .Y(n7532), .A0(n6552), .A1(n6553) );
  inv02 U5309 ( .Y(n6554), .A(n7611) );
  inv01 U5310 ( .Y(n6555), .A(n7388) );
  inv01 U5311 ( .Y(n6556), .A(n7390) );
  inv01 U5312 ( .Y(n6557), .A(n7554) );
  inv01 U5313 ( .Y(n6558), .A(n7572) );
  nand02 U5314 ( .Y(n6559), .A0(n6556), .A1(n6560) );
  nand02 U5315 ( .Y(n6561), .A0(n6557), .A1(n6562) );
  nand02 U5316 ( .Y(n6563), .A0(n6558), .A1(n6564) );
  nand02 U5317 ( .Y(n6565), .A0(n6558), .A1(n6566) );
  nand02 U5318 ( .Y(n6567), .A0(n6554), .A1(n6555) );
  inv01 U5319 ( .Y(n6560), .A(n6567) );
  nand02 U5320 ( .Y(n6568), .A0(n6554), .A1(n6555) );
  inv01 U5321 ( .Y(n6562), .A(n6568) );
  nand02 U5322 ( .Y(n6569), .A0(n6554), .A1(n6556) );
  inv01 U5323 ( .Y(n6564), .A(n6569) );
  nand02 U5324 ( .Y(n6570), .A0(n6554), .A1(n6557) );
  inv01 U5325 ( .Y(n6566), .A(n6570) );
  nand02 U5326 ( .Y(n6571), .A0(n6559), .A1(n6561) );
  inv01 U5327 ( .Y(n6552), .A(n6571) );
  nand02 U5328 ( .Y(n6572), .A0(n6563), .A1(n6565) );
  inv01 U5329 ( .Y(n6553), .A(n6572) );
  ao221 U5330 ( .Y(n6573), .A0(n7549), .A1(n7390), .B0(n7562), .B1(n7388), 
        .C0(n7605) );
  inv01 U5331 ( .Y(n6574), .A(n6573) );
  inv02 U5332 ( .Y(n6576), .A(n6575) );
  inv01 U5333 ( .Y(n7526), .A(n6577) );
  nor02 U5334 ( .Y(n6578), .A0(n7395), .A1(n7582) );
  nor02 U5335 ( .Y(n6579), .A0(n7404), .A1(n7591) );
  inv01 U5336 ( .Y(n6580), .A(n7670) );
  nor02 U5337 ( .Y(n6577), .A0(n6580), .A1(n6581) );
  nor02 U5338 ( .Y(n6582), .A0(n6578), .A1(n6579) );
  inv01 U5339 ( .Y(n6581), .A(n6582) );
  inv02 U5340 ( .Y(n7674), .A(c_0_) );
  nor02 U5341 ( .Y(n6584), .A0(n7395), .A1(n7480) );
  nor02 U5342 ( .Y(n6585), .A0(n7404), .A1(n7493) );
  inv01 U5343 ( .Y(n6586), .A(n7668) );
  nor02 U5344 ( .Y(n6583), .A0(n6586), .A1(n6587) );
  nor02 U5345 ( .Y(n6588), .A0(n6584), .A1(n6585) );
  inv01 U5346 ( .Y(n6587), .A(n6588) );
  nor02 U5347 ( .Y(n6590), .A0(n7394), .A1(n7492) );
  nor02 U5348 ( .Y(n6591), .A0(n7403), .A1(n7498) );
  inv01 U5349 ( .Y(n6592), .A(n7499) );
  nor02 U5350 ( .Y(n6589), .A0(n6592), .A1(n6593) );
  nor02 U5351 ( .Y(n6594), .A0(n6590), .A1(n6591) );
  inv01 U5352 ( .Y(n6593), .A(n6594) );
  nor02 U5353 ( .Y(n6596), .A0(n7393), .A1(n7474) );
  nor02 U5354 ( .Y(n6597), .A0(n7403), .A1(n7480) );
  inv01 U5355 ( .Y(n6598), .A(n3557) );
  nor02 U5356 ( .Y(n6595), .A0(n6598), .A1(n6599) );
  nor02 U5357 ( .Y(n6600), .A0(n6596), .A1(n6597) );
  inv01 U5358 ( .Y(n6599), .A(n6600) );
  nor02 U5359 ( .Y(n6602), .A0(n7395), .A1(n7493) );
  nor02 U5360 ( .Y(n6603), .A0(n7403), .A1(n7492) );
  inv01 U5361 ( .Y(n6604), .A(n3463) );
  nor02 U5362 ( .Y(n6601), .A0(n6604), .A1(n6605) );
  nor02 U5363 ( .Y(n6606), .A0(n6602), .A1(n6603) );
  inv01 U5364 ( .Y(n6605), .A(n6606) );
  inv02 U5365 ( .Y(n7493), .A(r0_43_) );
  inv02 U5366 ( .Y(n7480), .A(r0_44_) );
  inv02 U5367 ( .Y(n7492), .A(r0_42_) );
  inv02 U5368 ( .Y(n7474), .A(r0_45_) );
  inv01 U5369 ( .Y(n7530), .A(n6607) );
  nor02 U5370 ( .Y(n6608), .A0(n7393), .A1(n7550) );
  nor02 U5371 ( .Y(n6609), .A0(n7403), .A1(n7556) );
  inv01 U5372 ( .Y(n6610), .A(n7672) );
  nor02 U5373 ( .Y(n6607), .A0(n6610), .A1(n6611) );
  nor02 U5374 ( .Y(n6612), .A0(n6608), .A1(n6609) );
  inv01 U5375 ( .Y(n6611), .A(n6612) );
  inv02 U5376 ( .Y(n7568), .A(n7390) );
  nand02 U5377 ( .Y(n7584), .A0(n6613), .A1(n6614) );
  inv02 U5378 ( .Y(n6615), .A(n7390) );
  inv02 U5379 ( .Y(n6616), .A(n7384) );
  inv02 U5380 ( .Y(n6617), .A(n7388) );
  inv02 U5381 ( .Y(n6618), .A(n7608) );
  inv02 U5382 ( .Y(n6619), .A(n7635) );
  inv02 U5383 ( .Y(n6620), .A(n7609) );
  nand02 U5384 ( .Y(n6621), .A0(n6617), .A1(n6622) );
  nand02 U5385 ( .Y(n6623), .A0(n6618), .A1(n6624) );
  nand02 U5386 ( .Y(n6625), .A0(n6619), .A1(n6626) );
  nand02 U5387 ( .Y(n6627), .A0(n6619), .A1(n6628) );
  nand02 U5388 ( .Y(n6629), .A0(n6620), .A1(n6630) );
  nand02 U5389 ( .Y(n6631), .A0(n6620), .A1(n6632) );
  nand02 U5390 ( .Y(n6633), .A0(n6620), .A1(n6634) );
  nand02 U5391 ( .Y(n6635), .A0(n6620), .A1(n6636) );
  nand02 U5392 ( .Y(n6637), .A0(n6615), .A1(n6616) );
  inv01 U5393 ( .Y(n6622), .A(n6637) );
  nand02 U5394 ( .Y(n6638), .A0(n6615), .A1(n6616) );
  inv01 U5395 ( .Y(n6624), .A(n6638) );
  nand02 U5396 ( .Y(n6639), .A0(n6615), .A1(n6617) );
  inv01 U5397 ( .Y(n6626), .A(n6639) );
  nand02 U5398 ( .Y(n6640), .A0(n6615), .A1(n6618) );
  inv01 U5399 ( .Y(n6628), .A(n6640) );
  nand02 U5400 ( .Y(n6641), .A0(n6616), .A1(n6617) );
  inv01 U5401 ( .Y(n6630), .A(n6641) );
  nand02 U5402 ( .Y(n6642), .A0(n6616), .A1(n6618) );
  inv01 U5403 ( .Y(n6632), .A(n6642) );
  nand02 U5404 ( .Y(n6643), .A0(n6617), .A1(n6619) );
  inv01 U5405 ( .Y(n6634), .A(n6643) );
  nand02 U5406 ( .Y(n6644), .A0(n6618), .A1(n6619) );
  inv01 U5407 ( .Y(n6636), .A(n6644) );
  nand02 U5408 ( .Y(n6645), .A0(n6621), .A1(n6623) );
  inv01 U5409 ( .Y(n6646), .A(n6645) );
  nand02 U5410 ( .Y(n6647), .A0(n6625), .A1(n6627) );
  inv01 U5411 ( .Y(n6648), .A(n6647) );
  nand02 U5412 ( .Y(n6649), .A0(n6646), .A1(n6648) );
  inv01 U5413 ( .Y(n6613), .A(n6649) );
  nand02 U5414 ( .Y(n6650), .A0(n6629), .A1(n6631) );
  inv01 U5415 ( .Y(n6651), .A(n6650) );
  nand02 U5416 ( .Y(n6652), .A0(n6633), .A1(n6635) );
  inv01 U5417 ( .Y(n6653), .A(n6652) );
  nand02 U5418 ( .Y(n6654), .A0(n6651), .A1(n6653) );
  inv01 U5419 ( .Y(n6614), .A(n6654) );
  nand02 U5420 ( .Y(n7435), .A0(n6655), .A1(n6656) );
  inv02 U5421 ( .Y(n6657), .A(n7390) );
  inv02 U5422 ( .Y(n6658), .A(n7600) );
  inv02 U5423 ( .Y(n6659), .A(n7388) );
  inv02 U5424 ( .Y(n6660), .A(n7599) );
  inv02 U5425 ( .Y(n6661), .A(n7384) );
  inv02 U5426 ( .Y(n6662), .A(n7601) );
  nand02 U5427 ( .Y(n6663), .A0(n6659), .A1(n6664) );
  nand02 U5428 ( .Y(n6665), .A0(n6660), .A1(n6666) );
  nand02 U5429 ( .Y(n6667), .A0(n6661), .A1(n6668) );
  nand02 U5430 ( .Y(n6669), .A0(n6661), .A1(n6670) );
  nand02 U5431 ( .Y(n6671), .A0(n6662), .A1(n6672) );
  nand02 U5432 ( .Y(n6673), .A0(n6662), .A1(n6674) );
  nand02 U5433 ( .Y(n6675), .A0(n6662), .A1(n6676) );
  nand02 U5434 ( .Y(n6677), .A0(n6662), .A1(n6678) );
  nand02 U5435 ( .Y(n6679), .A0(n6657), .A1(n6658) );
  inv01 U5436 ( .Y(n6664), .A(n6679) );
  nand02 U5437 ( .Y(n6680), .A0(n6657), .A1(n6658) );
  inv01 U5438 ( .Y(n6666), .A(n6680) );
  nand02 U5439 ( .Y(n6681), .A0(n6657), .A1(n6659) );
  inv01 U5440 ( .Y(n6668), .A(n6681) );
  nand02 U5441 ( .Y(n6682), .A0(n6657), .A1(n6660) );
  inv01 U5442 ( .Y(n6670), .A(n6682) );
  nand02 U5443 ( .Y(n6683), .A0(n6658), .A1(n6659) );
  inv01 U5444 ( .Y(n6672), .A(n6683) );
  nand02 U5445 ( .Y(n6684), .A0(n6658), .A1(n6660) );
  inv01 U5446 ( .Y(n6674), .A(n6684) );
  nand02 U5447 ( .Y(n6685), .A0(n6659), .A1(n6661) );
  inv01 U5448 ( .Y(n6676), .A(n6685) );
  nand02 U5449 ( .Y(n6686), .A0(n6660), .A1(n6661) );
  inv01 U5450 ( .Y(n6678), .A(n6686) );
  nand02 U5451 ( .Y(n6687), .A0(n6663), .A1(n6665) );
  inv01 U5452 ( .Y(n6688), .A(n6687) );
  nand02 U5453 ( .Y(n6689), .A0(n6667), .A1(n6669) );
  inv01 U5454 ( .Y(n6690), .A(n6689) );
  nand02 U5455 ( .Y(n6691), .A0(n6688), .A1(n6690) );
  inv01 U5456 ( .Y(n6655), .A(n6691) );
  nand02 U5457 ( .Y(n6692), .A0(n6671), .A1(n6673) );
  inv01 U5458 ( .Y(n6693), .A(n6692) );
  nand02 U5459 ( .Y(n6694), .A0(n6675), .A1(n6677) );
  inv01 U5460 ( .Y(n6695), .A(n6694) );
  nand02 U5461 ( .Y(n6696), .A0(n6693), .A1(n6695) );
  inv01 U5462 ( .Y(n6656), .A(n6696) );
  nand02 U5463 ( .Y(n7434), .A0(n6697), .A1(n6698) );
  inv02 U5464 ( .Y(n6699), .A(n7390) );
  inv02 U5465 ( .Y(n6700), .A(n7384) );
  inv02 U5466 ( .Y(n6701), .A(n7388) );
  inv02 U5467 ( .Y(n6702), .A(n7593) );
  inv02 U5468 ( .Y(n6703), .A(n7594) );
  inv02 U5469 ( .Y(n6704), .A(n7595) );
  nand02 U5470 ( .Y(n6705), .A0(n6701), .A1(n6706) );
  nand02 U5471 ( .Y(n6707), .A0(n6702), .A1(n6708) );
  nand02 U5472 ( .Y(n6709), .A0(n6703), .A1(n6710) );
  nand02 U5473 ( .Y(n6711), .A0(n6703), .A1(n6712) );
  nand02 U5474 ( .Y(n6713), .A0(n6704), .A1(n6714) );
  nand02 U5475 ( .Y(n6715), .A0(n6704), .A1(n6716) );
  nand02 U5476 ( .Y(n6717), .A0(n6704), .A1(n6718) );
  nand02 U5477 ( .Y(n6719), .A0(n6704), .A1(n6720) );
  nand02 U5478 ( .Y(n6721), .A0(n6699), .A1(n6700) );
  inv01 U5479 ( .Y(n6706), .A(n6721) );
  nand02 U5480 ( .Y(n6722), .A0(n6699), .A1(n6700) );
  inv01 U5481 ( .Y(n6708), .A(n6722) );
  nand02 U5482 ( .Y(n6723), .A0(n6699), .A1(n6701) );
  inv01 U5483 ( .Y(n6710), .A(n6723) );
  nand02 U5484 ( .Y(n6724), .A0(n6699), .A1(n6702) );
  inv01 U5485 ( .Y(n6712), .A(n6724) );
  nand02 U5486 ( .Y(n6725), .A0(n6700), .A1(n6701) );
  inv01 U5487 ( .Y(n6714), .A(n6725) );
  nand02 U5488 ( .Y(n6726), .A0(n6700), .A1(n6702) );
  inv01 U5489 ( .Y(n6716), .A(n6726) );
  nand02 U5490 ( .Y(n6727), .A0(n6701), .A1(n6703) );
  inv01 U5491 ( .Y(n6718), .A(n6727) );
  nand02 U5492 ( .Y(n6728), .A0(n6702), .A1(n6703) );
  inv01 U5493 ( .Y(n6720), .A(n6728) );
  nand02 U5494 ( .Y(n6729), .A0(n6705), .A1(n6707) );
  inv01 U5495 ( .Y(n6730), .A(n6729) );
  nand02 U5496 ( .Y(n6731), .A0(n6709), .A1(n6711) );
  inv01 U5497 ( .Y(n6732), .A(n6731) );
  nand02 U5498 ( .Y(n6733), .A0(n6730), .A1(n6732) );
  inv01 U5499 ( .Y(n6697), .A(n6733) );
  nand02 U5500 ( .Y(n6734), .A0(n6713), .A1(n6715) );
  inv01 U5501 ( .Y(n6735), .A(n6734) );
  nand02 U5502 ( .Y(n6736), .A0(n6717), .A1(n6719) );
  inv01 U5503 ( .Y(n6737), .A(n6736) );
  nand02 U5504 ( .Y(n6738), .A0(n6735), .A1(n6737) );
  inv01 U5505 ( .Y(n6698), .A(n6738) );
  nand02 U5506 ( .Y(n7575), .A0(n6739), .A1(n6740) );
  inv02 U5507 ( .Y(n6741), .A(n7388) );
  inv02 U5508 ( .Y(n6742), .A(c_3_) );
  inv02 U5509 ( .Y(n6743), .A(n7390) );
  inv02 U5510 ( .Y(n6744), .A(n7597) );
  inv02 U5511 ( .Y(n6745), .A(n7617) );
  inv02 U5512 ( .Y(n6746), .A(n7601) );
  nand02 U5513 ( .Y(n6747), .A0(n6743), .A1(n6748) );
  nand02 U5514 ( .Y(n6749), .A0(n6744), .A1(n6750) );
  nand02 U5515 ( .Y(n6751), .A0(n6745), .A1(n6752) );
  nand02 U5516 ( .Y(n6753), .A0(n6745), .A1(n6754) );
  nand02 U5517 ( .Y(n6755), .A0(n6746), .A1(n6756) );
  nand02 U5518 ( .Y(n6757), .A0(n6746), .A1(n6758) );
  nand02 U5519 ( .Y(n6759), .A0(n6746), .A1(n6760) );
  nand02 U5520 ( .Y(n6761), .A0(n6746), .A1(n6762) );
  nand02 U5521 ( .Y(n6763), .A0(n6741), .A1(n6742) );
  inv01 U5522 ( .Y(n6748), .A(n6763) );
  nand02 U5523 ( .Y(n6764), .A0(n6741), .A1(n6742) );
  inv01 U5524 ( .Y(n6750), .A(n6764) );
  nand02 U5525 ( .Y(n6765), .A0(n6741), .A1(n6743) );
  inv01 U5526 ( .Y(n6752), .A(n6765) );
  nand02 U5527 ( .Y(n6766), .A0(n6741), .A1(n6744) );
  inv01 U5528 ( .Y(n6754), .A(n6766) );
  nand02 U5529 ( .Y(n6767), .A0(n6742), .A1(n6743) );
  inv01 U5530 ( .Y(n6756), .A(n6767) );
  nand02 U5531 ( .Y(n6768), .A0(n6742), .A1(n6744) );
  inv01 U5532 ( .Y(n6758), .A(n6768) );
  nand02 U5533 ( .Y(n6769), .A0(n6743), .A1(n6745) );
  inv01 U5534 ( .Y(n6760), .A(n6769) );
  nand02 U5535 ( .Y(n6770), .A0(n6744), .A1(n6745) );
  inv01 U5536 ( .Y(n6762), .A(n6770) );
  nand02 U5537 ( .Y(n6771), .A0(n6747), .A1(n6749) );
  inv01 U5538 ( .Y(n6772), .A(n6771) );
  nand02 U5539 ( .Y(n6773), .A0(n6751), .A1(n6753) );
  inv01 U5540 ( .Y(n6774), .A(n6773) );
  nand02 U5541 ( .Y(n6775), .A0(n6772), .A1(n6774) );
  inv01 U5542 ( .Y(n6739), .A(n6775) );
  nand02 U5543 ( .Y(n6776), .A0(n6755), .A1(n6757) );
  inv01 U5544 ( .Y(n6777), .A(n6776) );
  nand02 U5545 ( .Y(n6778), .A0(n6759), .A1(n6761) );
  inv01 U5546 ( .Y(n6779), .A(n6778) );
  nand02 U5547 ( .Y(n6780), .A0(n6777), .A1(n6779) );
  inv01 U5548 ( .Y(n6740), .A(n6780) );
  buf02 U5549 ( .Y(n6781), .A(s_rad_i_51_) );
  buf02 U5550 ( .Y(n6783), .A(s_rad_i_51_) );
  buf02 U5551 ( .Y(n6782), .A(s_rad_i_51_) );
  nand02 U5552 ( .Y(n7579), .A0(n6784), .A1(n6785) );
  inv02 U5553 ( .Y(n6786), .A(n7390) );
  inv02 U5554 ( .Y(n6787), .A(n7384) );
  inv02 U5555 ( .Y(n6788), .A(n7388) );
  inv02 U5556 ( .Y(n6789), .A(n7604) );
  inv02 U5557 ( .Y(n6790), .A(n7621) );
  inv02 U5558 ( .Y(n6791), .A(n7606) );
  nand02 U5559 ( .Y(n6792), .A0(n6788), .A1(n6793) );
  nand02 U5560 ( .Y(n6794), .A0(n6789), .A1(n6795) );
  nand02 U5561 ( .Y(n6796), .A0(n6790), .A1(n6797) );
  nand02 U5562 ( .Y(n6798), .A0(n6790), .A1(n6799) );
  nand02 U5563 ( .Y(n6800), .A0(n6791), .A1(n6801) );
  nand02 U5564 ( .Y(n6802), .A0(n6791), .A1(n6803) );
  nand02 U5565 ( .Y(n6804), .A0(n6791), .A1(n6805) );
  nand02 U5566 ( .Y(n6806), .A0(n6791), .A1(n6807) );
  nand02 U5567 ( .Y(n6808), .A0(n6786), .A1(n6787) );
  inv01 U5568 ( .Y(n6793), .A(n6808) );
  nand02 U5569 ( .Y(n6809), .A0(n6786), .A1(n6787) );
  inv01 U5570 ( .Y(n6795), .A(n6809) );
  nand02 U5571 ( .Y(n6810), .A0(n6786), .A1(n6788) );
  inv01 U5572 ( .Y(n6797), .A(n6810) );
  nand02 U5573 ( .Y(n6811), .A0(n6786), .A1(n6789) );
  inv01 U5574 ( .Y(n6799), .A(n6811) );
  nand02 U5575 ( .Y(n6812), .A0(n6787), .A1(n6788) );
  inv01 U5576 ( .Y(n6801), .A(n6812) );
  nand02 U5577 ( .Y(n6813), .A0(n6787), .A1(n6789) );
  inv01 U5578 ( .Y(n6803), .A(n6813) );
  nand02 U5579 ( .Y(n6814), .A0(n6788), .A1(n6790) );
  inv01 U5580 ( .Y(n6805), .A(n6814) );
  nand02 U5581 ( .Y(n6815), .A0(n6789), .A1(n6790) );
  inv01 U5582 ( .Y(n6807), .A(n6815) );
  nand02 U5583 ( .Y(n6816), .A0(n6792), .A1(n6794) );
  inv01 U5584 ( .Y(n6817), .A(n6816) );
  nand02 U5585 ( .Y(n6818), .A0(n6796), .A1(n6798) );
  inv01 U5586 ( .Y(n6819), .A(n6818) );
  nand02 U5587 ( .Y(n6820), .A0(n6817), .A1(n6819) );
  inv01 U5588 ( .Y(n6784), .A(n6820) );
  nand02 U5589 ( .Y(n6821), .A0(n6800), .A1(n6802) );
  inv01 U5590 ( .Y(n6822), .A(n6821) );
  nand02 U5591 ( .Y(n6823), .A0(n6804), .A1(n6806) );
  inv01 U5592 ( .Y(n6824), .A(n6823) );
  nand02 U5593 ( .Y(n6825), .A0(n6822), .A1(n6824) );
  inv01 U5594 ( .Y(n6785), .A(n6825) );
  ao21 U5595 ( .Y(n6826), .A0(n6950), .A1(n7676), .B0(n7419) );
  inv02 U5596 ( .Y(n6827), .A(n6826) );
  ao221 U5597 ( .Y(n6828), .A0(n7609), .A1(n7374), .B0(n7570), .B1(n7390), 
        .C0(n7610) );
  inv02 U5598 ( .Y(n6829), .A(n6828) );
  inv02 U5599 ( .Y(n7566), .A(n7526) );
  inv02 U5600 ( .Y(n7570), .A(n6856) );
  nor02 U5601 ( .Y(n6857), .A0(n7394), .A1(n7607) );
  nor02 U5602 ( .Y(n6858), .A0(n7404), .A1(n7613) );
  inv01 U5603 ( .Y(n6859), .A(n7671) );
  nor02 U5604 ( .Y(n6856), .A0(n6859), .A1(n6860) );
  nor02 U5605 ( .Y(n6861), .A0(n6857), .A1(n6858) );
  inv01 U5606 ( .Y(n6860), .A(n6861) );
  inv02 U5607 ( .Y(n7586), .A(n7570) );
  inv02 U5608 ( .Y(n7599), .A(n6862) );
  nor02 U5609 ( .Y(n6863), .A0(n7641), .A1(n7393) );
  nor02 U5610 ( .Y(n6864), .A0(n7652), .A1(n7404) );
  inv01 U5611 ( .Y(n6865), .A(n7653) );
  nor02 U5612 ( .Y(n6862), .A0(n6865), .A1(n6866) );
  nor02 U5613 ( .Y(n6867), .A0(n6863), .A1(n6864) );
  inv01 U5614 ( .Y(n6866), .A(n6867) );
  inv02 U5615 ( .Y(n7486), .A(n6894) );
  nor02 U5616 ( .Y(n6895), .A0(n7394), .A1(n7504) );
  nor02 U5617 ( .Y(n6896), .A0(n7403), .A1(n7515) );
  inv01 U5618 ( .Y(n6897), .A(n3794) );
  nor02 U5619 ( .Y(n6894), .A0(n6897), .A1(n6898) );
  nor02 U5620 ( .Y(n6899), .A0(n6895), .A1(n6896) );
  inv01 U5621 ( .Y(n6898), .A(n6899) );
  inv02 U5622 ( .Y(n7528), .A(n6900) );
  nor02 U5623 ( .Y(n6901), .A0(n7395), .A1(n7563) );
  nor02 U5624 ( .Y(n6902), .A0(n7403), .A1(n7574) );
  inv01 U5625 ( .Y(n6903), .A(n7673) );
  nor02 U5626 ( .Y(n6900), .A0(n6903), .A1(n6904) );
  nor02 U5627 ( .Y(n6905), .A0(n6901), .A1(n6902) );
  inv01 U5628 ( .Y(n6904), .A(n6905) );
  inv04 U5629 ( .Y(n7658), .A(r0_0_) );
  inv02 U5630 ( .Y(n7621), .A(n6907) );
  nor02 U5631 ( .Y(n6908), .A0(n7652), .A1(n7395) );
  nor02 U5632 ( .Y(n6909), .A0(n7658), .A1(n7404) );
  inv01 U5633 ( .Y(n6910), .A(n7659) );
  nor02 U5634 ( .Y(n6907), .A0(n6910), .A1(n6911) );
  nor02 U5635 ( .Y(n6912), .A0(n6908), .A1(n6909) );
  inv01 U5636 ( .Y(n6911), .A(n6912) );
  inv02 U5637 ( .Y(n7471), .A(n6913) );
  nor02 U5638 ( .Y(n6914), .A0(n7394), .A1(n7514) );
  nor02 U5639 ( .Y(n6915), .A0(n7404), .A1(n7520) );
  inv01 U5640 ( .Y(n6916), .A(n3756) );
  nor02 U5641 ( .Y(n6913), .A0(n6916), .A1(n6917) );
  nor02 U5642 ( .Y(n6918), .A0(n6914), .A1(n6915) );
  inv01 U5643 ( .Y(n6917), .A(n6918) );
  inv02 U5644 ( .Y(n7461), .A(n6919) );
  nor02 U5645 ( .Y(n6920), .A0(n7395), .A1(n7515) );
  nor02 U5646 ( .Y(n6921), .A0(n7404), .A1(n7514) );
  inv01 U5647 ( .Y(n6922), .A(n3637) );
  nor02 U5648 ( .Y(n6919), .A0(n6922), .A1(n6923) );
  nor02 U5649 ( .Y(n6924), .A0(n6920), .A1(n6921) );
  inv01 U5650 ( .Y(n6923), .A(n6924) );
  inv02 U5651 ( .Y(n7593), .A(n6925) );
  nor02 U5652 ( .Y(n6926), .A0(n7393), .A1(n7642) );
  nor02 U5653 ( .Y(n6927), .A0(n7404), .A1(n7641) );
  inv01 U5654 ( .Y(n6928), .A(n7643) );
  nor02 U5655 ( .Y(n6925), .A0(n6928), .A1(n6929) );
  nor02 U5656 ( .Y(n6930), .A0(n6926), .A1(n6927) );
  inv01 U5657 ( .Y(n6929), .A(n6930) );
  inv02 U5658 ( .Y(n7514), .A(r0_38_) );
  inv02 U5659 ( .Y(n7515), .A(r0_39_) );
  inv02 U5660 ( .Y(n7447), .A(n6931) );
  nor02 U5661 ( .Y(n6932), .A0(n7393), .A1(n7498) );
  nor02 U5662 ( .Y(n6933), .A0(n7403), .A1(n7504) );
  inv01 U5663 ( .Y(n6934), .A(n7505) );
  nor02 U5664 ( .Y(n6931), .A0(n6934), .A1(n6935) );
  nor02 U5665 ( .Y(n6936), .A0(n6932), .A1(n6933) );
  inv01 U5666 ( .Y(n6935), .A(n6936) );
  inv02 U5667 ( .Y(n7504), .A(r0_40_) );
  inv02 U5668 ( .Y(n7498), .A(r0_41_) );
  inv02 U5669 ( .Y(n7510), .A(n6937) );
  nor02 U5670 ( .Y(n6938), .A0(n7393), .A1(n7524) );
  nor02 U5671 ( .Y(n6939), .A0(n7404), .A1(n7535) );
  inv01 U5672 ( .Y(n6940), .A(n3663) );
  nor02 U5673 ( .Y(n6937), .A0(n6940), .A1(n6941) );
  nor02 U5674 ( .Y(n6942), .A0(n6938), .A1(n6939) );
  inv01 U5675 ( .Y(n6941), .A(n6942) );
  inv04 U5676 ( .Y(n6943), .A(c_1_) );
  inv02 U5677 ( .Y(n6944), .A(n6943) );
  inv08 U5678 ( .Y(n6946), .A(n6943) );
  inv02 U5679 ( .Y(n6945), .A(n6943) );
  inv04 U5680 ( .Y(n6948), .A(n6947) );
  inv02 U5681 ( .Y(n6950), .A(n6949) );
  or02 U5682 ( .Y(n6951), .A0(n7421), .A1(n7676) );
  inv02 U5683 ( .Y(n6952), .A(n6951) );
  inv01 U5684 ( .Y(n6953), .A(s_op2_6_) );
  inv01 U5685 ( .Y(n6954), .A(n6953) );
  inv02 U5686 ( .Y(n6955), .A(n6953) );
  inv02 U5687 ( .Y(s_op2_7_), .A(n6956) );
  nor02 U5688 ( .Y(n6957), .A0(n7438), .A1(n7439) );
  nor02 U5689 ( .Y(n6958), .A0(n7436), .A1(n7437) );
  nor02 U5690 ( .Y(n6956), .A0(n6957), .A1(n6958) );
  inv01 U5691 ( .Y(n6959), .A(s_op2_5_) );
  inv01 U5692 ( .Y(n6960), .A(n6959) );
  inv02 U5693 ( .Y(n6961), .A(n6959) );
  inv02 U5694 ( .Y(s_op2_18_), .A(n6962) );
  nor02 U5695 ( .Y(n6963), .A0(n7378), .A1(n7551) );
  nor02 U5696 ( .Y(n6964), .A0(n7364), .A1(n7367) );
  nor02 U5697 ( .Y(n6962), .A0(n6963), .A1(n6964) );
  inv02 U5698 ( .Y(s_op2_16_), .A(n6965) );
  nor02 U5699 ( .Y(n6966), .A0(n7627), .A1(n7367) );
  nor02 U5700 ( .Y(n6967), .A0(n7378), .A1(n6503) );
  nor02 U5701 ( .Y(n6965), .A0(n6966), .A1(n6967) );
  inv02 U5702 ( .Y(n7378), .A(n7376) );
  inv02 U5703 ( .Y(s_op2_19_), .A(n6968) );
  nor02 U5704 ( .Y(n6969), .A0(n7378), .A1(n6501) );
  nor02 U5705 ( .Y(n6970), .A0(n7438), .A1(n7367) );
  nor02 U5706 ( .Y(n6968), .A0(n6969), .A1(n6970) );
  inv02 U5707 ( .Y(s_op2_17_), .A(n6971) );
  nor02 U5708 ( .Y(n6972), .A0(n7378), .A1(n7552) );
  nor02 U5709 ( .Y(n6973), .A0(n7366), .A1(n7367) );
  nor02 U5710 ( .Y(n6971), .A0(n6972), .A1(n6973) );
  nor02 U5711 ( .Y(n6975), .A0(n7482), .A1(n5486) );
  nor02 U5712 ( .Y(n6976), .A0(n7507), .A1(n7372) );
  inv01 U5713 ( .Y(n6977), .A(n7508) );
  nor02 U5714 ( .Y(n6974), .A0(n6977), .A1(n6978) );
  nor02 U5715 ( .Y(n6979), .A0(n6975), .A1(n6976) );
  inv01 U5716 ( .Y(n6978), .A(n6979) );
  inv02 U5717 ( .Y(n7507), .A(n7528) );
  nor02 U5718 ( .Y(n6981), .A0(n7502), .A1(n7387) );
  nor02 U5719 ( .Y(n6982), .A0(n7501), .A1(n7372) );
  inv01 U5720 ( .Y(n6983), .A(n7503) );
  nor02 U5721 ( .Y(n6980), .A0(n6983), .A1(n6984) );
  nor02 U5722 ( .Y(n6985), .A0(n6981), .A1(n6982) );
  inv01 U5723 ( .Y(n6984), .A(n6985) );
  inv02 U5724 ( .Y(s_op2_40_), .A(n6986) );
  nor02 U5725 ( .Y(n6987), .A0(n7518), .A1(n7387) );
  nor02 U5726 ( .Y(n6988), .A0(n7517), .A1(n7372) );
  inv01 U5727 ( .Y(n6989), .A(n7519) );
  nor02 U5728 ( .Y(n6986), .A0(n6989), .A1(n6990) );
  nor02 U5729 ( .Y(n6991), .A0(n6987), .A1(n6988) );
  inv01 U5730 ( .Y(n6990), .A(n6991) );
  inv02 U5731 ( .Y(s_op2_51_), .A(n6992) );
  nor02 U5732 ( .Y(n6993), .A0(n7444), .A1(n7387) );
  nor02 U5733 ( .Y(n6994), .A0(n7443), .A1(n7372) );
  inv01 U5734 ( .Y(n6995), .A(n7445) );
  nor02 U5735 ( .Y(n6992), .A0(n6995), .A1(n6996) );
  nor02 U5736 ( .Y(n6997), .A0(n6993), .A1(n6994) );
  inv01 U5737 ( .Y(n6996), .A(n6997) );
  inv04 U5738 ( .Y(n7372), .A(n7371) );
  nor02 U5739 ( .Y(n6999), .A0(n6409), .A1(n7387) );
  nor02 U5740 ( .Y(n7000), .A0(n7459), .A1(n7372) );
  inv01 U5741 ( .Y(n7001), .A(n7460) );
  nor02 U5742 ( .Y(n6998), .A0(n7001), .A1(n7002) );
  nor02 U5743 ( .Y(n7003), .A0(n6999), .A1(n7000) );
  inv01 U5744 ( .Y(n7002), .A(n7003) );
  inv02 U5745 ( .Y(s_op2_44_), .A(n7004) );
  nor02 U5746 ( .Y(n7005), .A0(n7496), .A1(n7387) );
  nor02 U5747 ( .Y(n7006), .A0(n7495), .A1(n7372) );
  inv01 U5748 ( .Y(n7007), .A(n7497) );
  nor02 U5749 ( .Y(n7004), .A0(n7007), .A1(n7008) );
  nor02 U5750 ( .Y(n7009), .A0(n7005), .A1(n7006) );
  inv01 U5751 ( .Y(n7008), .A(n7009) );
  inv02 U5752 ( .Y(s_op2_45_), .A(n7010) );
  nor02 U5753 ( .Y(n7011), .A0(n7490), .A1(n7387) );
  nor02 U5754 ( .Y(n7012), .A0(n7489), .A1(n7372) );
  inv01 U5755 ( .Y(n7013), .A(n7491) );
  nor02 U5756 ( .Y(n7010), .A0(n7013), .A1(n7014) );
  nor02 U5757 ( .Y(n7015), .A0(n7011), .A1(n7012) );
  inv01 U5758 ( .Y(n7014), .A(n7015) );
  inv02 U5759 ( .Y(s_op2_47_), .A(n7016) );
  nor02 U5760 ( .Y(n7017), .A0(n7478), .A1(n7387) );
  nor02 U5761 ( .Y(n7018), .A0(n7477), .A1(n7372) );
  inv01 U5762 ( .Y(n7019), .A(n7479) );
  nor02 U5763 ( .Y(n7016), .A0(n7019), .A1(n7020) );
  nor02 U5764 ( .Y(n7021), .A0(n7017), .A1(n7018) );
  inv01 U5765 ( .Y(n7020), .A(n7021) );
  nor02 U5766 ( .Y(n7023), .A0(n6365), .A1(n7387) );
  nor02 U5767 ( .Y(n7024), .A0(n7665), .A1(n5486) );
  inv01 U5768 ( .Y(n7025), .A(n7666) );
  nor02 U5769 ( .Y(n7022), .A0(n7025), .A1(n7026) );
  nor02 U5770 ( .Y(n7027), .A0(n7023), .A1(n7024) );
  inv01 U5771 ( .Y(n7026), .A(n7027) );
  inv02 U5772 ( .Y(s_op2_36_), .A(n7028) );
  nor02 U5773 ( .Y(n7029), .A0(n7539), .A1(n7387) );
  nor02 U5774 ( .Y(n7030), .A0(n7538), .A1(n7372) );
  inv01 U5775 ( .Y(n7031), .A(n7540) );
  nor02 U5776 ( .Y(n7028), .A0(n7031), .A1(n7032) );
  nor02 U5777 ( .Y(n7033), .A0(n7029), .A1(n7030) );
  inv01 U5778 ( .Y(n7032), .A(n7033) );
  inv02 U5779 ( .Y(s_op2_48_), .A(n7034) );
  nor02 U5780 ( .Y(n7035), .A0(n7469), .A1(n7387) );
  nor02 U5781 ( .Y(n7036), .A0(n7468), .A1(n7372) );
  inv01 U5782 ( .Y(n7037), .A(n7470) );
  nor02 U5783 ( .Y(n7034), .A0(n7037), .A1(n7038) );
  nor02 U5784 ( .Y(n7039), .A0(n7035), .A1(n7036) );
  inv01 U5785 ( .Y(n7038), .A(n7039) );
  inv02 U5786 ( .Y(s_op2_41_), .A(n7040) );
  nor02 U5787 ( .Y(n7041), .A0(n7512), .A1(n7387) );
  nor02 U5788 ( .Y(n7042), .A0(n7511), .A1(n7372) );
  inv01 U5789 ( .Y(n7043), .A(n7513) );
  nor02 U5790 ( .Y(n7040), .A0(n7043), .A1(n7044) );
  nor02 U5791 ( .Y(n7045), .A0(n7041), .A1(n7042) );
  inv01 U5792 ( .Y(n7044), .A(n7045) );
  inv02 U5793 ( .Y(s_op2_39_), .A(n7046) );
  nor02 U5794 ( .Y(n7047), .A0(n6574), .A1(n7387) );
  nor02 U5795 ( .Y(n7048), .A0(n7522), .A1(n7372) );
  inv01 U5796 ( .Y(n7049), .A(n7523) );
  nor02 U5797 ( .Y(n7046), .A0(n7049), .A1(n7050) );
  nor02 U5798 ( .Y(n7051), .A0(n7047), .A1(n7048) );
  inv01 U5799 ( .Y(n7050), .A(n7051) );
  inv02 U5800 ( .Y(s_op2_37_), .A(n7052) );
  nor02 U5801 ( .Y(n7053), .A0(n7532), .A1(n7387) );
  nor02 U5802 ( .Y(n7054), .A0(n7531), .A1(n7372) );
  inv01 U5803 ( .Y(n7055), .A(n7533) );
  nor02 U5804 ( .Y(n7052), .A0(n7055), .A1(n7056) );
  nor02 U5805 ( .Y(n7057), .A0(n7053), .A1(n7054) );
  inv01 U5806 ( .Y(n7056), .A(n7057) );
  nor02 U5807 ( .Y(n7059), .A0(n7483), .A1(n5486) );
  nor02 U5808 ( .Y(n7060), .A0(n7482), .A1(n7372) );
  inv01 U5809 ( .Y(n7061), .A(n7485) );
  nor02 U5810 ( .Y(n7058), .A0(n7061), .A1(n7062) );
  nor02 U5811 ( .Y(n7063), .A0(n7059), .A1(n7060) );
  inv01 U5812 ( .Y(n7062), .A(n7063) );
  inv02 U5813 ( .Y(n7482), .A(n7530) );
  inv02 U5814 ( .Y(n7483), .A(n7510) );
  nor02 U5815 ( .Y(n7065), .A0(n7436), .A1(n7367) );
  nor02 U5816 ( .Y(n7066), .A0(n7438), .A1(n7602) );
  nor02 U5817 ( .Y(n7067), .A0(n7378), .A1(n6574) );
  nor02 U5818 ( .Y(n7064), .A0(n7067), .A1(n7068) );
  nor02 U5819 ( .Y(n7069), .A0(n7065), .A1(n7066) );
  inv01 U5820 ( .Y(n7068), .A(n7069) );
  inv02 U5821 ( .Y(n7438), .A(n7621) );
  nor02 U5822 ( .Y(n7071), .A0(n7442), .A1(n7367) );
  nor02 U5823 ( .Y(n7072), .A0(n7366), .A1(n7602) );
  nor02 U5824 ( .Y(n7073), .A0(n7378), .A1(n7532) );
  nor02 U5825 ( .Y(n7070), .A0(n7073), .A1(n7074) );
  nor02 U5826 ( .Y(n7075), .A0(n7071), .A1(n7072) );
  inv01 U5827 ( .Y(n7074), .A(n7075) );
  inv02 U5828 ( .Y(s_op2_38_), .A(n7076) );
  inv01 U5829 ( .Y(n7077), .A(n7446) );
  inv01 U5830 ( .Y(n7078), .A(n7528) );
  inv01 U5831 ( .Y(n7079), .A(n6108) );
  inv01 U5832 ( .Y(n7080), .A(n7526) );
  nor02 U5833 ( .Y(n7081), .A0(n7077), .A1(n7078) );
  nor02 U5834 ( .Y(n7082), .A0(n7079), .A1(n7080) );
  nor02 U5835 ( .Y(n7076), .A0(n7529), .A1(n7083) );
  nor02 U5836 ( .Y(n7084), .A0(n7081), .A1(n7082) );
  inv01 U5837 ( .Y(n7083), .A(n7084) );
  inv02 U5838 ( .Y(s_op2_22_), .A(n7085) );
  nor02 U5839 ( .Y(n7086), .A0(n7440), .A1(n7367) );
  nor02 U5840 ( .Y(n7087), .A0(n7364), .A1(n7602) );
  nor02 U5841 ( .Y(n7088), .A0(n7378), .A1(n6829) );
  nor02 U5842 ( .Y(n7085), .A0(n7088), .A1(n7089) );
  nor02 U5843 ( .Y(n7090), .A0(n7086), .A1(n7087) );
  inv01 U5844 ( .Y(n7089), .A(n7090) );
  inv02 U5845 ( .Y(n7366), .A(n7365) );
  inv02 U5846 ( .Y(n7442), .A(n7593) );
  ao22 U5847 ( .Y(n7091), .A0(n7551), .A1(n7377), .B0(n6365), .B1(n7387) );
  inv01 U5848 ( .Y(n7092), .A(n7091) );
  inv02 U5849 ( .Y(n7093), .A(n7091) );
  ao22 U5850 ( .Y(n7094), .A0(n6298), .A1(n7377), .B0(n7490), .B1(n7387) );
  inv02 U5851 ( .Y(n7095), .A(n7094) );
  ao22 U5852 ( .Y(n7096), .A0(n7584), .A1(n7377), .B0(n7585), .B1(n7387) );
  inv02 U5853 ( .Y(n7097), .A(n7096) );
  ao22 U5854 ( .Y(n7098), .A0(n7579), .A1(n7377), .B0(n7502), .B1(n7387) );
  inv02 U5855 ( .Y(n7099), .A(n7098) );
  ao22 U5856 ( .Y(n7100), .A0(n6300), .A1(n7380), .B0(n7565), .B1(n7387) );
  inv01 U5857 ( .Y(n7101), .A(n7100) );
  inv02 U5858 ( .Y(n7102), .A(n7100) );
  ao22 U5859 ( .Y(n7103), .A0(n6501), .A1(n7380), .B0(n7444), .B1(n7387) );
  inv02 U5860 ( .Y(n7104), .A(n7103) );
  ao22 U5861 ( .Y(n7105), .A0(n7614), .A1(n7380), .B0(n7539), .B1(n7387) );
  inv02 U5862 ( .Y(n7106), .A(n7105) );
  ao22 U5863 ( .Y(n7107), .A0(n6503), .A1(n7380), .B0(n7469), .B1(n7387) );
  inv02 U5864 ( .Y(n7108), .A(n7107) );
  ao22 U5865 ( .Y(n7109), .A0(n7435), .A1(n7379), .B0(n7518), .B1(n7387) );
  inv01 U5866 ( .Y(n7110), .A(n7109) );
  inv02 U5867 ( .Y(n7111), .A(n7109) );
  ao22 U5868 ( .Y(n7112), .A0(n7434), .A1(n7379), .B0(n7512), .B1(n7387) );
  inv02 U5869 ( .Y(n7113), .A(n7112) );
  ao22 U5870 ( .Y(n7114), .A0(n7575), .A1(n7379), .B0(n7496), .B1(n7387) );
  inv02 U5871 ( .Y(n7115), .A(n7114) );
  ao22 U5872 ( .Y(n7116), .A0(n7552), .A1(n7379), .B0(n6409), .B1(n7387) );
  inv02 U5873 ( .Y(n7117), .A(n7116) );
  ao22 U5874 ( .Y(n7118), .A0(n6296), .A1(n7379), .B0(n7478), .B1(n7387) );
  inv02 U5875 ( .Y(n7119), .A(n7118) );
  inv02 U5876 ( .Y(n7641), .A(r0_2_) );
  inv04 U5877 ( .Y(n7122), .A(n7582) );
  inv02 U5878 ( .Y(n7608), .A(n7126) );
  nor02 U5879 ( .Y(n7127), .A0(n7660), .A1(n7393) );
  nor02 U5880 ( .Y(n7128), .A0(n7404), .A1(n7642) );
  inv01 U5881 ( .Y(n7129), .A(n7664) );
  nor02 U5882 ( .Y(n7126), .A0(n7129), .A1(n7130) );
  nor02 U5883 ( .Y(n7131), .A0(n7127), .A1(n7128) );
  inv01 U5884 ( .Y(n7130), .A(n7131) );
  inv02 U5885 ( .Y(n7525), .A(n7132) );
  nor02 U5886 ( .Y(n7133), .A0(n7393), .A1(n7578) );
  nor02 U5887 ( .Y(n7134), .A0(n7404), .A1(n7582) );
  inv01 U5888 ( .Y(n7135), .A(n7583) );
  nor02 U5889 ( .Y(n7132), .A0(n7135), .A1(n7136) );
  nor02 U5890 ( .Y(n7137), .A0(n7133), .A1(n7134) );
  inv01 U5891 ( .Y(n7136), .A(n7137) );
  inv02 U5892 ( .Y(n7440), .A(n7608) );
  inv02 U5893 ( .Y(n7642), .A(r0_3_) );
  inv02 U5894 ( .Y(n7582), .A(r0_24_) );
  inv02 U5895 ( .Y(n7604), .A(n7138) );
  nor02 U5896 ( .Y(n7139), .A0(n7649), .A1(n7394) );
  nor02 U5897 ( .Y(n7140), .A0(n7660), .A1(n7404) );
  inv01 U5898 ( .Y(n7141), .A(n7661) );
  nor02 U5899 ( .Y(n7138), .A0(n7141), .A1(n7142) );
  nor02 U5900 ( .Y(n7143), .A0(n7139), .A1(n7140) );
  inv01 U5901 ( .Y(n7142), .A(n7143) );
  inv02 U5902 ( .Y(n7436), .A(n7604) );
  inv02 U5903 ( .Y(n7660), .A(r0_4_) );
  inv08 U5904 ( .Y(n7145), .A(n7144) );
  inv02 U5905 ( .Y(n7521), .A(n7146) );
  nor02 U5906 ( .Y(n7147), .A0(n7394), .A1(n7573) );
  nor02 U5907 ( .Y(n7148), .A0(n7403), .A1(n7578) );
  inv01 U5908 ( .Y(n7149), .A(n3543) );
  nor02 U5909 ( .Y(n7146), .A0(n7149), .A1(n7150) );
  nor02 U5910 ( .Y(n7151), .A0(n7147), .A1(n7148) );
  inv01 U5911 ( .Y(n7150), .A(n7151) );
  inv02 U5912 ( .Y(n7506), .A(n7152) );
  nor02 U5913 ( .Y(n7153), .A0(n7393), .A1(n7559) );
  nor02 U5914 ( .Y(n7154), .A0(n7403), .A1(n7563) );
  inv01 U5915 ( .Y(n7155), .A(n7564) );
  nor02 U5916 ( .Y(n7152), .A0(n7155), .A1(n7156) );
  nor02 U5917 ( .Y(n7157), .A0(n7153), .A1(n7154) );
  inv01 U5918 ( .Y(n7156), .A(n7157) );
  inv02 U5919 ( .Y(n7516), .A(n7158) );
  nor02 U5920 ( .Y(n7159), .A0(n7395), .A1(n7574) );
  nor02 U5921 ( .Y(n7160), .A0(n7404), .A1(n7573) );
  inv01 U5922 ( .Y(n7161), .A(n3501) );
  nor02 U5923 ( .Y(n7158), .A0(n7161), .A1(n7162) );
  nor02 U5924 ( .Y(n7163), .A0(n7159), .A1(n7160) );
  inv01 U5925 ( .Y(n7162), .A(n7163) );
  inv02 U5926 ( .Y(n7578), .A(r0_25_) );
  inv02 U5927 ( .Y(n7573), .A(r0_26_) );
  inv02 U5928 ( .Y(n7563), .A(r0_28_) );
  inv02 U5929 ( .Y(n7574), .A(r0_27_) );
  inv04 U5930 ( .Y(n7652), .A(r0_1_) );
  inv02 U5931 ( .Y(n7166), .A(r0_23_) );
  inv02 U5932 ( .Y(n7537), .A(n7168) );
  nor02 U5933 ( .Y(n7169), .A0(n7395), .A1(n7591) );
  nor02 U5934 ( .Y(n7170), .A0(n7403), .A1(n7590) );
  inv01 U5935 ( .Y(n7171), .A(n7592) );
  nor02 U5936 ( .Y(n7168), .A0(n7171), .A1(n7172) );
  nor02 U5937 ( .Y(n7173), .A0(n7169), .A1(n7170) );
  inv01 U5938 ( .Y(n7172), .A(n7173) );
  inv02 U5939 ( .Y(n7543), .A(n7174) );
  nor02 U5940 ( .Y(n7175), .A0(n7394), .A1(n7590) );
  nor02 U5941 ( .Y(n7176), .A0(n7403), .A1(n7598) );
  inv01 U5942 ( .Y(n7177), .A(n3597) );
  nor02 U5943 ( .Y(n7174), .A0(n7177), .A1(n7178) );
  nor02 U5944 ( .Y(n7179), .A0(n7175), .A1(n7176) );
  inv01 U5945 ( .Y(n7178), .A(n7179) );
  inv02 U5946 ( .Y(n7590), .A(r0_22_) );
  inv02 U5947 ( .Y(n7591), .A(r0_23_) );
  inv02 U5948 ( .Y(n7500), .A(n7180) );
  nor02 U5949 ( .Y(n7181), .A0(n7394), .A1(n7555) );
  nor02 U5950 ( .Y(n7182), .A0(n7403), .A1(n7559) );
  inv01 U5951 ( .Y(n7183), .A(n7560) );
  nor02 U5952 ( .Y(n7180), .A0(n7183), .A1(n7184) );
  nor02 U5953 ( .Y(n7185), .A0(n7181), .A1(n7182) );
  inv01 U5954 ( .Y(n7184), .A(n7185) );
  inv02 U5955 ( .Y(n7559), .A(r0_29_) );
  inv02 U5956 ( .Y(n7481), .A(n7188) );
  nor02 U5957 ( .Y(n7189), .A0(n7393), .A1(n7541) );
  nor02 U5958 ( .Y(n7190), .A0(n7403), .A1(n7550) );
  inv01 U5959 ( .Y(n7191), .A(n3571) );
  nor02 U5960 ( .Y(n7188), .A0(n7191), .A1(n7192) );
  nor02 U5961 ( .Y(n7193), .A0(n7189), .A1(n7190) );
  inv01 U5962 ( .Y(n7192), .A(n7193) );
  inv02 U5963 ( .Y(n7494), .A(n7194) );
  nor02 U5964 ( .Y(n7195), .A0(n7395), .A1(n7556) );
  nor02 U5965 ( .Y(n7196), .A0(n7403), .A1(n7555) );
  inv01 U5966 ( .Y(n7197), .A(n3503) );
  nor02 U5967 ( .Y(n7194), .A0(n7197), .A1(n7198) );
  nor02 U5968 ( .Y(n7199), .A0(n7195), .A1(n7196) );
  inv01 U5969 ( .Y(n7198), .A(n7199) );
  inv02 U5970 ( .Y(n7550), .A(r0_32_) );
  inv02 U5971 ( .Y(n7555), .A(r0_30_) );
  inv02 U5972 ( .Y(n7556), .A(r0_31_) );
  inv02 U5973 ( .Y(n7589), .A(n7215) );
  nor02 U5974 ( .Y(n7216), .A0(n7395), .A1(n7636) );
  nor02 U5975 ( .Y(n7217), .A0(n7404), .A1(n7644) );
  inv01 U5976 ( .Y(n7218), .A(n7645) );
  nor02 U5977 ( .Y(n7215), .A0(n7218), .A1(n7219) );
  nor02 U5978 ( .Y(n7220), .A0(n7216), .A1(n7217) );
  inv01 U5979 ( .Y(n7219), .A(n7220) );
  inv02 U5980 ( .Y(n7601), .A(n7221) );
  nor02 U5981 ( .Y(n7222), .A0(n7393), .A1(n7646) );
  nor02 U5982 ( .Y(n7223), .A0(n7649), .A1(n7404) );
  inv01 U5983 ( .Y(n7224), .A(n7650) );
  nor02 U5984 ( .Y(n7221), .A0(n7224), .A1(n7225) );
  nor02 U5985 ( .Y(n7226), .A0(n7222), .A1(n7223) );
  inv01 U5986 ( .Y(n7225), .A(n7226) );
  inv02 U5987 ( .Y(n7649), .A(r0_5_) );
  buf08 U5988 ( .Y(n7393), .A(n7454) );
  inv02 U5989 ( .Y(n7609), .A(n7227) );
  nor02 U5990 ( .Y(n7228), .A0(n7393), .A1(n7656) );
  nor02 U5991 ( .Y(n7229), .A0(n7404), .A1(n7647) );
  inv01 U5992 ( .Y(n7230), .A(n7662) );
  nor02 U5993 ( .Y(n7227), .A0(n7230), .A1(n7231) );
  nor02 U5994 ( .Y(n7232), .A0(n7228), .A1(n7229) );
  inv01 U5995 ( .Y(n7231), .A(n7232) );
  inv02 U5996 ( .Y(n7558), .A(n7233) );
  nor02 U5997 ( .Y(n7234), .A0(n7394), .A1(n7612) );
  nor02 U5998 ( .Y(n7235), .A0(n7403), .A1(n7616) );
  inv01 U5999 ( .Y(n7236), .A(n3701) );
  nor02 U6000 ( .Y(n7233), .A0(n7236), .A1(n7237) );
  nor02 U6001 ( .Y(n7238), .A0(n7234), .A1(n7235) );
  inv01 U6002 ( .Y(n7237), .A(n7238) );
  inv02 U6003 ( .Y(n7562), .A(n7239) );
  nor02 U6004 ( .Y(n7240), .A0(n7393), .A1(n7616) );
  nor02 U6005 ( .Y(n7241), .A0(n7403), .A1(n7620) );
  inv01 U6006 ( .Y(n7242), .A(n3517) );
  nor02 U6007 ( .Y(n7239), .A0(n7242), .A1(n7243) );
  nor02 U6008 ( .Y(n7244), .A0(n7240), .A1(n7241) );
  inv01 U6009 ( .Y(n7243), .A(n7244) );
  inv02 U6010 ( .Y(n7549), .A(n7245) );
  nor02 U6011 ( .Y(n7246), .A0(n7393), .A1(n7598) );
  nor02 U6012 ( .Y(n7247), .A0(n7403), .A1(n7607) );
  inv01 U6013 ( .Y(n7248), .A(n3798) );
  nor02 U6014 ( .Y(n7245), .A0(n7248), .A1(n7249) );
  nor02 U6015 ( .Y(n7250), .A0(n7246), .A1(n7247) );
  inv01 U6016 ( .Y(n7249), .A(n7250) );
  inv02 U6017 ( .Y(n7616), .A(r0_17_) );
  inv02 U6018 ( .Y(n7607), .A(r0_20_) );
  inv02 U6019 ( .Y(n7598), .A(r0_21_) );
  inv02 U6020 ( .Y(n7581), .A(n7251) );
  nor02 U6021 ( .Y(n7252), .A0(n7395), .A1(n7629) );
  nor02 U6022 ( .Y(n7253), .A0(n7404), .A1(n7632) );
  inv01 U6023 ( .Y(n7254), .A(n7633) );
  nor02 U6024 ( .Y(n7251), .A0(n7254), .A1(n7255) );
  nor02 U6025 ( .Y(n7256), .A0(n7252), .A1(n7253) );
  inv01 U6026 ( .Y(n7255), .A(n7256) );
  inv02 U6027 ( .Y(n7606), .A(n7257) );
  nor02 U6028 ( .Y(n7258), .A0(n7394), .A1(n7654) );
  nor02 U6029 ( .Y(n7259), .A0(n7404), .A1(n7656) );
  inv01 U6030 ( .Y(n7260), .A(n7657) );
  nor02 U6031 ( .Y(n7257), .A0(n7260), .A1(n7261) );
  nor02 U6032 ( .Y(n7262), .A0(n7258), .A1(n7259) );
  inv01 U6033 ( .Y(n7261), .A(n7262) );
  inv02 U6034 ( .Y(n7554), .A(n7263) );
  nor02 U6035 ( .Y(n7264), .A0(n7395), .A1(n7613) );
  nor02 U6036 ( .Y(n7265), .A0(n7403), .A1(n7612) );
  inv01 U6037 ( .Y(n7266), .A(n3635) );
  nor02 U6038 ( .Y(n7263), .A0(n7266), .A1(n7267) );
  nor02 U6039 ( .Y(n7268), .A0(n7264), .A1(n7265) );
  inv01 U6040 ( .Y(n7267), .A(n7268) );
  inv02 U6041 ( .Y(n7656), .A(r0_8_) );
  inv02 U6042 ( .Y(n7612), .A(r0_18_) );
  inv02 U6043 ( .Y(n7613), .A(r0_19_) );
  inv02 U6044 ( .Y(n7597), .A(n7269) );
  nor02 U6045 ( .Y(n7270), .A0(n7395), .A1(n7644) );
  nor02 U6046 ( .Y(n7271), .A0(n7404), .A1(n7654) );
  inv01 U6047 ( .Y(n7272), .A(n7655) );
  nor02 U6048 ( .Y(n7269), .A0(n7272), .A1(n7273) );
  nor02 U6049 ( .Y(n7274), .A0(n7270), .A1(n7271) );
  inv01 U6050 ( .Y(n7273), .A(n7274) );
  inv02 U6051 ( .Y(n7654), .A(r0_9_) );
  inv02 U6052 ( .Y(n7644), .A(r0_10_) );
  inv02 U6053 ( .Y(n7595), .A(n7275) );
  nor02 U6054 ( .Y(n7276), .A0(n7394), .A1(n7647) );
  nor02 U6055 ( .Y(n7277), .A0(n7404), .A1(n7646) );
  inv01 U6056 ( .Y(n7278), .A(n7648) );
  nor02 U6057 ( .Y(n7275), .A0(n7278), .A1(n7279) );
  nor02 U6058 ( .Y(n7280), .A0(n7276), .A1(n7277) );
  inv01 U6059 ( .Y(n7279), .A(n7280) );
  inv02 U6060 ( .Y(n7646), .A(r0_6_) );
  inv02 U6061 ( .Y(n7647), .A(r0_7_) );
  inv02 U6062 ( .Y(n7587), .A(n7281) );
  nor02 U6063 ( .Y(n7282), .A0(n7394), .A1(n7632) );
  nor02 U6064 ( .Y(n7283), .A0(n7404), .A1(n7636) );
  inv01 U6065 ( .Y(n7284), .A(n7637) );
  nor02 U6066 ( .Y(n7281), .A0(n7284), .A1(n7285) );
  nor02 U6067 ( .Y(n7286), .A0(n7282), .A1(n7283) );
  inv01 U6068 ( .Y(n7285), .A(n7286) );
  inv02 U6069 ( .Y(n7476), .A(n7287) );
  nor02 U6070 ( .Y(n7288), .A0(n7394), .A1(n7534) );
  nor02 U6071 ( .Y(n7289), .A0(n7403), .A1(n7541) );
  inv01 U6072 ( .Y(n7290), .A(n7542) );
  nor02 U6073 ( .Y(n7287), .A0(n7290), .A1(n7291) );
  nor02 U6074 ( .Y(n7292), .A0(n7288), .A1(n7289) );
  inv01 U6075 ( .Y(n7291), .A(n7292) );
  inv02 U6076 ( .Y(n7458), .A(n7293) );
  nor02 U6077 ( .Y(n7294), .A0(n7393), .A1(n7520) );
  nor02 U6078 ( .Y(n7295), .A0(n7403), .A1(n7524) );
  inv01 U6079 ( .Y(n7296), .A(n3730) );
  nor02 U6080 ( .Y(n7293), .A0(n7296), .A1(n7297) );
  nor02 U6081 ( .Y(n7298), .A0(n7294), .A1(n7295) );
  inv01 U6082 ( .Y(n7297), .A(n7298) );
  inv02 U6083 ( .Y(n7467), .A(n7299) );
  nor02 U6084 ( .Y(n7300), .A0(n7395), .A1(n7535) );
  nor02 U6085 ( .Y(n7301), .A0(n7403), .A1(n7534) );
  inv01 U6086 ( .Y(n7302), .A(n7536) );
  nor02 U6087 ( .Y(n7299), .A0(n7302), .A1(n7303) );
  nor02 U6088 ( .Y(n7304), .A0(n7300), .A1(n7301) );
  inv01 U6089 ( .Y(n7303), .A(n7304) );
  inv02 U6090 ( .Y(n7636), .A(r0_11_) );
  inv02 U6091 ( .Y(n7632), .A(r0_12_) );
  inv02 U6092 ( .Y(n7541), .A(r0_33_) );
  inv02 U6093 ( .Y(n7534), .A(r0_34_) );
  inv02 U6094 ( .Y(n7524), .A(r0_36_) );
  inv02 U6095 ( .Y(n7520), .A(r0_37_) );
  inv02 U6096 ( .Y(n7535), .A(r0_35_) );
  inv02 U6097 ( .Y(n7572), .A(n7305) );
  nor02 U6098 ( .Y(n7306), .A0(n7394), .A1(n7623) );
  nor02 U6099 ( .Y(n7307), .A0(n7404), .A1(n7625) );
  inv01 U6100 ( .Y(n7308), .A(n7626) );
  nor02 U6101 ( .Y(n7305), .A0(n7308), .A1(n7309) );
  nor02 U6102 ( .Y(n7310), .A0(n7306), .A1(n7307) );
  inv01 U6103 ( .Y(n7309), .A(n7310) );
  inv02 U6104 ( .Y(n7577), .A(n7311) );
  nor02 U6105 ( .Y(n7312), .A0(n7393), .A1(n7625) );
  nor02 U6106 ( .Y(n7313), .A0(n7404), .A1(n7629) );
  inv01 U6107 ( .Y(n7314), .A(n7630) );
  nor02 U6108 ( .Y(n7311), .A0(n7314), .A1(n7315) );
  nor02 U6109 ( .Y(n7316), .A0(n7312), .A1(n7313) );
  inv01 U6110 ( .Y(n7315), .A(n7316) );
  inv02 U6111 ( .Y(n7625), .A(r0_14_) );
  inv02 U6112 ( .Y(n7629), .A(r0_13_) );
  inv02 U6113 ( .Y(n7569), .A(n7317) );
  nor02 U6114 ( .Y(n7318), .A0(n7395), .A1(n7620) );
  nor02 U6115 ( .Y(n7319), .A0(n7404), .A1(n7623) );
  inv01 U6116 ( .Y(n7320), .A(n3796) );
  nor02 U6117 ( .Y(n7317), .A0(n7320), .A1(n7321) );
  nor02 U6118 ( .Y(n7322), .A0(n7318), .A1(n7319) );
  inv01 U6119 ( .Y(n7321), .A(n7322) );
  inv02 U6120 ( .Y(n7623), .A(r0_15_) );
  inv02 U6121 ( .Y(n7620), .A(r0_16_) );
  or02 U6122 ( .Y(n7323), .A0(n7364), .A1(n7437) );
  inv02 U6123 ( .Y(n7324), .A(n7323) );
  or02 U6124 ( .Y(n7325), .A0(n7366), .A1(n7437) );
  inv02 U6125 ( .Y(n7326), .A(n7325) );
  nor02 U6126 ( .Y(n7327), .A0(n7438), .A1(n7437) );
  or02 U6127 ( .Y(n7328), .A0(n7627), .A1(n7437) );
  inv02 U6128 ( .Y(n7329), .A(n7328) );
  inv01 U6129 ( .Y(n7330), .A(n7328) );
  or02 U6130 ( .Y(n7331), .A0(n7380), .A1(n6298) );
  inv02 U6131 ( .Y(n7332), .A(n7331) );
  or02 U6132 ( .Y(n7333), .A0(n7377), .A1(n6296) );
  inv02 U6133 ( .Y(n7334), .A(n7333) );
  or02 U6134 ( .Y(n7335), .A0(n7377), .A1(n6300) );
  inv02 U6135 ( .Y(n7336), .A(n7335) );
  or02 U6136 ( .Y(n7337), .A0(n7379), .A1(n7584) );
  inv01 U6137 ( .Y(n7338), .A(n7337) );
  inv02 U6138 ( .Y(n7339), .A(n7337) );
  or02 U6139 ( .Y(n7340), .A0(n7379), .A1(n7435) );
  inv02 U6140 ( .Y(n7341), .A(n7340) );
  or02 U6141 ( .Y(n7342), .A0(n7380), .A1(n7434) );
  inv02 U6142 ( .Y(n7343), .A(n7342) );
  or02 U6143 ( .Y(n7344), .A0(n7379), .A1(n7575) );
  inv02 U6144 ( .Y(n7345), .A(n7344) );
  or02 U6145 ( .Y(n7346), .A0(n7380), .A1(n7579) );
  inv02 U6146 ( .Y(n7347), .A(n7346) );
  inv01 U6147 ( .Y(n7349), .A(n8007) );
  inv01 U6148 ( .Y(n7350), .A(s_count_1_) );
  inv01 U6149 ( .Y(n7351), .A(s_count_0_) );
  nand02 U6150 ( .Y(n7348), .A0(n7351), .A1(n7352) );
  nand02 U6151 ( .Y(n7353), .A0(n7349), .A1(n7350) );
  inv01 U6152 ( .Y(n7352), .A(n7353) );
  inv02 U6153 ( .Y(n7677), .A(n7676) );
  inv02 U6154 ( .Y(s_op2_4_), .A(n7354) );
  inv01 U6155 ( .Y(n7355), .A(c_3_) );
  inv01 U6156 ( .Y(n7356), .A(n7379) );
  inv01 U6157 ( .Y(n7357), .A(n3079) );
  nand02 U6158 ( .Y(n7354), .A0(n7357), .A1(n7358) );
  nand02 U6159 ( .Y(n7359), .A0(n7355), .A1(n7356) );
  inv01 U6160 ( .Y(n7358), .A(n7359) );
  or02 U6161 ( .Y(n7360), .A0(n7421), .A1(n6950) );
  inv01 U6162 ( .Y(n7361), .A(n7360) );
  inv01 U6163 ( .Y(n7363), .A(n7360) );
  inv01 U6164 ( .Y(n7362), .A(n7360) );
  buf02 U6165 ( .Y(n7364), .A(n7441) );
  ao22 U6166 ( .Y(n7365), .A0(n7399), .A1(n7164), .B0(n7401), .B1(r0_0_) );
  buf04 U6167 ( .Y(n7367), .A(n7603) );
  buf08 U6168 ( .Y(n7370), .A(n7450) );
  inv04 U6169 ( .Y(n7437), .A(n7369) );
  buf02 U6170 ( .Y(n7371), .A(n6108) );
  inv02 U6171 ( .Y(n7373), .A(n7548) );
  inv04 U6172 ( .Y(n7374), .A(n7373) );
  inv04 U6173 ( .Y(n7375), .A(n7373) );
  inv08 U6174 ( .Y(n7376), .A(c_4_) );
  inv04 U6175 ( .Y(n7380), .A(n7376) );
  inv04 U6176 ( .Y(n7379), .A(n7376) );
  inv12 U6177 ( .Y(n7771), .A(n6204) );
  nand02 U6178 ( .Y(n7381), .A0(n____return1071), .A1(n7382) );
  nand02 U6179 ( .Y(n7383), .A0(n7385), .A1(n7787) );
  inv01 U6180 ( .Y(n7382), .A(n7383) );
  inv02 U6181 ( .Y(n7787), .A(n7420) );
  buf08 U6182 ( .Y(n7384), .A(n7547) );
  buf12 U6183 ( .Y(n7385), .A(n7769) );
  buf02 U6184 ( .Y(n7386), .A(n7379) );
  buf12 U6185 ( .Y(n7388), .A(n7545) );
  buf12 U6186 ( .Y(n7389), .A(n4257) );
  buf12 U6187 ( .Y(n7390), .A(n7544) );
  nand02 U6188 ( .Y(n7391), .A0(n6944), .A1(n7674) );
  nand02 U6189 ( .Y(n7392), .A0(n6944), .A1(n7674) );
  nor02 U6190 ( .Y(n7396), .A0(n6945), .A1(c_0_) );
  nor02 U6191 ( .Y(n7397), .A0(n6945), .A1(c_0_) );
  buf08 U6192 ( .Y(n7398), .A(n7457) );
  buf08 U6193 ( .Y(n7400), .A(n7397) );
  buf16 U6194 ( .Y(n7401), .A(n4161) );
  inv04 U6195 ( .Y(n7402), .A(n7452) );
  nand02 U6196 ( .Y(n7405), .A0(n____return912), .A1(n7428) );
  nand02 U6197 ( .Y(n7406), .A0(n____return912), .A1(n7428) );
  buf16 U6198 ( .Y(n7407), .A(n7789) );
  buf16 U6199 ( .Y(n7408), .A(n7405) );
  buf16 U6200 ( .Y(n7409), .A(n7406) );
  inv16 U6201 ( .Y(n7411), .A(n6107) );
  inv16 U6202 ( .Y(n7413), .A(n6107) );
  inv16 U6203 ( .Y(n7412), .A(n6107) );
  inv12 U6204 ( .Y(n7414), .A(n6203) );
  inv12 U6205 ( .Y(n7415), .A(n7414) );
  inv12 U6206 ( .Y(n7417), .A(n7414) );
  inv12 U6207 ( .Y(n7416), .A(n7414) );
  inv08 U6208 ( .Y(n7418), .A(s_state110) );
  inv12 U6209 ( .Y(n7419), .A(n7418) );
  inv12 U6210 ( .Y(n7421), .A(n7418) );
  inv12 U6211 ( .Y(n7420), .A(n7418) );
  inv16 U6212 ( .Y(n7423), .A(n7422) );
  inv16 U6213 ( .Y(n7425), .A(n6106) );
  inv16 U6214 ( .Y(n7424), .A(n6106) );
  buf12 U6215 ( .Y(n7426), .A(n7788) );
  inv16 U6216 ( .Y(n7427), .A(n7426) );
  inv16 U6217 ( .Y(n7429), .A(n7426) );
  inv16 U6218 ( .Y(n7428), .A(n7426) );
  buf12 U6219 ( .Y(n7430), .A(n7361) );
  inv16 U6220 ( .Y(n7431), .A(n7430) );
  inv16 U6221 ( .Y(n7433), .A(n7430) );
  inv16 U6222 ( .Y(n7432), .A(n7430) );
  inv01 U6223 ( .Y(n7443), .A(n7458) );
  inv01 U6224 ( .Y(n7459), .A(n7467) );
  inv01 U6225 ( .Y(n7468), .A(n7476) );
  inv01 U6226 ( .Y(n7477), .A(n7481) );
  inv01 U6227 ( .Y(n7489), .A(n7494) );
  inv01 U6228 ( .Y(n7495), .A(n7500) );
  inv01 U6229 ( .Y(n7501), .A(n7506) );
  inv01 U6230 ( .Y(n7511), .A(n7516) );
  inv01 U6231 ( .Y(n7517), .A(n7521) );
  nor02 U6232 ( .Y(s_op2_3_), .A0(n7438), .A1(n7437) );
  inv01 U6233 ( .Y(n7522), .A(n7525) );
  inv01 U6234 ( .Y(n7531), .A(n7537) );
  inv01 U6235 ( .Y(n7538), .A(n7543) );
  ao22 U6236 ( .Y(n7546), .A0(n7384), .A1(n7525), .B0(n7374), .B1(n7549) );
  ao22 U6237 ( .Y(n7553), .A0(n7384), .A1(n7537), .B0(n7375), .B1(n7554) );
  ao22 U6238 ( .Y(n7557), .A0(n7384), .A1(n7543), .B0(n7375), .B1(n7558) );
  ao22 U6239 ( .Y(n7561), .A0(n7384), .A1(n7549), .B0(n7374), .B1(n7562) );
  inv01 U6240 ( .Y(n7565), .A(n7487) );
  ao22 U6241 ( .Y(n7571), .A0(n7384), .A1(n7554), .B0(n7375), .B1(n7572) );
  ao22 U6242 ( .Y(n7576), .A0(n7384), .A1(n7558), .B0(n7374), .B1(n7577) );
  ao22 U6243 ( .Y(n7580), .A0(n7384), .A1(n7562), .B0(n7375), .B1(n7581) );
  inv01 U6244 ( .Y(n7585), .A(n7509) );
  ao22 U6245 ( .Y(n7588), .A0(n7384), .A1(n7572), .B0(n7374), .B1(n7589) );
  inv01 U6246 ( .Y(n7594), .A(n7366) );
  ao22 U6247 ( .Y(n7596), .A0(n7384), .A1(n7577), .B0(n7375), .B1(n7597) );
  ao22 U6248 ( .Y(n7605), .A0(n7384), .A1(n7581), .B0(n7375), .B1(n7606) );
  ao22 U6249 ( .Y(n7610), .A0(n7388), .A1(n7569), .B0(n7384), .B1(n7587) );
  nand02 U6250 ( .Y(n7602), .A0(n7379), .A1(n7388) );
  ao22 U6251 ( .Y(n7611), .A0(n7374), .A1(n7595), .B0(n7384), .B1(n7589) );
  ao22 U6252 ( .Y(n7615), .A0(n7384), .A1(n7597), .B0(n7375), .B1(n7601) );
  nand02 U6253 ( .Y(n7614), .A0(n7617), .A1(n7618) );
  ao22 U6254 ( .Y(n7619), .A0(n7374), .A1(n7604), .B0(n7384), .B1(n7606) );
  ao22 U6255 ( .Y(n7622), .A0(n7374), .A1(n7608), .B0(n7384), .B1(n7609) );
  ao22 U6256 ( .Y(n7624), .A0(n7390), .A1(n7572), .B0(n7375), .B1(n7593) );
  nand02 U6257 ( .Y(n7603), .A0(n7380), .A1(n7390) );
  ao22 U6258 ( .Y(n7628), .A0(n7390), .A1(n7577), .B0(n7375), .B1(n7599) );
  ao22 U6259 ( .Y(n7631), .A0(n7384), .A1(n7604), .B0(n7388), .B1(n7606) );
  ao22 U6260 ( .Y(n7634), .A0(n7390), .A1(n7587), .B0(n7375), .B1(n7635) );
  inv01 U6261 ( .Y(n7617), .A(n3079) );
  inv01 U6262 ( .Y(n7600), .A(n7627) );
  inv01 U6263 ( .Y(n7635), .A(n7364) );
  nand02 U6264 ( .Y(n7627), .A0(n7398), .A1(n6906) );
  nor02 U6265 ( .Y(n7450), .A0(n7567), .A1(n7380) );
  nor02 U6266 ( .Y(n7448), .A0(n7568), .A1(n7377) );
  nor02 U6267 ( .Y(n7527), .A0(n7639), .A1(n7380) );
  nor02 U6268 ( .Y(n7548), .A0(n7651), .A1(n7618) );
  nor02 U6269 ( .Y(n7544), .A0(c_3_), .A1(c_2_) );
  nor02 U6270 ( .Y(n7545), .A0(n7651), .A1(c_3_) );
  nor02 U6271 ( .Y(n7446), .A0(n7640), .A1(n7379) );
  nor02 U6272 ( .Y(n7547), .A0(n7618), .A1(c_2_) );
  inv01 U6273 ( .Y(n7665), .A(n7486) );
  nor02 U6274 ( .Y(n7457), .A0(n6945), .A1(c_0_) );
  nand02 U6275 ( .Y(n7454), .A0(n6944), .A1(n7674) );
  nand02 U6276 ( .Y(n7452), .A0(n6944), .A1(c_0_) );
  nand04 U6277 ( .Y(n7681), .A0(n6110), .A1(n7682), .A2(n6144), .A3(n7683) );
  xor2 U6278 ( .Y(n7687), .A0(n____return1382_37_), .A1(s_rad_i_37_) );
  xor2 U6279 ( .Y(n7686), .A0(n____return1382_39_), .A1(s_rad_i_39_) );
  xor2 U6280 ( .Y(n7685), .A0(n____return1382_38_), .A1(n6272) );
  nand04 U6281 ( .Y(n7684), .A0(n4105), .A1(n4115), .A2(n4137), .A3(n4147) );
  xor2 U6282 ( .Y(n7691), .A0(n____return1382_42_), .A1(n6293) );
  xor2 U6283 ( .Y(n7690), .A0(n____return1382_44_), .A1(n6266) );
  xor2 U6284 ( .Y(n7689), .A0(n____return1382_43_), .A1(s_rad_i_43_) );
  nand03 U6285 ( .Y(n7688), .A0(n4053), .A1(n4069), .A2(n4101) );
  xor2 U6286 ( .Y(n7695), .A0(n____return1382_4_), .A1(n6284) );
  xor2 U6287 ( .Y(n7694), .A0(n____return1382_5_), .A1(s_rad_i_5_) );
  xor2 U6288 ( .Y(n7693), .A0(n____return1382_50_), .A1(n6275) );
  nand04 U6289 ( .Y(n7692), .A0(n4107), .A1(n4119), .A2(n4133), .A3(n4149) );
  xor2 U6290 ( .Y(n7699), .A0(n____return1382_9_), .A1(n6269) );
  xor2 U6291 ( .Y(n7698), .A0(n1384_51_), .A1(n6782) );
  xor2 U6292 ( .Y(n7697), .A0(n1384_49_), .A1(s_rad_i_49_) );
  nand03 U6293 ( .Y(n7696), .A0(n4059), .A1(n4051), .A2(n4091) );
  nand04 U6294 ( .Y(n7680), .A0(n6112), .A1(n7700), .A2(n6142), .A3(n7701) );
  xor2 U6295 ( .Y(n7705), .A0(n____return1382_13_), .A1(s_rad_i_13_) );
  xor2 U6296 ( .Y(n7704), .A0(n____return1382_15_), .A1(s_rad_i_15_) );
  xor2 U6297 ( .Y(n7703), .A0(n____return1382_14_), .A1(n6287) );
  nand04 U6298 ( .Y(n7702), .A0(n4083), .A1(n4113), .A2(n4129), .A3(n4159) );
  xor2 U6299 ( .Y(n7709), .A0(n____return1382_19_), .A1(s_rad_i_19_) );
  xor2 U6300 ( .Y(n7708), .A0(n____return1382_20_), .A1(n6278) );
  xor2 U6301 ( .Y(n7707), .A0(n____return1382_1_), .A1(s_rad_i_1_) );
  nand03 U6302 ( .Y(n7706), .A0(n4061), .A1(n4079), .A2(n4093) );
  xor2 U6303 ( .Y(n7713), .A0(n____return1382_25_), .A1(s_rad_i_25_) );
  xor2 U6304 ( .Y(n7712), .A0(n____return1382_27_), .A1(s_rad_i_27_) );
  xor2 U6305 ( .Y(n7711), .A0(n____return1382_26_), .A1(n6290) );
  nand04 U6306 ( .Y(n7710), .A0(n4085), .A1(n4127), .A2(n4139), .A3(n4155) );
  xor2 U6307 ( .Y(n7717), .A0(n____return1382_30_), .A1(s_rad_i_30_) );
  xor2 U6308 ( .Y(n7716), .A0(n____return1382_32_), .A1(n6281) );
  xor2 U6309 ( .Y(n7715), .A0(n____return1382_31_), .A1(s_rad_i_31_) );
  nand03 U6310 ( .Y(n7714), .A0(n4065), .A1(n4073), .A2(n4089) );
  nand04 U6311 ( .Y(n7679), .A0(n7718), .A1(n7719), .A2(n7720), .A3(n7721) );
  xnor2 U6312 ( .Y(n7723), .A0(n6271), .A1(n7726) );
  nand04 U6313 ( .Y(n7722), .A0(n4109), .A1(n4121), .A2(n4141), .A3(n4145) );
  xnor2 U6314 ( .Y(n7729), .A0(n6292), .A1(n7730) );
  xnor2 U6315 ( .Y(n7728), .A0(n6265), .A1(n7731) );
  nand03 U6316 ( .Y(n7727), .A0(n4055), .A1(n4067), .A2(n4103) );
  xnor2 U6317 ( .Y(n7735), .A0(n6274), .A1(n7737) );
  xnor2 U6318 ( .Y(n7734), .A0(n6283), .A1(n7738) );
  nand04 U6319 ( .Y(n7733), .A0(n4111), .A1(n4125), .A2(n4135), .A3(n4151) );
  xnor2 U6320 ( .Y(n7741), .A0(n6268), .A1(n7743) );
  xnor2 U6321 ( .Y(n7740), .A0(n6255), .A1(n7744) );
  nand03 U6322 ( .Y(n7739), .A0(n3800), .A1(n4071), .A2(n4099) );
  nand04 U6323 ( .Y(n7678), .A0(n7745), .A1(n7746), .A2(n7747), .A3(n7748) );
  xnor2 U6324 ( .Y(n7750), .A0(n6286), .A1(n7753) );
  nand04 U6325 ( .Y(n7749), .A0(n4087), .A1(n4123), .A2(n4131), .A3(n4157) );
  xnor2 U6326 ( .Y(n7755), .A0(n6277), .A1(n7757) );
  nand03 U6327 ( .Y(n7754), .A0(n4057), .A1(n4077), .A2(n4097) );
  xnor2 U6328 ( .Y(n7760), .A0(n6289), .A1(n7763) );
  nand04 U6329 ( .Y(n7759), .A0(n4081), .A1(n4117), .A2(n4143), .A3(n4153) );
  xnor2 U6330 ( .Y(n7765), .A0(n6280), .A1(n7767) );
  nand03 U6331 ( .Y(n7764), .A0(n4063), .A1(n4075), .A2(n4095) );
  inv01 U6332 ( .Y(n7769), .A(n6952) );
  ao21 U6333 ( .Y(n3049), .A0(n6950), .A1(n7677), .B0(n7420) );
  inv01 U6334 ( .Y(n7793), .A(r1_2_0_) );
  inv01 U6335 ( .Y(n7798), .A(r1_2_2_) );
  inv01 U6336 ( .Y(n7801), .A(r1_2_3_) );
  inv01 U6337 ( .Y(n7806), .A(r1_2_5_) );
  inv01 U6338 ( .Y(n7809), .A(r1_2_6_) );
  inv01 U6339 ( .Y(n7818), .A(r1_2_10_) );
  inv01 U6340 ( .Y(n7821), .A(r1_2_11_) );
  inv01 U6341 ( .Y(n7824), .A(r1_2_12_) );
  inv01 U6342 ( .Y(n7833), .A(r1_2_16_) );
  inv01 U6343 ( .Y(n7836), .A(r1_2_17_) );
  inv01 U6344 ( .Y(n7839), .A(r1_2_18_) );
  inv01 U6345 ( .Y(n7846), .A(r1_2_21_) );
  inv01 U6346 ( .Y(n7849), .A(r1_2_22_) );
  inv01 U6347 ( .Y(n7852), .A(r1_2_23_) );
  inv01 U6348 ( .Y(n7855), .A(r1_2_24_) );
  inv01 U6349 ( .Y(n7864), .A(r1_2_28_) );
  inv01 U6350 ( .Y(n7867), .A(r1_2_29_) );
  inv01 U6351 ( .Y(n7876), .A(r1_2_33_) );
  inv01 U6352 ( .Y(n7879), .A(r1_2_34_) );
  inv01 U6353 ( .Y(n7882), .A(r1_2_35_) );
  inv01 U6354 ( .Y(n7885), .A(r1_2_36_) );
  inv01 U6355 ( .Y(n7894), .A(r1_2_40_) );
  inv01 U6356 ( .Y(n7897), .A(r1_2_41_) );
  inv01 U6357 ( .Y(n7906), .A(r1_2_45_) );
  inv01 U6358 ( .Y(n7909), .A(r1_2_46_) );
  inv01 U6359 ( .Y(n7912), .A(r1_2_47_) );
  inv01 U6360 ( .Y(n7915), .A(r1_2_48_) );
  inv01 U6361 ( .Y(n7922), .A(r1_2_51_) );
  inv01 U6362 ( .Y(n7925), .A(r1_0_) );
  inv01 U6363 ( .Y(n7928), .A(r1_1_) );
  inv01 U6364 ( .Y(n7931), .A(r1_2_) );
  inv01 U6365 ( .Y(n7934), .A(r1_3_) );
  inv01 U6366 ( .Y(n7937), .A(r1_4_) );
  inv01 U6367 ( .Y(n7940), .A(r1_5_) );
  inv01 U6368 ( .Y(n7943), .A(r1_6_) );
  inv01 U6369 ( .Y(n7946), .A(r1_7_) );
  inv01 U6370 ( .Y(n7949), .A(r1_8_) );
  inv01 U6371 ( .Y(n7952), .A(r1_9_) );
  inv01 U6372 ( .Y(n7955), .A(r1_10_) );
  inv01 U6373 ( .Y(n7958), .A(r1_11_) );
  inv01 U6374 ( .Y(n7961), .A(r1_12_) );
  inv01 U6375 ( .Y(n7964), .A(r1_13_) );
  inv01 U6376 ( .Y(n7967), .A(r1_14_) );
  inv01 U6377 ( .Y(n7970), .A(r1_15_) );
  inv01 U6378 ( .Y(n7973), .A(r1_16_) );
  inv01 U6379 ( .Y(n7976), .A(r1_17_) );
  inv01 U6380 ( .Y(n7979), .A(r1_18_) );
  inv01 U6381 ( .Y(n7982), .A(r1_19_) );
  inv01 U6382 ( .Y(n7985), .A(r1_20_) );
  inv01 U6383 ( .Y(n7988), .A(r1_21_) );
  inv01 U6384 ( .Y(n7991), .A(r1_22_) );
  inv01 U6385 ( .Y(n7994), .A(r1_23_) );
  inv01 U6386 ( .Y(n7997), .A(r1_24_) );
  inv01 U6387 ( .Y(n8000), .A(r1_25_) );
  nand02 U6388 ( .Y(n7791), .A0(n7428), .A1(n8001) );
  nand02 U6389 ( .Y(n7789), .A0(n____return912), .A1(n7428) );
  nand02 U6390 ( .Y(n7788), .A0(n6950), .A1(n7787) );
  inv01 U6391 ( .Y(n7792), .A(s_sum2b[0]) );
  inv01 U6392 ( .Y(n7790), .A(s_sum1b[0]) );
  inv01 U6393 ( .Y(n7795), .A(s_sum2b[1]) );
  inv01 U6394 ( .Y(n7794), .A(s_sum1b[1]) );
  inv01 U6395 ( .Y(n7797), .A(s_sum2b[2]) );
  inv01 U6396 ( .Y(n7796), .A(s_sum1b[2]) );
  inv01 U6397 ( .Y(n7800), .A(s_sum2b[3]) );
  inv01 U6398 ( .Y(n7799), .A(s_sum1b[3]) );
  inv01 U6399 ( .Y(n7803), .A(s_sum2b[4]) );
  inv01 U6400 ( .Y(n7802), .A(s_sum1b[4]) );
  inv01 U6401 ( .Y(n7805), .A(s_sum2b[5]) );
  inv01 U6402 ( .Y(n7804), .A(s_sum1b[5]) );
  inv01 U6403 ( .Y(n7808), .A(s_sum2b[6]) );
  inv01 U6404 ( .Y(n7807), .A(s_sum1b[6]) );
  inv01 U6405 ( .Y(n7811), .A(s_sum2b[7]) );
  inv01 U6406 ( .Y(n7810), .A(s_sum1b[7]) );
  inv01 U6407 ( .Y(n7813), .A(s_sum2b[8]) );
  inv01 U6408 ( .Y(n7812), .A(s_sum1b[8]) );
  inv01 U6409 ( .Y(n7815), .A(s_sum2b[9]) );
  inv01 U6410 ( .Y(n7814), .A(s_sum1b[9]) );
  inv01 U6411 ( .Y(n7817), .A(s_sum2b[10]) );
  inv01 U6412 ( .Y(n7816), .A(s_sum1b[10]) );
  inv01 U6413 ( .Y(n7820), .A(s_sum2b[11]) );
  inv01 U6414 ( .Y(n7819), .A(s_sum1b[11]) );
  inv01 U6415 ( .Y(n7823), .A(s_sum2b[12]) );
  inv01 U6416 ( .Y(n7822), .A(s_sum1b[12]) );
  inv01 U6417 ( .Y(n7826), .A(s_sum2b[13]) );
  inv01 U6418 ( .Y(n7825), .A(s_sum1b[13]) );
  inv01 U6419 ( .Y(n7828), .A(s_sum2b[14]) );
  inv01 U6420 ( .Y(n7827), .A(s_sum1b[14]) );
  inv01 U6421 ( .Y(n7830), .A(s_sum2b[15]) );
  inv01 U6422 ( .Y(n7829), .A(s_sum1b[15]) );
  inv01 U6423 ( .Y(n7832), .A(s_sum2b[16]) );
  inv01 U6424 ( .Y(n7831), .A(s_sum1b[16]) );
  inv01 U6425 ( .Y(n7835), .A(s_sum2b[17]) );
  inv01 U6426 ( .Y(n7834), .A(s_sum1b[17]) );
  inv01 U6427 ( .Y(n7838), .A(s_sum2b[18]) );
  inv01 U6428 ( .Y(n7837), .A(s_sum1b[18]) );
  inv01 U6429 ( .Y(n7841), .A(s_sum2b[19]) );
  inv01 U6430 ( .Y(n7840), .A(s_sum1b[19]) );
  inv01 U6431 ( .Y(n7843), .A(s_sum2b[20]) );
  inv01 U6432 ( .Y(n7842), .A(s_sum1b[20]) );
  inv01 U6433 ( .Y(n7845), .A(s_sum2b[21]) );
  inv01 U6434 ( .Y(n7844), .A(s_sum1b[21]) );
  inv01 U6435 ( .Y(n7848), .A(s_sum2b[22]) );
  inv01 U6436 ( .Y(n7847), .A(s_sum1b[22]) );
  inv01 U6437 ( .Y(n7851), .A(s_sum2b[23]) );
  inv01 U6438 ( .Y(n7850), .A(s_sum1b[23]) );
  inv01 U6439 ( .Y(n7854), .A(s_sum2b[24]) );
  inv01 U6440 ( .Y(n7853), .A(s_sum1b[24]) );
  inv01 U6441 ( .Y(n7857), .A(s_sum2b[25]) );
  inv01 U6442 ( .Y(n7856), .A(s_sum1b[25]) );
  inv01 U6443 ( .Y(n7859), .A(s_sum2b[26]) );
  inv01 U6444 ( .Y(n7858), .A(s_sum1b[26]) );
  inv01 U6445 ( .Y(n7861), .A(s_sum2b[27]) );
  inv01 U6446 ( .Y(n7860), .A(s_sum1b[27]) );
  inv01 U6447 ( .Y(n7863), .A(s_sum2b[28]) );
  inv01 U6448 ( .Y(n7862), .A(s_sum1b[28]) );
  inv01 U6449 ( .Y(n7866), .A(s_sum2b[29]) );
  inv01 U6450 ( .Y(n7865), .A(s_sum1b[29]) );
  inv01 U6451 ( .Y(n7869), .A(s_sum2b[30]) );
  inv01 U6452 ( .Y(n7868), .A(s_sum1b[30]) );
  inv01 U6453 ( .Y(n7871), .A(s_sum2b[31]) );
  inv01 U6454 ( .Y(n7870), .A(s_sum1b[31]) );
  inv01 U6455 ( .Y(n7873), .A(s_sum2b[32]) );
  inv01 U6456 ( .Y(n7872), .A(s_sum1b[32]) );
  inv01 U6457 ( .Y(n7875), .A(s_sum2b[33]) );
  inv01 U6458 ( .Y(n7874), .A(s_sum1b[33]) );
  inv01 U6459 ( .Y(n7878), .A(s_sum2b[34]) );
  inv01 U6460 ( .Y(n7877), .A(s_sum1b[34]) );
  inv01 U6461 ( .Y(n7881), .A(s_sum2b[35]) );
  inv01 U6462 ( .Y(n7880), .A(s_sum1b[35]) );
  inv01 U6463 ( .Y(n7884), .A(s_sum2b[36]) );
  inv01 U6464 ( .Y(n7883), .A(s_sum1b[36]) );
  inv01 U6465 ( .Y(n7887), .A(s_sum2b[37]) );
  inv01 U6466 ( .Y(n7886), .A(s_sum1b[37]) );
  inv01 U6467 ( .Y(n7889), .A(s_sum2b[38]) );
  inv01 U6468 ( .Y(n7888), .A(s_sum1b[38]) );
  inv01 U6469 ( .Y(n7891), .A(s_sum2b[39]) );
  inv01 U6470 ( .Y(n7890), .A(s_sum1b[39]) );
  inv01 U6471 ( .Y(n7893), .A(s_sum2b[40]) );
  inv01 U6472 ( .Y(n7892), .A(s_sum1b[40]) );
  inv01 U6473 ( .Y(n7896), .A(s_sum2b[41]) );
  inv01 U6474 ( .Y(n7895), .A(s_sum1b[41]) );
  inv01 U6475 ( .Y(n7899), .A(s_sum2b[42]) );
  inv01 U6476 ( .Y(n7898), .A(s_sum1b[42]) );
  inv01 U6477 ( .Y(n7901), .A(s_sum2b[43]) );
  inv01 U6478 ( .Y(n7900), .A(s_sum1b[43]) );
  inv01 U6479 ( .Y(n7903), .A(s_sum2b[44]) );
  inv01 U6480 ( .Y(n7902), .A(s_sum1b[44]) );
  inv01 U6481 ( .Y(n7905), .A(s_sum2b[45]) );
  inv01 U6482 ( .Y(n7904), .A(s_sum1b[45]) );
  inv01 U6483 ( .Y(n7908), .A(s_sum2b[46]) );
  inv01 U6484 ( .Y(n7907), .A(s_sum1b[46]) );
  inv01 U6485 ( .Y(n7911), .A(s_sum2b[47]) );
  inv01 U6486 ( .Y(n7910), .A(s_sum1b[47]) );
  inv01 U6487 ( .Y(n7914), .A(s_sum2b[48]) );
  inv01 U6488 ( .Y(n7913), .A(s_sum1b[48]) );
  inv01 U6489 ( .Y(n7917), .A(s_sum2b[49]) );
  inv01 U6490 ( .Y(n7916), .A(s_sum1b[49]) );
  inv01 U6491 ( .Y(n7919), .A(s_sum2b[50]) );
  inv01 U6492 ( .Y(n7918), .A(s_sum1b[50]) );
  inv01 U6493 ( .Y(n7921), .A(s_sum2b[51]) );
  inv01 U6494 ( .Y(n7920), .A(s_sum1b[51]) );
  inv01 U6495 ( .Y(n7924), .A(s_sum2a_0_) );
  inv01 U6496 ( .Y(n7923), .A(s_sum1a_0_) );
  inv01 U6497 ( .Y(n7927), .A(s_sum2a_1_) );
  inv01 U6498 ( .Y(n7926), .A(s_sum1a_1_) );
  inv01 U6499 ( .Y(n7930), .A(s_sum2a_2_) );
  inv01 U6500 ( .Y(n7929), .A(s_sum1a_2_) );
  inv01 U6501 ( .Y(n7933), .A(s_sum2a_3_) );
  inv01 U6502 ( .Y(n7932), .A(s_sum1a_3_) );
  inv01 U6503 ( .Y(n7936), .A(s_sum2a_4_) );
  inv01 U6504 ( .Y(n7935), .A(s_sum1a_4_) );
  inv01 U6505 ( .Y(n7939), .A(s_sum2a_5_) );
  inv01 U6506 ( .Y(n7938), .A(s_sum1a_5_) );
  inv01 U6507 ( .Y(n7942), .A(s_sum2a_6_) );
  inv01 U6508 ( .Y(n7941), .A(s_sum1a_6_) );
  inv01 U6509 ( .Y(n7945), .A(s_sum2a_7_) );
  inv01 U6510 ( .Y(n7944), .A(s_sum1a_7_) );
  inv01 U6511 ( .Y(n7948), .A(s_sum2a_8_) );
  inv01 U6512 ( .Y(n7947), .A(s_sum1a_8_) );
  inv01 U6513 ( .Y(n7951), .A(s_sum2a_9_) );
  inv01 U6514 ( .Y(n7950), .A(s_sum1a_9_) );
  inv01 U6515 ( .Y(n7954), .A(s_sum2a_10_) );
  inv01 U6516 ( .Y(n7953), .A(s_sum1a_10_) );
  inv01 U6517 ( .Y(n7957), .A(s_sum2a_11_) );
  inv01 U6518 ( .Y(n7956), .A(s_sum1a_11_) );
  inv01 U6519 ( .Y(n7960), .A(s_sum2a_12_) );
  inv01 U6520 ( .Y(n7959), .A(s_sum1a_12_) );
  inv01 U6521 ( .Y(n7963), .A(s_sum2a_13_) );
  inv01 U6522 ( .Y(n7962), .A(s_sum1a_13_) );
  inv01 U6523 ( .Y(n7966), .A(s_sum2a_14_) );
  inv01 U6524 ( .Y(n7965), .A(s_sum1a_14_) );
  inv01 U6525 ( .Y(n7969), .A(s_sum2a_15_) );
  inv01 U6526 ( .Y(n7968), .A(s_sum1a_15_) );
  inv01 U6527 ( .Y(n7972), .A(s_sum2a_16_) );
  inv01 U6528 ( .Y(n7971), .A(s_sum1a_16_) );
  inv01 U6529 ( .Y(n7975), .A(s_sum2a_17_) );
  inv01 U6530 ( .Y(n7974), .A(s_sum1a_17_) );
  inv01 U6531 ( .Y(n7978), .A(s_sum2a_18_) );
  inv01 U6532 ( .Y(n7977), .A(s_sum1a_18_) );
  inv01 U6533 ( .Y(n7981), .A(s_sum2a_19_) );
  inv01 U6534 ( .Y(n7980), .A(s_sum1a_19_) );
  inv01 U6535 ( .Y(n7984), .A(s_sum2a_20_) );
  inv01 U6536 ( .Y(n7983), .A(s_sum1a_20_) );
  inv01 U6537 ( .Y(n7987), .A(s_sum2a_21_) );
  inv01 U6538 ( .Y(n7986), .A(s_sum1a_21_) );
  inv01 U6539 ( .Y(n7990), .A(s_sum2a_22_) );
  inv01 U6540 ( .Y(n7989), .A(s_sum1a_22_) );
  inv01 U6541 ( .Y(n7993), .A(s_sum2a_23_) );
  inv01 U6542 ( .Y(n7992), .A(s_sum1a_23_) );
  inv01 U6543 ( .Y(n7996), .A(s_sum2a_24_) );
  inv01 U6544 ( .Y(n7995), .A(s_sum1a_24_) );
  nand03 U6545 ( .Y(n8003), .A0(n8001), .A1(n7787), .A2(n7433) );
  inv01 U6546 ( .Y(n8001), .A(n____return912) );
  inv01 U6547 ( .Y(n7999), .A(s_sum2a_25_) );
  nand03 U6548 ( .Y(n8002), .A0(n7431), .A1(n7787), .A2(n____return912) );
  inv01 U6549 ( .Y(n7998), .A(s_sum1a_25_) );
  inv01 U6550 ( .Y(n7455), .A(r0_49_) );
  and02 U6551 ( .Y(n2843), .A0(r0_50_), .A1(n7363) );
  and02 U6552 ( .Y(n2842), .A0(r0_51_), .A1(n7361) );
  nand02 U6553 ( .Y(n2841), .A0(n8004), .A1(n6827) );
  mux21 U6554 ( .Y(n8004), .A0(s_count_4_), .A1(sum181_4_), .S0(s_state) );
  nand02 U6555 ( .Y(n2840), .A0(n8005), .A1(n6827) );
  mux21 U6556 ( .Y(n8005), .A0(s_count_3_), .A1(sum181_3_), .S0(s_state) );
  ao32 U6557 ( .Y(n2839), .A0(s_state), .A1(n6952), .A2(sum181_2_), .B0(
        s_count_2_), .B1(n7363) );
  nand02 U6558 ( .Y(n2838), .A0(n8006), .A1(n6827) );
  mux21 U6559 ( .Y(n8006), .A0(s_count_1_), .A1(sum181_1_), .S0(s_state) );
  ao32 U6560 ( .Y(n2837), .A0(s_state), .A1(n6952), .A2(sum181_0_), .B0(
        s_count_0_), .B1(n7362) );
  or03 U6561 ( .Y(n8007), .A0(s_count_2_), .A1(s_count_4_), .A2(s_count_3_) );
  or02 U6562 ( .Y(c222_4_), .A0(ARG260_4_), .A1(n7419) );
  or02 U6563 ( .Y(c222_3_), .A0(ARG260_3_), .A1(n7421) );
  and02 U6564 ( .Y(c222_2_), .A0(ARG260_2_), .A1(n7787) );
  or02 U6565 ( .Y(c222_1_), .A0(ARG260_1_), .A1(n7421) );
  and02 U6566 ( .Y(c222_0_), .A0(ARG260_0_), .A1(n7787) );
  nand02 U6567 ( .Y(b206_25_), .A0(n7787), .A1(n1906) );
  sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_inc_52_0 add_0_root_add_199_plus_plus ( .A({
        n____return1344_51_, n____return1344_50_, n1346_49_, 
        n____return1344_48_, n____return1344_47_, n____return1344_46_, 
        n____return1344_45_, n____return1344_44_, n____return1344_43_, 
        n____return1344_42_, n____return1344_41_, n____return1344_40_, 
        n____return1344_39_, n____return1344_38_, n____return1344_37_, 
        n____return1344_36_, n____return1344_35_, n____return1344_34_, 
        n____return1344_33_, n____return1344_32_, n____return1344_31_, 
        n____return1344_30_, n____return1344_29_, n____return1344_28_, 
        n____return1344_27_, n____return1344_26_, n____return1344_25_, 
        n____return1344_24_, n____return1344_23_, n____return1344_22_, 
        n____return1344_21_, n____return1344_20_, n____return1344_19_, 
        n____return1344_18_, n____return1344_17_, n____return1344_16_, 
        n____return1344_15_, n____return1344_14_, n____return1344_13_, 
        n____return1344_12_, n____return1344_11_, n____return1344_10_, 
        n____return1344_9_, n____return1344_8_, n____return1344_7_, 
        n____return1344_6_, n____return1344_5_, n____return1344_4_, 
        n____return1344_3_, n____return1344_2_, n____return1344_1_, 
        n____return1344_0_}), .SUM({n1384_51_, n____return1382_50_, n1384_49_, 
        n____return1382_48_, n____return1382_47_, n____return1382_46_, 
        n____return1382_45_, n____return1382_44_, n____return1382_43_, 
        n____return1382_42_, n____return1382_41_, n____return1382_40_, 
        n____return1382_39_, n____return1382_38_, n____return1382_37_, 
        n____return1382_36_, n____return1382_35_, n____return1382_34_, 
        n____return1382_33_, n____return1382_32_, n____return1382_31_, 
        n____return1382_30_, n____return1382_29_, n____return1382_28_, 
        n____return1382_27_, n____return1382_26_, n____return1382_25_, 
        n____return1382_24_, n____return1382_23_, n____return1382_22_, 
        n____return1382_21_, n____return1382_20_, n____return1382_19_, 
        n____return1382_18_, n____return1382_17_, n____return1382_16_, 
        n____return1382_15_, n____return1382_14_, n____return1382_13_, 
        n____return1382_12_, n____return1382_11_, n____return1382_10_, 
        n____return1382_9_, n____return1382_8_, n____return1382_7_, 
        n____return1382_6_, n____return1382_5_, n____return1382_4_, 
        n____return1382_3_, n____return1382_2_, n____return1382_1_, 
        n____return1382_0_}) );
  sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_sub_52_1 sub_1_root_add_199_plus_plus ( .A({
        n6948, r1_2_50_, r1_2_49_, n6891, n6845, n6883, n6831, r1_2_44_, 
        r1_2_43_, r1_2_42_, n6843, n6873, r1_2_39_, r1_2_38_, r1_2_37_, n6893, 
        n6835, n6879, n6849, r1_2_32_, r1_2_31_, r1_2_30_, n6855, n6875, 
        r1_2_27_, r1_2_26_, r1_2_25_, n6887, n6847, n6869, n6837, r1_2_20_, 
        r1_2_19_, n6881, n6851, n6877, r1_2_15_, r1_2_14_, r1_2_13_, n6889, 
        n6839, n6853, r1_2_9_, r1_2_8_, r1_2_7_, n6885, n6833, r1_2_4_, n6841, 
        n6871, r1_2_1_, r1_2_0_}), .B({r1_50_, r1_49_, r1_48_, r1_47_, r1_46_, 
        r1_45_, r1_44_, r1_43_, r1_42_, r1_41_, r1_40_, r1_39_, r1_38_, r1_37_, 
        r1_36_, r1_35_, r1_34_, r1_33_, r1_32_, r1_31_, r1_30_, r1_29_, r1_28_, 
        r1_27_, r1_26_, r1_25_, r1_24_, r1_23_, r1_22_, r1_21_, r1_20_, r1_19_, 
        r1_18_, r1_17_, r1_16_, r1_15_, r1_14_, r1_13_, r1_12_, r1_11_, r1_10_, 
        r1_9_, r1_8_, r1_7_, r1_6_, r1_5_, r1_4_, r1_3_, r1_2_, r1_1_, r1_0_, 
        1'b0}), .CI(1'b0), .DIFF({n____return1344_51_, n____return1344_50_, 
        n1346_49_, n____return1344_48_, n____return1344_47_, 
        n____return1344_46_, n____return1344_45_, n____return1344_44_, 
        n____return1344_43_, n____return1344_42_, n____return1344_41_, 
        n____return1344_40_, n____return1344_39_, n____return1344_38_, 
        n____return1344_37_, n____return1344_36_, n____return1344_35_, 
        n____return1344_34_, n____return1344_33_, n____return1344_32_, 
        n____return1344_31_, n____return1344_30_, n____return1344_29_, 
        n____return1344_28_, n____return1344_27_, n____return1344_26_, 
        n____return1344_25_, n____return1344_24_, n____return1344_23_, 
        n____return1344_22_, n____return1344_21_, n____return1344_20_, 
        n____return1344_19_, n____return1344_18_, n____return1344_17_, 
        n____return1344_16_, n____return1344_15_, n____return1344_14_, 
        n____return1344_13_, n____return1344_12_, n____return1344_11_, 
        n____return1344_10_, n____return1344_9_, n____return1344_8_, 
        n____return1344_7_, n____return1344_6_, n____return1344_5_, 
        n____return1344_4_, n____return1344_3_, n____return1344_2_, 
        n____return1344_1_, n____return1344_0_}) );
  sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_dec_26_0 sub_185_sub_169_minus ( .A({r1_25_, 
        r1_24_, r1_23_, r1_22_, r1_21_, r1_20_, r1_19_, r1_18_, r1_17_, r1_16_, 
        r1_15_, r1_14_, r1_13_, r1_12_, r1_11_, r1_10_, r1_9_, r1_8_, r1_7_, 
        r1_6_, r1_5_, r1_4_, r1_3_, r1_2_, r1_1_, n4391}), .SUM({ARG1118_25_, 
        ARG1118_24_, ARG1118_23_, ARG1118_22_, ARG1118_21_, ARG1118_20_, 
        ARG1118_19_, ARG1118_18_, ARG1118_17_, ARG1118_16_, ARG1118_15_, 
        ARG1118_14_, ARG1118_13_, ARG1118_12_, ARG1118_11_, ARG1118_10_, 
        ARG1118_9_, ARG1118_8_, ARG1118_7_, ARG1118_6_, ARG1118_5_, ARG1118_4_, 
        ARG1118_3_, ARG1118_2_, ARG1118_1_, ARG1118_0_}) );
  sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_cmp2_52_1 gt_184_gt_gt ( .A({n6782, n6276, 
        s_rad_i_49_, s_rad_i_48_, s_rad_i_47_, s_rad_i_46_, s_rad_i_45_, n6267, 
        s_rad_i_43_, n6294, s_rad_i_41_, s_rad_i_40_, s_rad_i_39_, n6273, 
        s_rad_i_37_, s_rad_i_36_, s_rad_i_35_, s_rad_i_34_, s_rad_i_33_, n6282, 
        s_rad_i_31_, s_rad_i_30_, s_rad_i_29_, s_rad_i_28_, s_rad_i_27_, n6290, 
        s_rad_i_25_, n6261, s_rad_i_23_, s_rad_i_22_, s_rad_i_21_, n6279, 
        s_rad_i_19_, s_rad_i_18_, s_rad_i_17_, s_rad_i_16_, s_rad_i_15_, n6287, 
        s_rad_i_13_, n6257, s_rad_i_11_, s_rad_i_10_, n6270, n6256, s_rad_i_7_, 
        s_rad_i_6_, s_rad_i_5_, n6285, s_rad_i_3_, s_rad_i_2_, s_rad_i_1_, 
        s_rad_i_0_}), .B({n6948, n6132, n6164, n6891, n6845, n6883, n6831, 
        n6246, n6172, n6240, n6843, n6873, n6180, n6236, n6170, n6893, n6835, 
        n6879, n6849, n6238, n6184, n6250, n6855, n6875, n6176, n6234, n6182, 
        n6887, n6847, n6869, n6837, n6244, n6168, n6881, n6851, n6877, n6174, 
        n6242, n6166, n6889, n6839, n6853, n6232, n6252, n6178, n6885, n6833, 
        n6248, n6841, n6871, r1_2_1_, r1_2_0_}), .LEQ(1'b0), .TC(1'b0), 
        .LT_LE(n____return1071) );
  sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_cmp2_52_0 gt_163_gt_gt ( .A({n6783, n6275, 
        s_rad_i_49_, s_rad_i_48_, s_rad_i_47_, s_rad_i_46_, s_rad_i_45_, n6266, 
        s_rad_i_43_, n6293, s_rad_i_41_, s_rad_i_40_, s_rad_i_39_, n6272, 
        s_rad_i_37_, s_rad_i_36_, s_rad_i_35_, s_rad_i_34_, s_rad_i_33_, n6281, 
        s_rad_i_31_, s_rad_i_30_, s_rad_i_29_, s_rad_i_28_, s_rad_i_27_, n6291, 
        s_rad_i_25_, n6264, s_rad_i_23_, s_rad_i_22_, s_rad_i_21_, n6278, 
        s_rad_i_19_, s_rad_i_18_, s_rad_i_17_, s_rad_i_16_, s_rad_i_15_, n6288, 
        s_rad_i_13_, n6260, s_rad_i_11_, s_rad_i_10_, n6269, n6253, s_rad_i_7_, 
        s_rad_i_6_, s_rad_i_5_, n6284, s_rad_i_3_, s_rad_i_2_, s_rad_i_1_, 
        s_rad_i_0_}), .B({r0_2_51_, r0_2_50_, r0_2_49_, r0_2_48_, r0_2_47_, 
        r0_2_46_, r0_2_45_, r0_2_44_, r0_2_43_, r0_2_42_, r0_2_41_, r0_2_40_, 
        r0_2_39_, r0_2_38_, r0_2_37_, r0_2_36_, r0_2_35_, r0_2_34_, r0_2_33_, 
        r0_2_32_, r0_2_31_, r0_2_30_, r0_2_29_, r0_2_28_, r0_2_27_, r0_2_26_, 
        r0_2_25_, r0_2_24_, r0_2_23_, r0_2_22_, r0_2_21_, r0_2_20_, r0_2_19_, 
        r0_2_18_, r0_2_17_, r0_2_16_, r0_2_15_, r0_2_14_, r0_2_13_, r0_2_12_, 
        r0_2_11_, r0_2_10_, r0_2_9_, r0_2_8_, r0_2_7_, r0_2_6_, r0_2_5_, 
        r0_2_4_, r0_2_3_, r0_2_2_, r0_2_1_, r0_2_0_}), .LEQ(1'b0), .TC(1'b0), 
        .LT_LE(n____return912) );
  sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_add_52_1 add_151_plus_plus ( .A({s_op1_51_, 
        s_op1_50_, s_op1_49_, s_op1_48_, s_op1_47_, s_op1_46_, s_op1_45_, 
        s_op1_44_, s_op1_43_, s_op1_42_, s_op1_41_, s_op1_40_, s_op1_39_, 
        s_op1_38_, s_op1_37_, s_op1_36_, s_op1_35_, s_op1_34_, s_op1_33_, 
        s_op1_32_, s_op1_31_, s_op1_30_, s_op1_29_, s_op1_28_, s_op1_27_, 
        s_op1_26_, s_op1_25_, s_op1_24_, s_op1_23_, s_op1_22_, s_op1_21_, 
        s_op1_20_, s_op1_19_, s_op1_18_, s_op1_17_, s_op1_16_, s_op1_15_, 
        s_op1_14_, s_op1_13_, s_op1_12_, s_op1_11_, s_op1_10_, s_op1_9_, 
        s_op1_8_, s_op1_7_, s_op1_6_, s_op1_5_, s_op1_4_, s_op1_3_, s_op1_2_, 
        s_op1_1_, s_op1_0_}), .B({s_op2_51_, result407_50_, s_op2_49_, 
        s_op2_48_, s_op2_47_, s_op2_46_, s_op2_45_, s_op2_44_, s_op2_43_, 
        s_op2_42_, s_op2_41_, s_op2_40_, s_op2_39_, s_op2_38_, s_op2_37_, 
        s_op2_36_, n7104, n7093, n7117, n7108, n7119, n7102, n7095, n7115, 
        n7099, n7097, n7113, n7111, s_op2_23_, s_op2_22_, s_op2_21_, n7106, 
        s_op2_19_, s_op2_18_, s_op2_17_, s_op2_16_, n7334, n7336, n7332, n7345, 
        n7347, n7339, n7343, n7341, s_op2_7_, n6955, n6961, s_op2_4_, s_op2_3_, 
        n7324, n7326, n7329}), .CI(1'b0), .SUM(s_sum2b) );
  sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_sub_52_0 sub_150_minus_minus ( .A({s_op1_51_, 
        s_op1_50_, s_op1_49_, s_op1_48_, s_op1_47_, s_op1_46_, s_op1_45_, 
        s_op1_44_, s_op1_43_, s_op1_42_, s_op1_41_, s_op1_40_, s_op1_39_, 
        s_op1_38_, s_op1_37_, s_op1_36_, s_op1_35_, s_op1_34_, s_op1_33_, 
        s_op1_32_, s_op1_31_, s_op1_30_, s_op1_29_, s_op1_28_, s_op1_27_, 
        s_op1_26_, s_op1_25_, s_op1_24_, s_op1_23_, s_op1_22_, s_op1_21_, 
        s_op1_20_, s_op1_19_, s_op1_18_, s_op1_17_, s_op1_16_, s_op1_15_, 
        s_op1_14_, s_op1_13_, s_op1_12_, s_op1_11_, s_op1_10_, s_op1_9_, 
        s_op1_8_, s_op1_7_, s_op1_6_, s_op1_5_, s_op1_4_, s_op1_3_, s_op1_2_, 
        s_op1_1_, s_op1_0_}), .B({s_op2_51_, result407_50_, s_op2_49_, 
        s_op2_48_, s_op2_47_, s_op2_46_, s_op2_45_, s_op2_44_, s_op2_43_, 
        s_op2_42_, s_op2_41_, s_op2_40_, s_op2_39_, s_op2_38_, s_op2_37_, 
        s_op2_36_, n7104, n7092, n7117, n7108, n7119, n7101, n7095, n7115, 
        n7099, n7097, n7113, n7110, s_op2_23_, s_op2_22_, s_op2_21_, n7106, 
        s_op2_19_, s_op2_18_, s_op2_17_, s_op2_16_, n7334, n7336, n7332, n7345, 
        n7347, n7338, n7343, n7341, s_op2_7_, n6954, n6960, s_op2_4_, n7327, 
        n7324, n7326, n7330}), .CI(1'b0), .DIFF(s_sum1b) );
  sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_add_26_0 add_149_plus_plus ( .A({n7145, 
        n7122, n7167, n7165, n7211, n7208, n7205, n7200, n7206, n7201, n7204, 
        n7187, n7207, n7210, n7203, n7209, n7213, n7214, n7202, n7186, n7212, 
        n7125, n7123, n7121, n7164, n6906}), .B({b_25_, b_24_, b_23_, b_22_, 
        b_21_, b_20_, b_19_, b_18_, b_17_, b_16_, b_15_, b_14_, b_13_, b_12_, 
        b_11_, b_10_, b_9_, b_8_, b_7_, b_6_, b_5_, b_4_, b_3_, b_2_, b_1_, 
        b_0_}), .CI(1'b0), .SUM({s_sum2a_25_, s_sum2a_24_, s_sum2a_23_, 
        s_sum2a_22_, s_sum2a_21_, s_sum2a_20_, s_sum2a_19_, s_sum2a_18_, 
        s_sum2a_17_, s_sum2a_16_, s_sum2a_15_, s_sum2a_14_, s_sum2a_13_, 
        s_sum2a_12_, s_sum2a_11_, s_sum2a_10_, s_sum2a_9_, s_sum2a_8_, 
        s_sum2a_7_, s_sum2a_6_, s_sum2a_5_, s_sum2a_4_, s_sum2a_3_, s_sum2a_2_, 
        s_sum2a_1_, s_sum2a_0_}) );
  sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_sub_26_0 sub_148_minus_minus ( .A({n7145, 
        n7122, n7167, n7165, n7211, n7208, n7205, n7200, n7206, n7201, n7204, 
        n7187, n7207, n7210, n7203, n7209, n7213, n7214, n7202, n7186, n7212, 
        n7125, n7123, n7121, n7164, n6906}), .B({b_25_, b_24_, b_23_, b_22_, 
        b_21_, b_20_, b_19_, b_18_, b_17_, b_16_, b_15_, b_14_, b_13_, b_12_, 
        b_11_, b_10_, b_9_, b_8_, b_7_, b_6_, b_5_, b_4_, b_3_, b_2_, b_1_, 
        b_0_}), .CI(1'b0), .DIFF({s_sum1a_25_, s_sum1a_24_, s_sum1a_23_, 
        s_sum1a_22_, s_sum1a_21_, s_sum1a_20_, s_sum1a_19_, s_sum1a_18_, 
        s_sum1a_17_, s_sum1a_16_, s_sum1a_15_, s_sum1a_14_, s_sum1a_13_, 
        s_sum1a_12_, s_sum1a_11_, s_sum1a_10_, s_sum1a_9_, s_sum1a_8_, 
        s_sum1a_7_, s_sum1a_6_, s_sum1a_5_, s_sum1a_4_, s_sum1a_3_, s_sum1a_2_, 
        s_sum1a_1_, s_sum1a_0_}) );
  sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_add_52_0 add_146_plus_plus ( .A({r0_2_51_, 
        r0_2_50_, r0_2_49_, r0_2_48_, r0_2_47_, r0_2_46_, r0_2_45_, r0_2_44_, 
        r0_2_43_, r0_2_42_, r0_2_41_, r0_2_40_, r0_2_39_, r0_2_38_, r0_2_37_, 
        r0_2_36_, r0_2_35_, r0_2_34_, r0_2_33_, r0_2_32_, r0_2_31_, r0_2_30_, 
        r0_2_29_, r0_2_28_, r0_2_27_, r0_2_26_, r0_2_25_, r0_2_24_, r0_2_23_, 
        r0_2_22_, r0_2_21_, r0_2_20_, r0_2_19_, r0_2_18_, r0_2_17_, r0_2_16_, 
        r0_2_15_, r0_2_14_, r0_2_13_, r0_2_12_, r0_2_11_, r0_2_10_, r0_2_9_, 
        r0_2_8_, r0_2_7_, r0_2_6_, r0_2_5_, r0_2_4_, r0_2_3_, r0_2_2_, r0_2_1_, 
        r0_2_0_}), .B(b_2), .CI(1'b0), .SUM({s_op1_51_, s_op1_50_, s_op1_49_, 
        s_op1_48_, s_op1_47_, s_op1_46_, s_op1_45_, s_op1_44_, s_op1_43_, 
        s_op1_42_, s_op1_41_, s_op1_40_, s_op1_39_, s_op1_38_, s_op1_37_, 
        s_op1_36_, s_op1_35_, s_op1_34_, s_op1_33_, s_op1_32_, s_op1_31_, 
        s_op1_30_, s_op1_29_, s_op1_28_, s_op1_27_, s_op1_26_, s_op1_25_, 
        s_op1_24_, s_op1_23_, s_op1_22_, s_op1_21_, s_op1_20_, s_op1_19_, 
        s_op1_18_, s_op1_17_, s_op1_16_, s_op1_15_, s_op1_14_, s_op1_13_, 
        s_op1_12_, s_op1_11_, s_op1_10_, s_op1_9_, s_op1_8_, s_op1_7_, 
        s_op1_6_, s_op1_5_, s_op1_4_, s_op1_3_, s_op1_2_, s_op1_1_, s_op1_0_})
         );
  sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_dec_5_1 sub_139_sub_169_minus ( .A({n7377, 
        n4177, c_2_, n6946, n6576}), .SUM({ARG260_4_, ARG260_3_, ARG260_2_, 
        ARG260_1_, ARG260_0_}) );
  sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_dec_5_0 sub_121 ( .A({s_count_4_, s_count_3_, 
        s_count_2_, s_count_1_, s_count_0_}), .SUM({sum181_4_, sum181_3_, 
        sum181_2_, sum181_1_, sum181_0_}) );
endmodule


module fpu_DW01_inc_32_0 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   carry_31_, carry_30_, carry_29_, carry_28_, carry_27_, carry_26_,
         carry_25_, carry_24_, carry_23_, carry_22_, carry_21_, carry_20_,
         carry_19_, carry_18_, carry_17_, carry_16_, carry_15_, carry_14_,
         carry_13_, carry_12_, carry_11_, carry_10_, carry_9_, carry_8_,
         carry_7_, carry_6_, carry_5_, carry_4_, carry_3_, carry_2_;

  inv01 U5 ( .Y(SUM[0]), .A(A[0]) );
  xor2 U6 ( .Y(SUM[31]), .A0(carry_31_), .A1(A[31]) );
  hadd1 U1_1_1 ( .S(SUM[1]), .CO(carry_2_), .A(A[1]), .B(A[0]) );
  hadd1 U1_1_2 ( .S(SUM[2]), .CO(carry_3_), .A(A[2]), .B(carry_2_) );
  hadd1 U1_1_3 ( .S(SUM[3]), .CO(carry_4_), .A(A[3]), .B(carry_3_) );
  hadd1 U1_1_4 ( .S(SUM[4]), .CO(carry_5_), .A(A[4]), .B(carry_4_) );
  hadd1 U1_1_5 ( .S(SUM[5]), .CO(carry_6_), .A(A[5]), .B(carry_5_) );
  hadd1 U1_1_6 ( .S(SUM[6]), .CO(carry_7_), .A(A[6]), .B(carry_6_) );
  hadd1 U1_1_7 ( .S(SUM[7]), .CO(carry_8_), .A(A[7]), .B(carry_7_) );
  hadd1 U1_1_8 ( .S(SUM[8]), .CO(carry_9_), .A(A[8]), .B(carry_8_) );
  hadd1 U1_1_9 ( .S(SUM[9]), .CO(carry_10_), .A(A[9]), .B(carry_9_) );
  hadd1 U1_1_10 ( .S(SUM[10]), .CO(carry_11_), .A(A[10]), .B(carry_10_) );
  hadd1 U1_1_11 ( .S(SUM[11]), .CO(carry_12_), .A(A[11]), .B(carry_11_) );
  hadd1 U1_1_12 ( .S(SUM[12]), .CO(carry_13_), .A(A[12]), .B(carry_12_) );
  hadd1 U1_1_13 ( .S(SUM[13]), .CO(carry_14_), .A(A[13]), .B(carry_13_) );
  hadd1 U1_1_14 ( .S(SUM[14]), .CO(carry_15_), .A(A[14]), .B(carry_14_) );
  hadd1 U1_1_15 ( .S(SUM[15]), .CO(carry_16_), .A(A[15]), .B(carry_15_) );
  hadd1 U1_1_16 ( .S(SUM[16]), .CO(carry_17_), .A(A[16]), .B(carry_16_) );
  hadd1 U1_1_17 ( .S(SUM[17]), .CO(carry_18_), .A(A[17]), .B(carry_17_) );
  hadd1 U1_1_18 ( .S(SUM[18]), .CO(carry_19_), .A(A[18]), .B(carry_18_) );
  hadd1 U1_1_19 ( .S(SUM[19]), .CO(carry_20_), .A(A[19]), .B(carry_19_) );
  hadd1 U1_1_20 ( .S(SUM[20]), .CO(carry_21_), .A(A[20]), .B(carry_20_) );
  hadd1 U1_1_21 ( .S(SUM[21]), .CO(carry_22_), .A(A[21]), .B(carry_21_) );
  hadd1 U1_1_22 ( .S(SUM[22]), .CO(carry_23_), .A(A[22]), .B(carry_22_) );
  hadd1 U1_1_23 ( .S(SUM[23]), .CO(carry_24_), .A(A[23]), .B(carry_23_) );
  hadd1 U1_1_24 ( .S(SUM[24]), .CO(carry_25_), .A(A[24]), .B(carry_24_) );
  hadd1 U1_1_25 ( .S(SUM[25]), .CO(carry_26_), .A(A[25]), .B(carry_25_) );
  hadd1 U1_1_26 ( .S(SUM[26]), .CO(carry_27_), .A(A[26]), .B(carry_26_) );
  hadd1 U1_1_27 ( .S(SUM[27]), .CO(carry_28_), .A(A[27]), .B(carry_27_) );
  hadd1 U1_1_28 ( .S(SUM[28]), .CO(carry_29_), .A(A[28]), .B(carry_28_) );
  hadd1 U1_1_29 ( .S(SUM[29]), .CO(carry_30_), .A(A[29]), .B(carry_29_) );
  hadd1 U1_1_30 ( .S(SUM[30]), .CO(carry_31_), .A(A[30]), .B(carry_30_) );
endmodule


module fpu ( clk_i, opa_i, opb_i, fpu_op_i, rmode_i, output_o, start_i, 
        ready_o, ine_o, overflow_o, underflow_o, div_zero_o, inf_o, zero_o, 
        qnan_o, snan_o );
  input [31:0] opa_i;
  input [31:0] opb_i;
  input [2:0] fpu_op_i;
  input [1:0] rmode_i;
  output [31:0] output_o;
  input clk_i, start_i;
  output ready_o, ine_o, overflow_o, underflow_o, div_zero_o, inf_o, zero_o,
         qnan_o, snan_o;
  wire   s_fpu_op_i_0_, addsub_sign_o, postnorm_addsub_ine_o, mul_24_sign,
         post_norm_mul_ine, serial_div_sign, post_norm_div_ine, sqrt_ine_o,
         post_norm_sqrt_ine_o, s_output_o_31_, s_output_o_30_, s_output_o_29_,
         s_output_o_28_, s_output_o_27_, s_output_o_26_, s_output_o_25_,
         s_output_o_24_, s_output_o_22_, s_output_o_21_, s_output_o_20_,
         s_output_o_19_, s_output_o_18_, s_output_o_17_, s_output_o_16_,
         s_output_o_15_, s_output_o_14_, s_output_o_13_, s_output_o_12_,
         s_output_o_11_, s_output_o_10_, s_output_o_9_, s_output_o_8_,
         s_output_o_7_, s_output_o_6_, s_output_o_5_, s_output_o_4_,
         s_output_o_3_, s_output_o_2_, s_output_o_1_, s_output_o_0_, s_ine_o,
         s_div_zero_o, s_inf_o, s_zero_o, s_qnan_o, s_snan_o, s_output1_31_,
         s_output1_23_, s_output1_22_, s_output1_21_, s_output1_20_,
         s_output1_19_, s_output1_18_, s_output1_17_, s_output1_16_,
         s_output1_11_, s_output1_10_, s_output1_9_, s_output1_8_,
         s_output1_7_, s_output1_6_, s_output1_5_, s_output1_4_, s_output1_3_,
         s_output1_2_, s_output1_1_, s_output1_0_, serial_div_div_zero,
         s_state, s_state213, s_count_31_, s_count_30_, s_count_29_,
         s_count_28_, s_count_27_, s_count_26_, s_count_25_, s_count_24_,
         s_count_23_, s_count_22_, s_count_21_, s_count_20_, s_count_19_,
         s_count_18_, s_count_17_, s_count_16_, s_count_15_, s_count_14_,
         s_count_13_, s_count_12_, s_count_11_, s_count_10_, s_count_9_,
         s_count_8_, s_count_7_, s_count_6_, s_count_5_, s_count_4_,
         s_count_3_, s_count_2_, s_count_1_, s_count_0_, sum339_31_,
         sum339_30_, sum339_29_, sum339_28_, sum339_27_, sum339_26_,
         sum339_25_, sum339_24_, sum339_23_, sum339_22_, sum339_21_,
         sum339_20_, sum339_19_, sum339_18_, sum339_17_, sum339_16_,
         sum339_15_, sum339_14_, sum339_13_, sum339_12_, sum339_11_,
         sum339_10_, sum339_9_, sum339_8_, sum339_7_, sum339_6_, sum339_5_,
         sum339_4_, sum339_3_, sum339_2_, sum339_1_, sum339_0_,
         s_output1408_31_, s_output1408_30_, s_output1408_29_,
         s_output1408_28_, s_output1408_27_, s_output1408_26_,
         s_output1408_25_, s_output1408_24_, s_output1408_23_,
         s_output1408_22_, s_output1408_21_, s_output1408_20_,
         s_output1408_19_, s_output1408_18_, s_output1408_17_,
         s_output1408_16_, s_output1408_15_, s_output1408_14_,
         s_output1408_13_, s_output1408_12_, s_output1408_11_,
         s_output1408_10_, s_output1408_9_, s_output1408_8_, s_output1408_7_,
         s_output1408_6_, s_output1408_5_, s_output1408_4_, s_output1408_3_,
         s_output1408_2_, s_output1408_1_, s_output1408_0_, s_ine_o415, n650,
         n651, n652, n653, n654, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n682, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104;
  wire   [31:0] s_opa_i;
  wire   [31:0] s_opb_i;
  wire   [27:0] prenorm_addsub_fracta_28_o;
  wire   [27:0] prenorm_addsub_fractb_28_o;
  wire   [7:0] prenorm_addsub_exp_o;
  wire   [27:0] addsub_fract_o;
  wire   [1:0] s_rmode_i;
  wire   [31:0] postnorm_addsub_output_o;
  wire   [9:0] pre_norm_mul_exp_10;
  wire   [23:0] pre_norm_mul_fracta_24;
  wire   [23:0] pre_norm_mul_fractb_24;
  wire   [31:0] post_norm_mul_output;
  wire   [9:0] pre_norm_div_exp;
  wire   [49:0] pre_norm_div_dvdnd;
  wire   [26:0] pre_norm_div_dvsor;
  wire   [26:0] serial_div_qutnt;
  wire   [26:0] serial_div_rmndr;
  wire   [31:0] post_norm_div_output;
  wire   [51:0] pre_norm_sqrt_fracta_o;
  wire   [7:0] pre_norm_sqrt_exp_o;
  wire   [25:0] sqrt_sqr_o;
  wire   [31:0] post_norm_sqrt_output;
  wire   [47:0] mul_fract_48;

  pre_norm_addsub i_prenorm_addsub ( .clk_i(clk_i), .opa_i({s_opa_i[31], n1315, 
        n1311, n1310, n1314, n1309, n1316, n1312, n1303, s_opa_i[22:21], n1305, 
        n1300, s_opa_i[18], n1301, s_opa_i[16:15], n1272, s_opa_i[13], n1292, 
        s_opa_i[11], n1280, n1278, n1276, n1291, s_opa_i[6:2], n1293, n1302}), 
        .opb_i({n1233, s_opb_i[30:28], n1277, s_opb_i[26:24], n1258, 
        s_opb_i[22], n1236, s_opb_i[20], n1237, s_opb_i[18:17], n1245, n1255, 
        s_opb_i[14], n1227, n1226, n1225, n1240, n1231, n1228, n1230, 
        s_opb_i[6], n1247, n1242, n1229, n1243, s_opb_i[1], n1251}), 
        .fracta_28_o(prenorm_addsub_fracta_28_o), .fractb_28_o(
        prenorm_addsub_fractb_28_o), .exp_o(prenorm_addsub_exp_o) );
  addsub_28 i_addsub ( .clk_i(clk_i), .fpu_op_i(s_fpu_op_i_0_), .fracta_i(
        prenorm_addsub_fracta_28_o), .fractb_i(prenorm_addsub_fractb_28_o), 
        .signa_i(n1265), .signb_i(n1234), .fract_o(addsub_fract_o), .sign_o(
        addsub_sign_o) );
  post_norm_addsub i_postnorm_addsub ( .clk_i(clk_i), .opa_i({s_opa_i[31], 
        n1315, n1311, n1310, n1314, n1309, n1316, n1312, n1303, s_opa_i[22], 
        n1298, s_opa_i[20], n1300, s_opa_i[18], n1301, s_opa_i[16], n1290, 
        s_opa_i[14], n1285, s_opa_i[12:5], n1274, n1270, n1275, n1293, 
        s_opa_i[0]}), .opb_i({n1234, n1288, s_opb_i[29:23], n1222, n1236, 
        n1224, s_opb_i[19:18], n1248, s_opb_i[16], n1255, s_opb_i[14], n1227, 
        n1226, s_opb_i[11], n1240, n1231, n1228, n1230, n1257, s_opb_i[5], 
        n1242, n1229, s_opb_i[2:1], n1250}), .fract_28_i(addsub_fract_o), 
        .exp_i(prenorm_addsub_exp_o), .sign_i(addsub_sign_o), .fpu_op_i(
        s_fpu_op_i_0_), .rmode_i({n1219, s_rmode_i[0]}), .output_o(
        postnorm_addsub_output_o), .ine_o(postnorm_addsub_ine_o) );
  pre_norm_mul i_pre_norm_mul ( .clk_i(clk_i), .opa_i({s_opa_i[31], n1315, 
        n1311, n1310, n1314, n1309, n1316, n1312, n1303, n1286, n1298, n1305, 
        s_opa_i[19], n1306, s_opa_i[17], n1308, n1290, n1272, n1285, 
        s_opa_i[12], n1287, n1280, n1278, n1276, s_opa_i[7], n1282, n1284, 
        n1274, s_opa_i[3], n1275, n1294, n1302}), .opb_i({n1233, n1288, n1267, 
        n1268, n1277, n1263, n1266, n1269, s_opb_i[23], n1222, s_opb_i[21:19], 
        n1238, n1248, s_opb_i[16:15], n1262, n1227, n1226, n1225, n1240, 
        s_opb_i[9], n1228, n1230, s_opb_i[6:4], n1229, s_opb_i[2], n1260, 
        n1253}), .exp_10_o(pre_norm_mul_exp_10), .fracta_24_o(
        pre_norm_mul_fracta_24), .fractb_24_o(pre_norm_mul_fractb_24) );
  post_norm_mul i_post_norm_mul ( .clk_i(clk_i), .opa_i({s_opa_i[31], n1315, 
        n1311, n1310, n1314, n1309, n1316, n1312, n1303, n1286, n1298, n1305, 
        n1300, s_opa_i[18], n1301, s_opa_i[16], n1290, s_opa_i[14:13], n1292, 
        s_opa_i[11], n1280, n1278, s_opa_i[8], n1291, n1282, n1284, n1274, 
        n1270, n1275, n1293, s_opa_i[0]}), .opb_i({n1233, s_opb_i[30:29], 
        n1268, n1277, n1263, n1266, s_opb_i[24:22], n1236, n1224, 
        s_opb_i[19:17], n1245, n1255, s_opb_i[14], n1227, n1226, 
        s_opb_i[11:10], n1231, n1228, n1230, n1257, s_opb_i[5], n1242, n1229, 
        s_opb_i[2:1], n1250}), .exp_10_i(pre_norm_mul_exp_10), .fract_48_i(
        mul_fract_48), .sign_i(mul_24_sign), .rmode_i({n1217, n1221}), 
        .output_o(post_norm_mul_output), .ine_o(post_norm_mul_ine) );
  pre_norm_div i_pre_norm_div ( .clk_i(clk_i), .opa_i({s_opa_i[31], n1315, 
        n1311, n1310, n1314, n1309, n1316, n1312, n1303, n1286, n1298, 
        s_opa_i[20], n1300, n1306, s_opa_i[17], n1308, s_opa_i[15], n1272, 
        n1285, n1292, n1287, n1280, s_opa_i[9], n1276, n1291, n1282, n1284, 
        n1274, n1270, n1275, n1296, s_opa_i[0]}), .opb_i({n1233, n1288, n1267, 
        s_opb_i[28:25], n1269, s_opb_i[23], n1222, n1236, n1224, n1237, n1238, 
        n1248, n1245, n1255, n1262, s_opb_i[13:11], n1240, s_opb_i[9:7], n1257, 
        n1247, n1242, s_opb_i[3], n1243, n1260, n1252}), .exp_10_o(
        pre_norm_div_exp), .dvdnd_50_o({pre_norm_div_dvdnd[49:26], 
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26}), .dvsor_27_o({SYNOPSYS_UNCONNECTED_27, 
        SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, 
        pre_norm_div_dvsor[23:0]}) );
  post_norm_div i_post_norm_div ( .clk_i(clk_i), .opa_i({s_opa_i[31], n1315, 
        n1311, n1310, n1314, n1309, n1316, n1312, n1303, s_opa_i[22:20], n1300, 
        s_opa_i[18], n1301, s_opa_i[16], n1290, s_opa_i[14:12], n1287, n1280, 
        s_opa_i[9:8], n1291, s_opa_i[6], n1284, n1274, s_opa_i[3:2], n1296, 
        n1302}), .opb_i({n1233, n1288, n1267, n1268, s_opb_i[27], n1263, n1266, 
        n1269, n1258, s_opb_i[22:21], n1224, n1237, s_opb_i[18:11], n1240, 
        n1231, s_opb_i[8:7], n1257, n1247, n1242, s_opb_i[3], n1243, 
        s_opb_i[1], n1251}), .qutnt_i(serial_div_qutnt), .rmndr_i(
        serial_div_rmndr), .exp_10_i(pre_norm_div_exp), .sign_i(
        serial_div_sign), .rmode_i({n1216, n1221}), .output_o(
        post_norm_div_output), .ine_o(post_norm_div_ine) );
  pre_norm_sqrt i_pre_norm_sqrt ( .clk_i(clk_i), .opa_i({s_opa_i[31], n1315, 
        n1311, n1310, n1314, n1309, n1316, n1312, n1303, n1286, n1298, n1305, 
        n1300, n1306, n1301, n1308, n1290, n1272, n1285, n1292, s_opa_i[11], 
        n1280, n1278, n1276, n1291, n1282, n1284, s_opa_i[4], n1270, n1275, 
        n1295, n1302}), .fracta_52_o({pre_norm_sqrt_fracta_o[51:27], 
        SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, 
        SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33, 
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, 
        SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, 
        SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49, 
        SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51, 
        SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53, 
        SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55, 
        SYNOPSYS_UNCONNECTED_56}), .exp_o(pre_norm_sqrt_exp_o) );
  post_norm_sqrt i_post_norm_sqrt ( .clk_i(clk_i), .opa_i({s_opa_i[31], n1315, 
        n1311, n1310, n1314, n1309, n1316, n1312, n1303, n1286, n1298, n1305, 
        n1300, n1306, n1301, n1308, s_opa_i[15], n1272, s_opa_i[13], n1292, 
        n1287, s_opa_i[10:5], n1274, n1270, n1275, n1293, n1302}), 
        .fract_26_i(sqrt_sqr_o), .exp_i(pre_norm_sqrt_exp_o), .ine_i(
        sqrt_ine_o), .rmode_i({n1218, n1221}), .output_o(post_norm_sqrt_output), .ine_o(post_norm_sqrt_ine_o) );
  mul_24 i_mul_24 ( .clk_i(clk_i), .fracta_i(pre_norm_mul_fracta_24), 
        .fractb_i(pre_norm_mul_fractb_24), .signa_i(n1265), .signb_i(n1234), 
        .start_i(start_i), .fract_o(mul_fract_48), .sign_o(mul_24_sign) );
  serial_mul i_serial_mul ( .clk_i(clk_i), .fracta_i(pre_norm_mul_fracta_24), 
        .fractb_i(pre_norm_mul_fractb_24), .signa_i(n1265), .signb_i(n1233), 
        .start_i(n1191), .fract_o({SYNOPSYS_UNCONNECTED_57, 
        SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59, 
        SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61, 
        SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63, 
        SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65, 
        SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67, 
        SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69, 
        SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71, 
        SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73, 
        SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75, 
        SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77, 
        SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79, 
        SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81, 
        SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83, 
        SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85, 
        SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87, 
        SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89, 
        SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91, 
        SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93, 
        SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95, 
        SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97, 
        SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101, 
        SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103, 
        SYNOPSYS_UNCONNECTED_104}) );
  serial_div i_serial_div ( .clk_i(clk_i), .dvdnd_i({pre_norm_div_dvdnd[49:26], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .dvsor_i({1'b0, 1'b0, 1'b0, pre_norm_div_dvsor[23:0]}), 
        .sign_dvd_i(n1265), .sign_div_i(n1233), .start_i(n1191), .qutnt_o(
        serial_div_qutnt), .rmndr_o(serial_div_rmndr), .sign_o(serial_div_sign), .div_zero_o(serial_div_div_zero) );
  sqrt_RD_WIDTH52_SQ_WIDTH26 i_sqrt ( .clk_i(clk_i), .rad_i({
        pre_norm_sqrt_fracta_o[51:27], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .start_i(n1191), .sqr_o(sqrt_sqr_o), .ine_o(sqrt_ine_o) );
  dff s_count_reg_0_ ( .Q(s_count_0_), .D(n903), .CLK(clk_i) );
  dff s_count_reg_1_ ( .Q(s_count_1_), .D(n904), .CLK(clk_i) );
  dff s_count_reg_2_ ( .Q(s_count_2_), .D(n905), .CLK(clk_i) );
  dff s_count_reg_3_ ( .Q(s_count_3_), .D(n906), .CLK(clk_i) );
  dff s_count_reg_4_ ( .Q(s_count_4_), .D(n907), .CLK(clk_i) );
  dff s_count_reg_5_ ( .Q(s_count_5_), .D(n908), .CLK(clk_i) );
  dff s_count_reg_6_ ( .Q(s_count_6_), .D(n909), .CLK(clk_i) );
  dff s_count_reg_7_ ( .Q(s_count_7_), .D(n910), .CLK(clk_i) );
  dff s_count_reg_8_ ( .Q(s_count_8_), .D(n911), .CLK(clk_i) );
  dff s_count_reg_9_ ( .Q(s_count_9_), .D(n912), .CLK(clk_i) );
  dff s_count_reg_10_ ( .Q(s_count_10_), .D(n913), .CLK(clk_i) );
  dff s_count_reg_11_ ( .Q(s_count_11_), .D(n914), .CLK(clk_i) );
  dff s_count_reg_12_ ( .Q(s_count_12_), .D(n915), .CLK(clk_i) );
  dff s_count_reg_13_ ( .Q(s_count_13_), .D(n916), .CLK(clk_i) );
  dff s_count_reg_14_ ( .Q(s_count_14_), .D(n917), .CLK(clk_i) );
  dff s_count_reg_15_ ( .Q(s_count_15_), .D(n918), .CLK(clk_i) );
  dff s_count_reg_16_ ( .Q(s_count_16_), .D(n919), .CLK(clk_i) );
  dff s_count_reg_17_ ( .Q(s_count_17_), .D(n920), .CLK(clk_i) );
  dff s_count_reg_18_ ( .Q(s_count_18_), .D(n921), .CLK(clk_i) );
  dff s_count_reg_19_ ( .Q(s_count_19_), .D(n922), .CLK(clk_i) );
  dff s_count_reg_20_ ( .Q(s_count_20_), .D(n923), .CLK(clk_i) );
  dff s_count_reg_21_ ( .Q(s_count_21_), .D(n924), .CLK(clk_i) );
  dff s_count_reg_22_ ( .Q(s_count_22_), .D(n925), .CLK(clk_i) );
  dff s_count_reg_23_ ( .Q(s_count_23_), .D(n926), .CLK(clk_i) );
  dff s_count_reg_24_ ( .Q(s_count_24_), .D(n927), .CLK(clk_i) );
  dff s_count_reg_25_ ( .Q(s_count_25_), .D(n928), .CLK(clk_i) );
  dff s_count_reg_26_ ( .Q(s_count_26_), .D(n929), .CLK(clk_i) );
  dff s_count_reg_27_ ( .Q(s_count_27_), .D(n930), .CLK(clk_i) );
  dff s_count_reg_28_ ( .Q(s_count_28_), .D(n931), .CLK(clk_i) );
  dff s_count_reg_29_ ( .Q(s_count_29_), .D(n932), .CLK(clk_i) );
  dff s_count_reg_30_ ( .Q(s_count_30_), .D(n933), .CLK(clk_i) );
  dff s_count_reg_31_ ( .Q(s_count_31_), .D(n934), .CLK(clk_i) );
  dff s_state_reg ( .Q(s_state), .D(n935), .CLK(clk_i) );
  dff ready_o_reg ( .Q(ready_o), .QB(n902), .D(n1104), .CLK(clk_i) );
  dff s_opa_i_reg_31_ ( .Q(s_opa_i[31]), .QB(n1264), .D(opa_i[31]), .CLK(clk_i) );
  dff s_opa_i_reg_30_ ( .Q(s_opa_i[30]), .QB(n952), .D(opa_i[30]), .CLK(clk_i)
         );
  dff s_opa_i_reg_29_ ( .Q(s_opa_i[29]), .QB(n951), .D(opa_i[29]), .CLK(clk_i)
         );
  dff s_opa_i_reg_28_ ( .Q(s_opa_i[28]), .QB(n950), .D(opa_i[28]), .CLK(clk_i)
         );
  dff s_opa_i_reg_27_ ( .Q(s_opa_i[27]), .QB(n949), .D(opa_i[27]), .CLK(clk_i)
         );
  dff s_opa_i_reg_26_ ( .Q(s_opa_i[26]), .QB(n948), .D(opa_i[26]), .CLK(clk_i)
         );
  dff s_opa_i_reg_25_ ( .Q(s_opa_i[25]), .QB(n947), .D(opa_i[25]), .CLK(clk_i)
         );
  dff s_opa_i_reg_24_ ( .Q(s_opa_i[24]), .QB(n946), .D(opa_i[24]), .CLK(clk_i)
         );
  dff s_opa_i_reg_23_ ( .Q(s_opa_i[23]), .QB(n945), .D(opa_i[23]), .CLK(clk_i)
         );
  dff s_opa_i_reg_22_ ( .Q(s_opa_i[22]), .QB(n682), .D(opa_i[22]), .CLK(clk_i)
         );
  dff s_opa_i_reg_21_ ( .Q(s_opa_i[21]), .D(opa_i[21]), .CLK(clk_i) );
  dff s_opa_i_reg_20_ ( .Q(s_opa_i[20]), .QB(n1304), .D(opa_i[20]), .CLK(clk_i) );
  dff s_opa_i_reg_19_ ( .Q(s_opa_i[19]), .QB(n1417), .D(opa_i[19]), .CLK(clk_i) );
  dff s_opa_i_reg_18_ ( .Q(s_opa_i[18]), .QB(n1416), .D(opa_i[18]), .CLK(clk_i) );
  dff s_opa_i_reg_17_ ( .Q(s_opa_i[17]), .QB(n1418), .D(opa_i[17]), .CLK(clk_i) );
  dff s_opa_i_reg_16_ ( .Q(s_opa_i[16]), .QB(n1307), .D(opa_i[16]), .CLK(clk_i) );
  dff s_opa_i_reg_15_ ( .Q(s_opa_i[15]), .QB(n1289), .D(opa_i[15]), .CLK(clk_i) );
  dff s_opa_i_reg_14_ ( .Q(s_opa_i[14]), .QB(n1271), .D(opa_i[14]), .CLK(clk_i) );
  dff s_opa_i_reg_13_ ( .Q(s_opa_i[13]), .QB(n678), .D(opa_i[13]), .CLK(clk_i)
         );
  dff s_opa_i_reg_12_ ( .Q(s_opa_i[12]), .QB(n677), .D(opa_i[12]), .CLK(clk_i)
         );
  dff s_opa_i_reg_11_ ( .Q(s_opa_i[11]), .QB(n676), .D(opa_i[11]), .CLK(clk_i)
         );
  dff s_opa_i_reg_10_ ( .Q(s_opa_i[10]), .QB(n1279), .D(opa_i[10]), .CLK(clk_i) );
  dff s_opa_i_reg_9_ ( .Q(s_opa_i[9]), .QB(n675), .D(opa_i[9]), .CLK(clk_i) );
  dff s_opa_i_reg_8_ ( .Q(s_opa_i[8]), .QB(n674), .D(opa_i[8]), .CLK(clk_i) );
  dff s_opa_i_reg_7_ ( .Q(s_opa_i[7]), .QB(n673), .D(opa_i[7]), .CLK(clk_i) );
  dff s_opa_i_reg_6_ ( .Q(s_opa_i[6]), .QB(n1281), .D(opa_i[6]), .CLK(clk_i)
         );
  dff s_opa_i_reg_5_ ( .Q(s_opa_i[5]), .QB(n1283), .D(opa_i[5]), .CLK(clk_i)
         );
  dff s_opa_i_reg_4_ ( .Q(s_opa_i[4]), .QB(n1273), .D(opa_i[4]), .CLK(clk_i)
         );
  dff s_opa_i_reg_3_ ( .Q(s_opa_i[3]), .QB(n672), .D(opa_i[3]), .CLK(clk_i) );
  dff s_opa_i_reg_2_ ( .Q(s_opa_i[2]), .QB(n671), .D(opa_i[2]), .CLK(clk_i) );
  dff s_opa_i_reg_1_ ( .Q(s_opa_i[1]), .D(opa_i[1]), .CLK(clk_i) );
  dff s_opa_i_reg_0_ ( .Q(s_opa_i[0]), .QB(n670), .D(opa_i[0]), .CLK(clk_i) );
  dff s_opb_i_reg_31_ ( .Q(s_opb_i[31]), .D(opb_i[31]), .CLK(clk_i) );
  dff s_opb_i_reg_30_ ( .Q(s_opb_i[30]), .QB(n944), .D(opb_i[30]), .CLK(clk_i)
         );
  dff s_opb_i_reg_29_ ( .Q(s_opb_i[29]), .QB(n943), .D(opb_i[29]), .CLK(clk_i)
         );
  dff s_opb_i_reg_28_ ( .Q(s_opb_i[28]), .QB(n942), .D(opb_i[28]), .CLK(clk_i)
         );
  dff s_opb_i_reg_27_ ( .Q(s_opb_i[27]), .QB(n941), .D(opb_i[27]), .CLK(clk_i)
         );
  dff s_opb_i_reg_26_ ( .Q(s_opb_i[26]), .QB(n940), .D(opb_i[26]), .CLK(clk_i)
         );
  dff s_opb_i_reg_25_ ( .Q(s_opb_i[25]), .QB(n939), .D(opb_i[25]), .CLK(clk_i)
         );
  dff s_opb_i_reg_24_ ( .Q(s_opb_i[24]), .QB(n938), .D(opb_i[24]), .CLK(clk_i)
         );
  dff s_opb_i_reg_23_ ( .Q(s_opb_i[23]), .QB(n937), .D(opb_i[23]), .CLK(clk_i)
         );
  dff s_opb_i_reg_22_ ( .Q(s_opb_i[22]), .QB(n669), .D(opb_i[22]), .CLK(clk_i)
         );
  dff s_opb_i_reg_21_ ( .Q(s_opb_i[21]), .QB(n1235), .D(opb_i[21]), .CLK(clk_i) );
  dff s_opb_i_reg_20_ ( .Q(s_opb_i[20]), .QB(n1223), .D(opb_i[20]), .CLK(clk_i) );
  dff s_opb_i_reg_19_ ( .Q(s_opb_i[19]), .QB(n1414), .D(opb_i[19]), .CLK(clk_i) );
  dff s_opb_i_reg_18_ ( .Q(s_opb_i[18]), .QB(n1413), .D(opb_i[18]), .CLK(clk_i) );
  dff s_opb_i_reg_17_ ( .Q(s_opb_i[17]), .QB(n1415), .D(opb_i[17]), .CLK(clk_i) );
  dff s_opb_i_reg_16_ ( .Q(s_opb_i[16]), .QB(n1244), .D(opb_i[16]), .CLK(clk_i) );
  dff s_opb_i_reg_15_ ( .Q(s_opb_i[15]), .QB(n1254), .D(opb_i[15]), .CLK(clk_i) );
  dff s_opb_i_reg_14_ ( .Q(s_opb_i[14]), .QB(n1261), .D(opb_i[14]), .CLK(clk_i) );
  dff s_opb_i_reg_13_ ( .Q(s_opb_i[13]), .QB(n665), .D(opb_i[13]), .CLK(clk_i)
         );
  dff s_opb_i_reg_12_ ( .Q(s_opb_i[12]), .QB(n664), .D(opb_i[12]), .CLK(clk_i)
         );
  dff s_opb_i_reg_11_ ( .Q(s_opb_i[11]), .QB(n663), .D(opb_i[11]), .CLK(clk_i)
         );
  dff s_opb_i_reg_10_ ( .Q(s_opb_i[10]), .QB(n1239), .D(opb_i[10]), .CLK(clk_i) );
  dff s_opb_i_reg_9_ ( .Q(s_opb_i[9]), .QB(n662), .D(opb_i[9]), .CLK(clk_i) );
  dff s_opb_i_reg_8_ ( .Q(s_opb_i[8]), .QB(n661), .D(opb_i[8]), .CLK(clk_i) );
  dff s_opb_i_reg_7_ ( .Q(s_opb_i[7]), .QB(n660), .D(opb_i[7]), .CLK(clk_i) );
  dff s_opb_i_reg_6_ ( .Q(s_opb_i[6]), .QB(n1256), .D(opb_i[6]), .CLK(clk_i)
         );
  dff s_opb_i_reg_5_ ( .Q(s_opb_i[5]), .QB(n1246), .D(opb_i[5]), .CLK(clk_i)
         );
  dff s_opb_i_reg_4_ ( .Q(s_opb_i[4]), .QB(n1241), .D(opb_i[4]), .CLK(clk_i)
         );
  dff s_opb_i_reg_3_ ( .Q(s_opb_i[3]), .QB(n659), .D(opb_i[3]), .CLK(clk_i) );
  dff s_opb_i_reg_2_ ( .Q(s_opb_i[2]), .QB(n658), .D(opb_i[2]), .CLK(clk_i) );
  dff s_opb_i_reg_1_ ( .Q(s_opb_i[1]), .QB(n1259), .D(opb_i[1]), .CLK(clk_i)
         );
  dff s_opb_i_reg_0_ ( .Q(s_opb_i[0]), .QB(n657), .D(opb_i[0]), .CLK(clk_i) );
  dff s_fpu_op_i_reg_2_ ( .Q(n1411), .D(fpu_op_i[2]), .CLK(clk_i) );
  dff s_fpu_op_i_reg_1_ ( .Q(n1412), .D(fpu_op_i[1]), .CLK(clk_i) );
  dff s_fpu_op_i_reg_0_ ( .Q(s_fpu_op_i_0_), .QB(n654), .D(fpu_op_i[0]), .CLK(
        clk_i) );
  dff s_rmode_i_reg_1_ ( .Q(s_rmode_i[1]), .D(rmode_i[1]), .CLK(clk_i) );
  dff s_rmode_i_reg_0_ ( .Q(s_rmode_i[0]), .QB(n1220), .D(rmode_i[0]), .CLK(
        clk_i) );
  dff output_o_reg_31_ ( .Q(output_o[31]), .D(s_output_o_31_), .CLK(clk_i) );
  dff output_o_reg_30_ ( .Q(output_o[30]), .D(s_output_o_30_), .CLK(clk_i) );
  dff output_o_reg_29_ ( .Q(output_o[29]), .D(s_output_o_29_), .CLK(clk_i) );
  dff output_o_reg_28_ ( .Q(output_o[28]), .D(s_output_o_28_), .CLK(clk_i) );
  dff output_o_reg_27_ ( .Q(output_o[27]), .D(s_output_o_27_), .CLK(clk_i) );
  dff output_o_reg_26_ ( .Q(output_o[26]), .D(s_output_o_26_), .CLK(clk_i) );
  dff output_o_reg_25_ ( .Q(output_o[25]), .D(s_output_o_25_), .CLK(clk_i) );
  dff output_o_reg_24_ ( .Q(output_o[24]), .D(s_output_o_24_), .CLK(clk_i) );
  dff output_o_reg_23_ ( .Q(output_o[23]), .D(n959), .CLK(clk_i) );
  dff output_o_reg_22_ ( .Q(output_o[22]), .D(s_output_o_22_), .CLK(clk_i) );
  dff output_o_reg_21_ ( .Q(output_o[21]), .D(s_output_o_21_), .CLK(clk_i) );
  dff output_o_reg_20_ ( .Q(output_o[20]), .D(s_output_o_20_), .CLK(clk_i) );
  dff output_o_reg_19_ ( .Q(output_o[19]), .D(s_output_o_19_), .CLK(clk_i) );
  dff output_o_reg_18_ ( .Q(output_o[18]), .D(s_output_o_18_), .CLK(clk_i) );
  dff output_o_reg_17_ ( .Q(output_o[17]), .D(s_output_o_17_), .CLK(clk_i) );
  dff output_o_reg_16_ ( .Q(output_o[16]), .D(s_output_o_16_), .CLK(clk_i) );
  dff output_o_reg_15_ ( .Q(output_o[15]), .D(s_output_o_15_), .CLK(clk_i) );
  dff output_o_reg_14_ ( .Q(output_o[14]), .D(s_output_o_14_), .CLK(clk_i) );
  dff output_o_reg_13_ ( .Q(output_o[13]), .D(s_output_o_13_), .CLK(clk_i) );
  dff output_o_reg_12_ ( .Q(output_o[12]), .D(s_output_o_12_), .CLK(clk_i) );
  dff output_o_reg_11_ ( .Q(output_o[11]), .D(s_output_o_11_), .CLK(clk_i) );
  dff output_o_reg_10_ ( .Q(output_o[10]), .D(s_output_o_10_), .CLK(clk_i) );
  dff output_o_reg_9_ ( .Q(output_o[9]), .D(s_output_o_9_), .CLK(clk_i) );
  dff output_o_reg_8_ ( .Q(output_o[8]), .D(s_output_o_8_), .CLK(clk_i) );
  dff output_o_reg_7_ ( .Q(output_o[7]), .D(s_output_o_7_), .CLK(clk_i) );
  dff output_o_reg_6_ ( .Q(output_o[6]), .D(s_output_o_6_), .CLK(clk_i) );
  dff output_o_reg_5_ ( .Q(output_o[5]), .D(s_output_o_5_), .CLK(clk_i) );
  dff output_o_reg_4_ ( .Q(output_o[4]), .D(s_output_o_4_), .CLK(clk_i) );
  dff output_o_reg_3_ ( .Q(output_o[3]), .D(s_output_o_3_), .CLK(clk_i) );
  dff output_o_reg_2_ ( .Q(output_o[2]), .D(s_output_o_2_), .CLK(clk_i) );
  dff output_o_reg_1_ ( .Q(output_o[1]), .D(s_output_o_1_), .CLK(clk_i) );
  dff output_o_reg_0_ ( .Q(output_o[0]), .D(s_output_o_0_), .CLK(clk_i) );
  dff s_output1_reg_31_ ( .Q(s_output1_31_), .D(s_output1408_31_), .CLK(clk_i)
         );
  dff s_output1_reg_30_ ( .Q(s_output_o_30_), .D(s_output1408_30_), .CLK(clk_i) );
  dff s_output1_reg_29_ ( .Q(s_output_o_29_), .D(s_output1408_29_), .CLK(clk_i) );
  dff s_output1_reg_28_ ( .Q(s_output_o_28_), .D(s_output1408_28_), .CLK(clk_i) );
  dff s_output1_reg_27_ ( .Q(s_output_o_27_), .D(s_output1408_27_), .CLK(clk_i) );
  dff s_output1_reg_26_ ( .Q(s_output_o_26_), .D(s_output1408_26_), .CLK(clk_i) );
  dff s_output1_reg_25_ ( .Q(s_output_o_25_), .D(s_output1408_25_), .CLK(clk_i) );
  dff s_output1_reg_24_ ( .Q(s_output_o_24_), .D(s_output1408_24_), .CLK(clk_i) );
  dff s_output1_reg_23_ ( .Q(s_output1_23_), .D(s_output1408_23_), .CLK(clk_i)
         );
  dff s_output1_reg_22_ ( .Q(s_output1_22_), .D(s_output1408_22_), .CLK(clk_i)
         );
  dff s_output1_reg_21_ ( .Q(s_output1_21_), .D(s_output1408_21_), .CLK(clk_i)
         );
  dff s_output1_reg_20_ ( .Q(s_output1_20_), .D(s_output1408_20_), .CLK(clk_i)
         );
  dff s_output1_reg_19_ ( .Q(s_output1_19_), .D(s_output1408_19_), .CLK(clk_i)
         );
  dff s_output1_reg_18_ ( .Q(s_output1_18_), .D(s_output1408_18_), .CLK(clk_i)
         );
  dff s_output1_reg_17_ ( .Q(s_output1_17_), .D(s_output1408_17_), .CLK(clk_i)
         );
  dff s_output1_reg_16_ ( .Q(s_output1_16_), .D(s_output1408_16_), .CLK(clk_i)
         );
  dff s_output1_reg_15_ ( .Q(n653), .D(s_output1408_15_), .CLK(clk_i) );
  dff s_output1_reg_14_ ( .Q(n652), .D(s_output1408_14_), .CLK(clk_i) );
  dff s_output1_reg_13_ ( .Q(n651), .D(s_output1408_13_), .CLK(clk_i) );
  dff s_output1_reg_12_ ( .Q(n650), .D(s_output1408_12_), .CLK(clk_i) );
  dff s_output1_reg_11_ ( .Q(s_output1_11_), .D(s_output1408_11_), .CLK(clk_i)
         );
  dff s_output1_reg_10_ ( .Q(s_output1_10_), .D(s_output1408_10_), .CLK(clk_i)
         );
  dff s_output1_reg_9_ ( .Q(s_output1_9_), .D(s_output1408_9_), .CLK(clk_i) );
  dff s_output1_reg_8_ ( .Q(s_output1_8_), .D(s_output1408_8_), .CLK(clk_i) );
  dff s_output1_reg_7_ ( .Q(s_output1_7_), .D(s_output1408_7_), .CLK(clk_i) );
  dff s_output1_reg_6_ ( .Q(s_output1_6_), .D(s_output1408_6_), .CLK(clk_i) );
  dff s_output1_reg_5_ ( .Q(s_output1_5_), .D(s_output1408_5_), .CLK(clk_i) );
  dff s_output1_reg_4_ ( .Q(s_output1_4_), .D(s_output1408_4_), .CLK(clk_i) );
  dff s_output1_reg_3_ ( .Q(s_output1_3_), .D(s_output1408_3_), .CLK(clk_i) );
  dff s_output1_reg_2_ ( .Q(s_output1_2_), .D(s_output1408_2_), .CLK(clk_i) );
  dff s_output1_reg_1_ ( .Q(s_output1_1_), .D(s_output1408_1_), .CLK(clk_i) );
  dff s_output1_reg_0_ ( .Q(s_output1_0_), .D(s_output1408_0_), .CLK(clk_i) );
  dff s_start_i_reg ( .Q(s_state213), .QB(n1190), .D(start_i), .CLK(clk_i) );
  dff ine_o_reg ( .Q(ine_o), .D(s_ine_o), .CLK(clk_i) );
  dff overflow_o_reg ( .Q(overflow_o), .D(n961), .CLK(clk_i) );
  dff underflow_o_reg ( .Q(underflow_o), .D(n965), .CLK(clk_i) );
  dff div_zero_o_reg ( .Q(div_zero_o), .D(s_div_zero_o), .CLK(clk_i) );
  dff inf_o_reg ( .Q(inf_o), .D(s_inf_o), .CLK(clk_i) );
  dff zero_o_reg ( .Q(zero_o), .D(s_zero_o), .CLK(clk_i) );
  dff qnan_o_reg ( .Q(qnan_o), .D(s_qnan_o), .CLK(clk_i) );
  dff snan_o_reg ( .Q(snan_o), .D(s_snan_o), .CLK(clk_i) );
  dff s_ine_o_reg ( .Q(s_ine_o), .D(s_ine_o415), .CLK(clk_i) );
  buf04 U478 ( .Y(n1275), .A(s_opa_i[2]) );
  xor2 U479 ( .Y(n953), .A0(n1233), .A1(n654) );
  inv01 U480 ( .Y(n954), .A(n953) );
  inv01 U481 ( .Y(n1405), .A(n955) );
  nor02 U482 ( .Y(n956), .A0(n1317), .A1(n1325) );
  inv01 U483 ( .Y(n957), .A(n1195) );
  nor02 U484 ( .Y(n955), .A0(n956), .A1(n957) );
  or02 U485 ( .Y(n958), .A0(n1347), .A1(n1348) );
  inv01 U486 ( .Y(n959), .A(n958) );
  or02 U487 ( .Y(n960), .A0(n1329), .A1(n1189) );
  inv01 U488 ( .Y(n961), .A(n960) );
  ao21 U489 ( .Y(n962), .A0(s_rmode_i[0]), .A1(n1352), .B0(n966) );
  inv01 U490 ( .Y(n963), .A(n962) );
  or02 U491 ( .Y(n964), .A0(n1328), .A1(n1329) );
  inv01 U492 ( .Y(n965), .A(n964) );
  buf02 U493 ( .Y(n966), .A(n1372) );
  ao22 U494 ( .Y(n967), .A0(post_norm_div_output[23]), .A1(n1325), .B0(
        post_norm_sqrt_output[23]), .B1(n1317) );
  inv01 U495 ( .Y(n968), .A(n967) );
  ao22 U496 ( .Y(n969), .A0(post_norm_div_output[22]), .A1(n1325), .B0(
        post_norm_sqrt_output[22]), .B1(n1317) );
  inv01 U497 ( .Y(n970), .A(n969) );
  ao22 U498 ( .Y(n971), .A0(post_norm_div_output[24]), .A1(n1325), .B0(
        post_norm_sqrt_output[24]), .B1(n1317) );
  inv01 U499 ( .Y(n972), .A(n971) );
  ao22 U500 ( .Y(n973), .A0(post_norm_div_output[21]), .A1(n1325), .B0(
        post_norm_sqrt_output[21]), .B1(n1317) );
  inv01 U501 ( .Y(n974), .A(n973) );
  ao22 U502 ( .Y(n975), .A0(post_norm_div_output[25]), .A1(n1325), .B0(
        post_norm_sqrt_output[25]), .B1(n1317) );
  inv01 U503 ( .Y(n976), .A(n975) );
  ao22 U504 ( .Y(n977), .A0(post_norm_div_output[20]), .A1(n1325), .B0(
        post_norm_sqrt_output[20]), .B1(n1317) );
  inv01 U505 ( .Y(n978), .A(n977) );
  ao22 U506 ( .Y(n979), .A0(post_norm_div_output[26]), .A1(n1325), .B0(
        post_norm_sqrt_output[26]), .B1(n1317) );
  inv01 U507 ( .Y(n980), .A(n979) );
  ao22 U508 ( .Y(n981), .A0(post_norm_div_output[1]), .A1(n1325), .B0(
        post_norm_sqrt_output[1]), .B1(n1317) );
  inv01 U509 ( .Y(n982), .A(n981) );
  ao22 U510 ( .Y(n983), .A0(post_norm_div_output[27]), .A1(n1325), .B0(
        post_norm_sqrt_output[27]), .B1(n1317) );
  inv01 U511 ( .Y(n984), .A(n983) );
  ao22 U512 ( .Y(n985), .A0(post_norm_div_output[19]), .A1(n1325), .B0(
        post_norm_sqrt_output[19]), .B1(n1317) );
  inv01 U513 ( .Y(n986), .A(n985) );
  ao22 U514 ( .Y(n987), .A0(post_norm_div_output[28]), .A1(n1325), .B0(
        post_norm_sqrt_output[28]), .B1(n1317) );
  inv01 U515 ( .Y(n988), .A(n987) );
  ao22 U516 ( .Y(n989), .A0(post_norm_div_output[18]), .A1(n1325), .B0(
        post_norm_sqrt_output[18]), .B1(n1317) );
  inv01 U517 ( .Y(n990), .A(n989) );
  ao22 U518 ( .Y(n991), .A0(post_norm_div_output[29]), .A1(n1325), .B0(
        post_norm_sqrt_output[29]), .B1(n1317) );
  inv01 U519 ( .Y(n992), .A(n991) );
  ao22 U520 ( .Y(n993), .A0(post_norm_div_output[17]), .A1(n1325), .B0(
        post_norm_sqrt_output[17]), .B1(n1317) );
  inv01 U521 ( .Y(n994), .A(n993) );
  ao22 U522 ( .Y(n995), .A0(post_norm_div_output[2]), .A1(n1325), .B0(
        post_norm_sqrt_output[2]), .B1(n1317) );
  inv01 U523 ( .Y(n996), .A(n995) );
  ao22 U524 ( .Y(n997), .A0(post_norm_div_output[16]), .A1(n1325), .B0(
        post_norm_sqrt_output[16]), .B1(n1317) );
  inv01 U525 ( .Y(n998), .A(n997) );
  ao22 U526 ( .Y(n999), .A0(post_norm_div_output[30]), .A1(n1325), .B0(
        post_norm_sqrt_output[30]), .B1(n1317) );
  inv01 U527 ( .Y(n1000), .A(n999) );
  ao22 U528 ( .Y(n1001), .A0(post_norm_div_output[15]), .A1(n1325), .B0(
        post_norm_sqrt_output[15]), .B1(n1317) );
  inv01 U529 ( .Y(n1002), .A(n1001) );
  ao22 U530 ( .Y(n1003), .A0(post_norm_div_output[31]), .A1(n1325), .B0(
        post_norm_sqrt_output[31]), .B1(n1317) );
  inv01 U531 ( .Y(n1004), .A(n1003) );
  ao22 U532 ( .Y(n1005), .A0(post_norm_div_output[14]), .A1(n1325), .B0(
        post_norm_sqrt_output[14]), .B1(n1317) );
  inv01 U533 ( .Y(n1006), .A(n1005) );
  ao22 U534 ( .Y(n1007), .A0(post_norm_div_output[3]), .A1(n1325), .B0(
        post_norm_sqrt_output[3]), .B1(n1317) );
  inv01 U535 ( .Y(n1008), .A(n1007) );
  ao22 U536 ( .Y(n1009), .A0(post_norm_div_output[13]), .A1(n1325), .B0(
        post_norm_sqrt_output[13]), .B1(n1317) );
  inv01 U537 ( .Y(n1010), .A(n1009) );
  ao22 U538 ( .Y(n1011), .A0(post_norm_div_output[4]), .A1(n1325), .B0(
        post_norm_sqrt_output[4]), .B1(n1317) );
  inv01 U539 ( .Y(n1012), .A(n1011) );
  ao22 U540 ( .Y(n1013), .A0(post_norm_div_output[12]), .A1(n1325), .B0(
        post_norm_sqrt_output[12]), .B1(n1317) );
  inv01 U541 ( .Y(n1014), .A(n1013) );
  ao22 U542 ( .Y(n1015), .A0(post_norm_div_output[5]), .A1(n1325), .B0(
        post_norm_sqrt_output[5]), .B1(n1317) );
  inv01 U543 ( .Y(n1016), .A(n1015) );
  ao22 U544 ( .Y(n1017), .A0(post_norm_div_output[11]), .A1(n1325), .B0(
        post_norm_sqrt_output[11]), .B1(n1317) );
  inv01 U545 ( .Y(n1018), .A(n1017) );
  ao22 U546 ( .Y(n1019), .A0(post_norm_div_output[6]), .A1(n1325), .B0(
        post_norm_sqrt_output[6]), .B1(n1317) );
  inv01 U547 ( .Y(n1020), .A(n1019) );
  ao22 U548 ( .Y(n1021), .A0(post_norm_div_output[10]), .A1(n1325), .B0(
        post_norm_sqrt_output[10]), .B1(n1317) );
  inv01 U549 ( .Y(n1022), .A(n1021) );
  ao22 U550 ( .Y(n1023), .A0(post_norm_div_output[7]), .A1(n1325), .B0(
        post_norm_sqrt_output[7]), .B1(n1317) );
  inv01 U551 ( .Y(n1024), .A(n1023) );
  ao22 U552 ( .Y(n1025), .A0(post_norm_div_output[0]), .A1(n1325), .B0(
        post_norm_sqrt_output[0]), .B1(n1317) );
  inv01 U553 ( .Y(n1026), .A(n1025) );
  ao22 U554 ( .Y(n1027), .A0(post_norm_div_output[8]), .A1(n1325), .B0(
        post_norm_sqrt_output[8]), .B1(n1317) );
  inv01 U555 ( .Y(n1028), .A(n1027) );
  ao22 U556 ( .Y(n1029), .A0(post_norm_div_ine), .A1(n1325), .B0(
        post_norm_sqrt_ine_o), .B1(n1317) );
  inv01 U557 ( .Y(n1030), .A(n1029) );
  ao22 U558 ( .Y(n1031), .A0(post_norm_div_output[9]), .A1(n1325), .B0(
        post_norm_sqrt_output[9]), .B1(n1317) );
  inv01 U559 ( .Y(n1032), .A(n1031) );
  ao22 U560 ( .Y(n1033), .A0(postnorm_addsub_output_o[23]), .A1(n1326), .B0(
        post_norm_mul_output[23]), .B1(n1318) );
  inv01 U561 ( .Y(n1034), .A(n1033) );
  ao22 U562 ( .Y(n1035), .A0(postnorm_addsub_output_o[24]), .A1(n1326), .B0(
        post_norm_mul_output[24]), .B1(n1318) );
  inv01 U563 ( .Y(n1036), .A(n1035) );
  ao22 U564 ( .Y(n1037), .A0(postnorm_addsub_output_o[22]), .A1(n1326), .B0(
        post_norm_mul_output[22]), .B1(n1318) );
  inv01 U565 ( .Y(n1038), .A(n1037) );
  ao22 U566 ( .Y(n1039), .A0(postnorm_addsub_output_o[25]), .A1(n1326), .B0(
        post_norm_mul_output[25]), .B1(n1318) );
  inv01 U567 ( .Y(n1040), .A(n1039) );
  ao22 U568 ( .Y(n1041), .A0(postnorm_addsub_output_o[21]), .A1(n1326), .B0(
        post_norm_mul_output[21]), .B1(n1318) );
  inv01 U569 ( .Y(n1042), .A(n1041) );
  ao22 U570 ( .Y(n1043), .A0(postnorm_addsub_output_o[26]), .A1(n1326), .B0(
        post_norm_mul_output[26]), .B1(n1318) );
  inv01 U571 ( .Y(n1044), .A(n1043) );
  ao22 U572 ( .Y(n1045), .A0(postnorm_addsub_output_o[20]), .A1(n1326), .B0(
        post_norm_mul_output[20]), .B1(n1318) );
  inv01 U573 ( .Y(n1046), .A(n1045) );
  ao22 U574 ( .Y(n1047), .A0(postnorm_addsub_output_o[27]), .A1(n1326), .B0(
        post_norm_mul_output[27]), .B1(n1318) );
  inv01 U575 ( .Y(n1048), .A(n1047) );
  ao22 U576 ( .Y(n1049), .A0(postnorm_addsub_output_o[1]), .A1(n1326), .B0(
        post_norm_mul_output[1]), .B1(n1318) );
  inv01 U577 ( .Y(n1050), .A(n1049) );
  ao22 U578 ( .Y(n1051), .A0(postnorm_addsub_output_o[28]), .A1(n1326), .B0(
        post_norm_mul_output[28]), .B1(n1318) );
  inv01 U579 ( .Y(n1052), .A(n1051) );
  ao22 U580 ( .Y(n1053), .A0(postnorm_addsub_output_o[19]), .A1(n1326), .B0(
        post_norm_mul_output[19]), .B1(n1318) );
  inv01 U581 ( .Y(n1054), .A(n1053) );
  ao22 U582 ( .Y(n1055), .A0(postnorm_addsub_output_o[29]), .A1(n1326), .B0(
        post_norm_mul_output[29]), .B1(n1318) );
  inv01 U583 ( .Y(n1056), .A(n1055) );
  ao22 U584 ( .Y(n1057), .A0(postnorm_addsub_output_o[18]), .A1(n1326), .B0(
        post_norm_mul_output[18]), .B1(n1318) );
  inv01 U585 ( .Y(n1058), .A(n1057) );
  ao22 U586 ( .Y(n1059), .A0(postnorm_addsub_output_o[2]), .A1(n1326), .B0(
        post_norm_mul_output[2]), .B1(n1318) );
  inv01 U587 ( .Y(n1060), .A(n1059) );
  ao22 U588 ( .Y(n1061), .A0(postnorm_addsub_output_o[17]), .A1(n1326), .B0(
        post_norm_mul_output[17]), .B1(n1318) );
  inv01 U589 ( .Y(n1062), .A(n1061) );
  ao22 U590 ( .Y(n1063), .A0(postnorm_addsub_output_o[30]), .A1(n1326), .B0(
        post_norm_mul_output[30]), .B1(n1318) );
  inv01 U591 ( .Y(n1064), .A(n1063) );
  ao22 U592 ( .Y(n1065), .A0(postnorm_addsub_output_o[16]), .A1(n1326), .B0(
        post_norm_mul_output[16]), .B1(n1318) );
  inv01 U593 ( .Y(n1066), .A(n1065) );
  ao22 U594 ( .Y(n1067), .A0(postnorm_addsub_output_o[31]), .A1(n1326), .B0(
        post_norm_mul_output[31]), .B1(n1318) );
  inv01 U595 ( .Y(n1068), .A(n1067) );
  ao22 U596 ( .Y(n1069), .A0(postnorm_addsub_output_o[15]), .A1(n1326), .B0(
        post_norm_mul_output[15]), .B1(n1318) );
  inv01 U597 ( .Y(n1070), .A(n1069) );
  ao22 U598 ( .Y(n1071), .A0(postnorm_addsub_output_o[3]), .A1(n1326), .B0(
        post_norm_mul_output[3]), .B1(n1318) );
  inv01 U599 ( .Y(n1072), .A(n1071) );
  ao22 U600 ( .Y(n1073), .A0(postnorm_addsub_output_o[14]), .A1(n1326), .B0(
        post_norm_mul_output[14]), .B1(n1318) );
  inv01 U601 ( .Y(n1074), .A(n1073) );
  ao22 U602 ( .Y(n1075), .A0(postnorm_addsub_output_o[4]), .A1(n1326), .B0(
        post_norm_mul_output[4]), .B1(n1318) );
  inv01 U603 ( .Y(n1076), .A(n1075) );
  ao22 U604 ( .Y(n1077), .A0(postnorm_addsub_output_o[13]), .A1(n1326), .B0(
        post_norm_mul_output[13]), .B1(n1318) );
  inv01 U605 ( .Y(n1078), .A(n1077) );
  ao22 U606 ( .Y(n1079), .A0(postnorm_addsub_output_o[5]), .A1(n1326), .B0(
        post_norm_mul_output[5]), .B1(n1318) );
  inv01 U607 ( .Y(n1080), .A(n1079) );
  ao22 U608 ( .Y(n1081), .A0(postnorm_addsub_output_o[12]), .A1(n1326), .B0(
        post_norm_mul_output[12]), .B1(n1318) );
  inv01 U609 ( .Y(n1082), .A(n1081) );
  ao22 U610 ( .Y(n1083), .A0(postnorm_addsub_output_o[6]), .A1(n1326), .B0(
        post_norm_mul_output[6]), .B1(n1318) );
  inv01 U611 ( .Y(n1084), .A(n1083) );
  ao22 U612 ( .Y(n1085), .A0(postnorm_addsub_output_o[11]), .A1(n1326), .B0(
        post_norm_mul_output[11]), .B1(n1318) );
  inv01 U613 ( .Y(n1086), .A(n1085) );
  ao22 U614 ( .Y(n1087), .A0(postnorm_addsub_output_o[7]), .A1(n1326), .B0(
        post_norm_mul_output[7]), .B1(n1318) );
  inv01 U615 ( .Y(n1088), .A(n1087) );
  ao22 U616 ( .Y(n1089), .A0(postnorm_addsub_output_o[10]), .A1(n1326), .B0(
        post_norm_mul_output[10]), .B1(n1318) );
  inv01 U617 ( .Y(n1090), .A(n1089) );
  ao22 U618 ( .Y(n1091), .A0(postnorm_addsub_output_o[8]), .A1(n1326), .B0(
        post_norm_mul_output[8]), .B1(n1318) );
  inv01 U619 ( .Y(n1092), .A(n1091) );
  ao22 U620 ( .Y(n1093), .A0(postnorm_addsub_output_o[0]), .A1(n1326), .B0(
        post_norm_mul_output[0]), .B1(n1318) );
  inv01 U621 ( .Y(n1094), .A(n1093) );
  ao22 U622 ( .Y(n1095), .A0(postnorm_addsub_output_o[9]), .A1(n1326), .B0(
        post_norm_mul_output[9]), .B1(n1318) );
  inv01 U623 ( .Y(n1096), .A(n1095) );
  ao22 U624 ( .Y(n1097), .A0(postnorm_addsub_ine_o), .A1(n1326), .B0(
        post_norm_mul_ine), .B1(n1318) );
  inv01 U625 ( .Y(n1098), .A(n1097) );
  ao22 U626 ( .Y(n1099), .A0(n1351), .A1(n1352), .B0(n1350), .B1(n1217) );
  inv01 U627 ( .Y(n1100), .A(n1099) );
  or03 U628 ( .Y(n1101), .A0(n1342), .A1(n1103), .A2(n1344) );
  inv01 U629 ( .Y(n1102), .A(n1101) );
  nand02 U630 ( .Y(n1103), .A0(n1216), .A1(s_rmode_i[0]) );
  buf02 U631 ( .Y(n1104), .A(n936) );
  inv01 U632 ( .Y(n1347), .A(n1105) );
  inv01 U633 ( .Y(n1106), .A(n1344) );
  inv01 U634 ( .Y(n1107), .A(n1332) );
  inv01 U635 ( .Y(n1108), .A(n1349) );
  nand02 U636 ( .Y(n1105), .A0(n1108), .A1(n1109) );
  nand02 U637 ( .Y(n1110), .A0(n1106), .A1(n1107) );
  inv01 U638 ( .Y(n1109), .A(n1110) );
  or03 U639 ( .Y(n1111), .A0(n1341), .A1(n1411), .A2(n1412) );
  inv01 U640 ( .Y(n1112), .A(n1111) );
  buf02 U641 ( .Y(n1113), .A(n1394) );
  buf02 U642 ( .Y(n1114), .A(n1394) );
  or03 U643 ( .Y(n1115), .A0(fpu_op_i[0]), .A1(fpu_op_i[2]), .A2(n1410) );
  inv01 U644 ( .Y(n1116), .A(n1115) );
  or03 U645 ( .Y(n1117), .A0(n1392), .A1(s_count_3_), .A2(n1194) );
  inv01 U646 ( .Y(n1118), .A(n1117) );
  buf02 U647 ( .Y(n1119), .A(n1330) );
  nor02 U648 ( .Y(n1376), .A0(n1406), .A1(n1120) );
  nor02 U649 ( .Y(n1121), .A0(fpu_op_i[0]), .A1(fpu_op_i[1]) );
  inv01 U650 ( .Y(n1120), .A(n1121) );
  inv02 U651 ( .Y(n1406), .A(fpu_op_i[2]) );
  inv08 U652 ( .Y(n1350), .A(s_output1_31_) );
  buf02 U653 ( .Y(n1122), .A(n1331) );
  or04 U654 ( .Y(n1123), .A0(s_count_6_), .A1(s_count_7_), .A2(s_count_8_), 
        .A3(s_count_9_) );
  inv01 U655 ( .Y(n1124), .A(n1123) );
  or04 U656 ( .Y(n1125), .A0(s_count_19_), .A1(s_count_20_), .A2(s_count_21_), 
        .A3(s_count_22_) );
  inv01 U657 ( .Y(n1126), .A(n1125) );
  or04 U658 ( .Y(n1127), .A0(n1400), .A1(s_count_16_), .A2(s_count_18_), .A3(
        s_count_17_) );
  inv01 U659 ( .Y(n1128), .A(n1127) );
  or04 U660 ( .Y(n1129), .A0(s_count_12_), .A1(s_count_13_), .A2(s_count_14_), 
        .A3(s_count_15_) );
  inv01 U661 ( .Y(n1130), .A(n1129) );
  or04 U662 ( .Y(n1131), .A0(n1399), .A1(s_count_23_), .A2(s_count_25_), .A3(
        s_count_24_) );
  inv01 U663 ( .Y(n1132), .A(n1131) );
  or04 U664 ( .Y(n1133), .A0(s_count_26_), .A1(s_count_27_), .A2(s_count_28_), 
        .A3(s_count_29_) );
  inv01 U665 ( .Y(n1134), .A(n1133) );
  or04 U666 ( .Y(n1135), .A0(n1398), .A1(s_count_30_), .A2(s_count_4_), .A3(
        s_count_31_) );
  inv01 U667 ( .Y(n1136), .A(n1135) );
  or04 U668 ( .Y(n1137), .A0(n949), .A1(n950), .A2(n951), .A3(n952) );
  inv01 U669 ( .Y(n1138), .A(n1137) );
  or04 U670 ( .Y(n1139), .A0(n1401), .A1(n1402), .A2(s_count_11_), .A3(
        s_count_10_) );
  inv01 U671 ( .Y(n1140), .A(n1139) );
  or04 U672 ( .Y(n1141), .A0(s_output_o_26_), .A1(s_output_o_25_), .A2(
        s_output_o_24_), .A3(s_output1_23_) );
  inv01 U673 ( .Y(n1142), .A(n1141) );
  or04 U674 ( .Y(n1143), .A0(n941), .A1(n942), .A2(n943), .A3(n944) );
  inv01 U675 ( .Y(n1144), .A(n1143) );
  or04 U676 ( .Y(n1145), .A0(n945), .A1(n946), .A2(n947), .A3(n948) );
  inv01 U677 ( .Y(n1146), .A(n1145) );
  or04 U678 ( .Y(n1147), .A0(s_output_o_30_), .A1(s_output_o_29_), .A2(
        s_output_o_28_), .A3(s_output_o_27_) );
  inv01 U679 ( .Y(n1148), .A(n1147) );
  or04 U680 ( .Y(n1149), .A0(n937), .A1(n938), .A2(n939), .A3(n940) );
  inv01 U681 ( .Y(n1150), .A(n1149) );
  inv01 U682 ( .Y(n1404), .A(n1151) );
  inv01 U683 ( .Y(n1152), .A(s_count_2_) );
  inv01 U684 ( .Y(n1153), .A(s_count_3_) );
  inv01 U685 ( .Y(n1154), .A(s_count_1_) );
  inv01 U686 ( .Y(n1155), .A(n1405) );
  nand02 U687 ( .Y(n1151), .A0(n1156), .A1(n1157) );
  nand02 U688 ( .Y(n1158), .A0(n1152), .A1(n1153) );
  inv01 U689 ( .Y(n1156), .A(n1158) );
  nand02 U690 ( .Y(n1159), .A0(n1154), .A1(n1155) );
  inv01 U691 ( .Y(n1157), .A(n1159) );
  or04 U692 ( .Y(n1160), .A0(n652), .A1(n1381), .A2(n651), .A3(n650) );
  inv01 U693 ( .Y(n1161), .A(n1160) );
  or04 U694 ( .Y(n1162), .A0(n1387), .A1(n657), .A2(s_opb_i[10]), .A3(n1369)
         );
  inv01 U695 ( .Y(n1163), .A(n1162) );
  or04 U696 ( .Y(n1164), .A0(n1391), .A1(n670), .A2(s_opa_i[10]), .A3(n1370)
         );
  inv01 U697 ( .Y(n1165), .A(n1164) );
  or04 U698 ( .Y(n1166), .A0(n1380), .A1(s_output1_10_), .A2(s_output1_16_), 
        .A3(s_output1_11_) );
  inv01 U699 ( .Y(n1167), .A(n1166) );
  or04 U700 ( .Y(n1168), .A0(s_output1_21_), .A1(n1379), .A2(s_output1_20_), 
        .A3(s_output1_1_) );
  inv01 U701 ( .Y(n1169), .A(n1168) );
  or04 U702 ( .Y(n1170), .A0(n1390), .A1(s_opa_i[14]), .A2(s_opa_i[16]), .A3(
        s_opa_i[15]) );
  inv01 U703 ( .Y(n1171), .A(n1170) );
  or04 U704 ( .Y(n1172), .A0(n1389), .A1(n1294), .A2(s_opa_i[21]), .A3(
        s_opa_i[20]) );
  inv01 U705 ( .Y(n1173), .A(n1172) );
  or04 U706 ( .Y(n1174), .A0(n1386), .A1(s_opb_i[14]), .A2(s_opb_i[16]), .A3(
        s_opb_i[15]) );
  inv01 U707 ( .Y(n1175), .A(n1174) );
  buf04 U708 ( .Y(n1176), .A(n1319) );
  or04 U709 ( .Y(n1177), .A0(n1385), .A1(s_opb_i[1]), .A2(s_opb_i[21]), .A3(
        s_opb_i[20]) );
  inv01 U710 ( .Y(n1178), .A(n1177) );
  or04 U711 ( .Y(n1179), .A0(n1378), .A1(s_output1_4_), .A2(s_output1_6_), 
        .A3(s_output1_5_) );
  inv01 U712 ( .Y(n1180), .A(n1179) );
  or04 U713 ( .Y(n1181), .A0(n1384), .A1(s_opb_i[4]), .A2(s_opb_i[6]), .A3(
        s_opb_i[5]) );
  inv01 U714 ( .Y(n1182), .A(n1181) );
  or04 U715 ( .Y(n1183), .A0(n1388), .A1(s_opa_i[4]), .A2(s_opa_i[6]), .A3(
        s_opa_i[5]) );
  inv01 U716 ( .Y(n1184), .A(n1183) );
  nand02 U717 ( .Y(n1344), .A0(n1185), .A1(n1186) );
  nand02 U718 ( .Y(n1187), .A0(n1368), .A1(n1369) );
  inv04 U719 ( .Y(n1185), .A(n1187) );
  nand02 U720 ( .Y(n1188), .A0(n1370), .A1(n1371) );
  inv02 U721 ( .Y(n1186), .A(n1188) );
  inv02 U722 ( .Y(n1189), .A(n1199) );
  inv04 U723 ( .Y(n1191), .A(n1190) );
  buf02 U724 ( .Y(n1192), .A(s_count_0_) );
  buf02 U725 ( .Y(n1195), .A(s_count_0_) );
  buf02 U726 ( .Y(n1193), .A(s_count_0_) );
  buf02 U727 ( .Y(n1194), .A(s_count_0_) );
  inv02 U728 ( .Y(s_qnan_o), .A(n1196) );
  inv01 U729 ( .Y(n1197), .A(n1353) );
  inv01 U730 ( .Y(n1198), .A(n1345) );
  inv01 U731 ( .Y(n1199), .A(n1332) );
  nand02 U732 ( .Y(n1196), .A0(n1199), .A1(n1200) );
  nand02 U733 ( .Y(n1201), .A0(n1197), .A1(n1198) );
  inv01 U734 ( .Y(n1200), .A(n1201) );
  inv02 U735 ( .Y(n1368), .A(s_qnan_o) );
  inv02 U736 ( .Y(s_zero_o), .A(n1202) );
  inv02 U737 ( .Y(n1203), .A(s_output1_22_) );
  inv01 U738 ( .Y(n1204), .A(n1328) );
  nand02 U739 ( .Y(n1202), .A0(n1204), .A1(n1205) );
  nand02 U740 ( .Y(n1206), .A0(n1198), .A1(n1203) );
  inv01 U741 ( .Y(n1205), .A(n1206) );
  inv02 U742 ( .Y(n1393), .A(n1207) );
  inv01 U743 ( .Y(n1208), .A(n1136) );
  inv01 U744 ( .Y(n1209), .A(n1132) );
  inv01 U745 ( .Y(n1210), .A(n1128) );
  inv01 U746 ( .Y(n1211), .A(n1140) );
  nor02 U747 ( .Y(n1207), .A0(n1212), .A1(n1213) );
  nor02 U748 ( .Y(n1214), .A0(n1208), .A1(n1209) );
  inv01 U749 ( .Y(n1212), .A(n1214) );
  nor02 U750 ( .Y(n1215), .A0(n1210), .A1(n1211) );
  inv01 U751 ( .Y(n1213), .A(n1215) );
  buf02 U752 ( .Y(n1216), .A(s_rmode_i[1]) );
  buf02 U753 ( .Y(n1219), .A(s_rmode_i[1]) );
  buf02 U754 ( .Y(n1217), .A(s_rmode_i[1]) );
  buf02 U755 ( .Y(n1218), .A(s_rmode_i[1]) );
  inv02 U756 ( .Y(n1221), .A(n1220) );
  inv04 U757 ( .Y(n1222), .A(n669) );
  inv04 U758 ( .Y(n1224), .A(n1223) );
  inv02 U759 ( .Y(n1225), .A(n663) );
  inv04 U760 ( .Y(n1226), .A(n664) );
  inv04 U761 ( .Y(n1227), .A(n665) );
  inv04 U762 ( .Y(n1228), .A(n661) );
  inv04 U763 ( .Y(n1229), .A(n659) );
  inv04 U764 ( .Y(n1230), .A(n660) );
  inv02 U765 ( .Y(n1231), .A(n662) );
  inv08 U766 ( .Y(n1232), .A(s_opb_i[31]) );
  inv16 U767 ( .Y(n1233), .A(n1232) );
  inv04 U768 ( .Y(n1234), .A(n1232) );
  inv02 U769 ( .Y(n1236), .A(n1235) );
  inv04 U770 ( .Y(n1237), .A(n1414) );
  inv04 U771 ( .Y(n1238), .A(n1413) );
  inv04 U772 ( .Y(n1240), .A(n1239) );
  inv04 U773 ( .Y(n1242), .A(n1241) );
  inv04 U774 ( .Y(n1243), .A(n658) );
  inv02 U775 ( .Y(n1245), .A(n1244) );
  inv02 U776 ( .Y(n1247), .A(n1246) );
  inv04 U777 ( .Y(n1248), .A(n1415) );
  inv08 U778 ( .Y(n1249), .A(s_opb_i[0]) );
  inv01 U779 ( .Y(n1250), .A(n1249) );
  inv02 U780 ( .Y(n1253), .A(n1249) );
  inv02 U781 ( .Y(n1251), .A(n1249) );
  inv02 U782 ( .Y(n1252), .A(n1249) );
  inv04 U783 ( .Y(n1255), .A(n1254) );
  inv04 U784 ( .Y(n1257), .A(n1256) );
  inv02 U785 ( .Y(n1258), .A(n937) );
  inv04 U786 ( .Y(n1260), .A(n1259) );
  inv04 U787 ( .Y(n1262), .A(n1261) );
  inv04 U788 ( .Y(n1263), .A(n940) );
  inv04 U789 ( .Y(n1265), .A(n1264) );
  inv04 U790 ( .Y(n1266), .A(n939) );
  inv04 U791 ( .Y(n1267), .A(n943) );
  inv04 U792 ( .Y(n1268), .A(n942) );
  inv04 U793 ( .Y(n1269), .A(n938) );
  inv04 U794 ( .Y(n1270), .A(n672) );
  inv04 U795 ( .Y(n1272), .A(n1271) );
  inv04 U796 ( .Y(n1274), .A(n1273) );
  inv04 U797 ( .Y(n1276), .A(n674) );
  inv04 U798 ( .Y(n1277), .A(n941) );
  inv04 U799 ( .Y(n1278), .A(n675) );
  inv04 U800 ( .Y(n1280), .A(n1279) );
  inv04 U801 ( .Y(n1282), .A(n1281) );
  inv04 U802 ( .Y(n1284), .A(n1283) );
  inv04 U803 ( .Y(n1285), .A(n678) );
  inv04 U804 ( .Y(n1286), .A(n682) );
  inv04 U805 ( .Y(n1287), .A(n676) );
  inv04 U806 ( .Y(n1288), .A(n944) );
  inv04 U807 ( .Y(n1290), .A(n1289) );
  inv04 U808 ( .Y(n1291), .A(n673) );
  inv04 U809 ( .Y(n1292), .A(n677) );
  buf02 U810 ( .Y(n1293), .A(s_opa_i[1]) );
  buf02 U811 ( .Y(n1296), .A(s_opa_i[1]) );
  buf02 U812 ( .Y(n1294), .A(s_opa_i[1]) );
  buf02 U813 ( .Y(n1295), .A(s_opa_i[1]) );
  inv02 U814 ( .Y(n1297), .A(s_opa_i[21]) );
  inv08 U815 ( .Y(n1298), .A(n1297) );
  inv04 U816 ( .Y(n1299), .A(s_opa_i[19]) );
  inv08 U817 ( .Y(n1300), .A(n1299) );
  inv04 U818 ( .Y(n1301), .A(n1418) );
  inv04 U819 ( .Y(n1302), .A(n670) );
  buf08 U820 ( .Y(n1303), .A(s_opa_i[23]) );
  inv08 U821 ( .Y(n1305), .A(n1304) );
  inv04 U822 ( .Y(n1306), .A(n1416) );
  inv04 U823 ( .Y(n1308), .A(n1307) );
  buf08 U824 ( .Y(n1309), .A(s_opa_i[26]) );
  buf08 U825 ( .Y(n1310), .A(s_opa_i[28]) );
  buf08 U826 ( .Y(n1311), .A(s_opa_i[29]) );
  buf08 U827 ( .Y(n1312), .A(s_opa_i[24]) );
  buf08 U828 ( .Y(n1313), .A(n1334) );
  buf08 U829 ( .Y(n1314), .A(s_opa_i[27]) );
  buf08 U830 ( .Y(n1315), .A(s_opa_i[30]) );
  buf08 U831 ( .Y(n1316), .A(s_opa_i[25]) );
  buf12 U832 ( .Y(n1317), .A(n1376) );
  buf12 U833 ( .Y(n1318), .A(n1116) );
  inv12 U834 ( .Y(n1396), .A(n1176) );
  inv01 U835 ( .Y(n1320), .A(n1327) );
  inv01 U836 ( .Y(n1321), .A(n1191) );
  inv02 U837 ( .Y(n1322), .A(n1397) );
  nand02 U838 ( .Y(n1319), .A0(n1322), .A1(n1323) );
  nand02 U839 ( .Y(n1324), .A0(n1320), .A1(n1321) );
  inv02 U840 ( .Y(n1323), .A(n1324) );
  buf12 U841 ( .Y(n1325), .A(n1375) );
  buf12 U842 ( .Y(n1326), .A(n1374) );
  buf12 U843 ( .Y(n1327), .A(n1395) );
  inv02 U844 ( .Y(n1374), .A(n1392) );
  nand02 U845 ( .Y(s_snan_o), .A0(n1119), .A1(n1122) );
  inv01 U846 ( .Y(n1329), .A(s_ine_o) );
  nand02 U847 ( .Y(s_output_o_9_), .A0(n1333), .A1(n1313) );
  nand02 U848 ( .Y(s_output_o_8_), .A0(n1335), .A1(n1313) );
  nand02 U849 ( .Y(s_output_o_7_), .A0(n1336), .A1(n1313) );
  nand02 U850 ( .Y(s_output_o_6_), .A0(n1337), .A1(n1313) );
  inv01 U851 ( .Y(n1337), .A(s_output1_6_) );
  nand02 U852 ( .Y(s_output_o_5_), .A0(n1338), .A1(n1313) );
  inv01 U853 ( .Y(n1338), .A(s_output1_5_) );
  nand02 U854 ( .Y(s_output_o_4_), .A0(n1339), .A1(n1313) );
  inv01 U855 ( .Y(n1339), .A(s_output1_4_) );
  nand02 U856 ( .Y(s_output_o_3_), .A0(n1340), .A1(n1313) );
  ao21 U857 ( .Y(s_output_o_31_), .A0(n1102), .A1(n1112), .B0(s_output1_31_)
         );
  nor02 U858 ( .Y(n1341), .A0(s_opa_i[31]), .A1(n954) );
  inv01 U859 ( .Y(n1342), .A(s_zero_o) );
  nand02 U860 ( .Y(n1328), .A0(n1142), .A1(n1148) );
  nand02 U861 ( .Y(s_output_o_2_), .A0(n1346), .A1(n1313) );
  inv01 U862 ( .Y(n1348), .A(s_output1_23_) );
  mux21 U863 ( .Y(n1349), .A0(n1350), .A1(n1100), .S0(n1343) );
  nand02 U864 ( .Y(s_output_o_22_), .A0(n1353), .A1(n1313) );
  nand02 U865 ( .Y(s_output_o_21_), .A0(n1354), .A1(n1313) );
  inv01 U866 ( .Y(n1354), .A(s_output1_21_) );
  nand02 U867 ( .Y(s_output_o_20_), .A0(n1355), .A1(n1313) );
  inv01 U868 ( .Y(n1355), .A(s_output1_20_) );
  nand02 U869 ( .Y(s_output_o_1_), .A0(n1356), .A1(n1313) );
  inv01 U870 ( .Y(n1356), .A(s_output1_1_) );
  nand02 U871 ( .Y(s_output_o_19_), .A0(n1357), .A1(n1313) );
  nand02 U872 ( .Y(s_output_o_18_), .A0(n1358), .A1(n1313) );
  nand02 U873 ( .Y(s_output_o_17_), .A0(n1359), .A1(n1313) );
  nand02 U874 ( .Y(s_output_o_16_), .A0(n1360), .A1(n1313) );
  inv01 U875 ( .Y(n1360), .A(s_output1_16_) );
  nand02 U876 ( .Y(s_output_o_15_), .A0(n1361), .A1(n1313) );
  nand02 U877 ( .Y(s_output_o_14_), .A0(n1362), .A1(n1313) );
  inv01 U878 ( .Y(n1362), .A(n652) );
  nand02 U879 ( .Y(s_output_o_13_), .A0(n1363), .A1(n1313) );
  inv01 U880 ( .Y(n1363), .A(n651) );
  nand02 U881 ( .Y(s_output_o_12_), .A0(n1364), .A1(n1313) );
  inv01 U882 ( .Y(n1364), .A(n650) );
  nand02 U883 ( .Y(s_output_o_11_), .A0(n1365), .A1(n1313) );
  inv01 U884 ( .Y(n1365), .A(s_output1_11_) );
  nand02 U885 ( .Y(s_output_o_10_), .A0(n1366), .A1(n1313) );
  inv01 U886 ( .Y(n1366), .A(s_output1_10_) );
  nand02 U887 ( .Y(s_output_o_0_), .A0(n1367), .A1(n1313) );
  or03 U888 ( .Y(n1334), .A0(n1332), .A1(n963), .A2(n1344) );
  aoi22 U889 ( .Y(n1372), .A0(n1343), .A1(n1350), .B0(n1373), .B1(
        s_output1_31_) );
  nand02 U890 ( .Y(n1373), .A0(n1218), .A1(n1351) );
  inv01 U891 ( .Y(n1351), .A(s_rmode_i[0]) );
  nand02 U892 ( .Y(n1343), .A0(n1216), .A1(s_rmode_i[0]) );
  inv01 U893 ( .Y(n1352), .A(n1219) );
  nand02 U894 ( .Y(s_output1408_9_), .A0(n1032), .A1(n1096) );
  nand02 U895 ( .Y(s_output1408_8_), .A0(n1028), .A1(n1092) );
  nand02 U896 ( .Y(s_output1408_7_), .A0(n1024), .A1(n1088) );
  nand02 U897 ( .Y(s_output1408_6_), .A0(n1020), .A1(n1084) );
  nand02 U898 ( .Y(s_output1408_5_), .A0(n1016), .A1(n1080) );
  nand02 U899 ( .Y(s_output1408_4_), .A0(n1012), .A1(n1076) );
  nand02 U900 ( .Y(s_output1408_3_), .A0(n1008), .A1(n1072) );
  nand02 U901 ( .Y(s_output1408_31_), .A0(n1004), .A1(n1068) );
  nand02 U902 ( .Y(s_output1408_30_), .A0(n1000), .A1(n1064) );
  nand02 U903 ( .Y(s_output1408_2_), .A0(n996), .A1(n1060) );
  nand02 U904 ( .Y(s_output1408_29_), .A0(n992), .A1(n1056) );
  nand02 U905 ( .Y(s_output1408_28_), .A0(n988), .A1(n1052) );
  nand02 U906 ( .Y(s_output1408_27_), .A0(n984), .A1(n1048) );
  nand02 U907 ( .Y(s_output1408_26_), .A0(n980), .A1(n1044) );
  nand02 U908 ( .Y(s_output1408_25_), .A0(n976), .A1(n1040) );
  nand02 U909 ( .Y(s_output1408_24_), .A0(n972), .A1(n1036) );
  nand02 U910 ( .Y(s_output1408_23_), .A0(n968), .A1(n1034) );
  nand02 U911 ( .Y(s_output1408_22_), .A0(n970), .A1(n1038) );
  nand02 U912 ( .Y(s_output1408_21_), .A0(n974), .A1(n1042) );
  nand02 U913 ( .Y(s_output1408_20_), .A0(n978), .A1(n1046) );
  nand02 U914 ( .Y(s_output1408_1_), .A0(n982), .A1(n1050) );
  nand02 U915 ( .Y(s_output1408_19_), .A0(n986), .A1(n1054) );
  nand02 U916 ( .Y(s_output1408_18_), .A0(n990), .A1(n1058) );
  nand02 U917 ( .Y(s_output1408_17_), .A0(n994), .A1(n1062) );
  nand02 U918 ( .Y(s_output1408_16_), .A0(n998), .A1(n1066) );
  nand02 U919 ( .Y(s_output1408_15_), .A0(n1002), .A1(n1070) );
  nand02 U920 ( .Y(s_output1408_14_), .A0(n1006), .A1(n1074) );
  nand02 U921 ( .Y(s_output1408_13_), .A0(n1010), .A1(n1078) );
  nand02 U922 ( .Y(s_output1408_12_), .A0(n1014), .A1(n1082) );
  nand02 U923 ( .Y(s_output1408_11_), .A0(n1018), .A1(n1086) );
  nand02 U924 ( .Y(s_output1408_10_), .A0(n1022), .A1(n1090) );
  nand02 U925 ( .Y(s_output1408_0_), .A0(n1026), .A1(n1094) );
  and04 U926 ( .Y(s_inf_o), .A0(n1119), .A1(n1122), .A2(n1368), .A3(n1377) );
  inv01 U927 ( .Y(n1377), .A(n1189) );
  inv01 U928 ( .Y(n1353), .A(s_output1_22_) );
  nand04 U929 ( .Y(n1345), .A0(n1161), .A1(n1167), .A2(n1169), .A3(n1180) );
  nand03 U930 ( .Y(n1378), .A0(n1335), .A1(n1333), .A2(n1336) );
  inv01 U931 ( .Y(n1336), .A(s_output1_7_) );
  inv01 U932 ( .Y(n1333), .A(s_output1_9_) );
  inv01 U933 ( .Y(n1335), .A(s_output1_8_) );
  nand02 U934 ( .Y(n1379), .A0(n1346), .A1(n1340) );
  inv01 U935 ( .Y(n1340), .A(s_output1_3_) );
  inv01 U936 ( .Y(n1346), .A(s_output1_2_) );
  nand03 U937 ( .Y(n1380), .A0(n1358), .A1(n1357), .A2(n1359) );
  inv01 U938 ( .Y(n1359), .A(s_output1_17_) );
  inv01 U939 ( .Y(n1357), .A(s_output1_19_) );
  inv01 U940 ( .Y(n1358), .A(s_output1_18_) );
  nand02 U941 ( .Y(n1381), .A0(n1361), .A1(n1367) );
  inv01 U942 ( .Y(n1367), .A(s_output1_0_) );
  inv01 U943 ( .Y(n1361), .A(n653) );
  nand02 U944 ( .Y(n1332), .A0(n1382), .A1(n1383) );
  and04 U945 ( .Y(n1383), .A0(s_output1_23_), .A1(s_output_o_24_), .A2(
        s_output_o_25_), .A3(s_output_o_26_) );
  and04 U946 ( .Y(n1382), .A0(s_output_o_27_), .A1(s_output_o_28_), .A2(
        s_output_o_29_), .A3(s_output_o_30_) );
  nand04 U947 ( .Y(n1331), .A0(n1163), .A1(n1175), .A2(n1178), .A3(n1182) );
  nand03 U948 ( .Y(n1384), .A0(n661), .A1(n662), .A2(n660) );
  nand03 U949 ( .Y(n1385), .A0(n658), .A1(n659), .A2(n669) );
  nand03 U950 ( .Y(n1386), .A0(n1413), .A1(n1414), .A2(n1415) );
  nand02 U951 ( .Y(n1369), .A0(n1144), .A1(n1150) );
  nand03 U952 ( .Y(n1387), .A0(n664), .A1(n665), .A2(n663) );
  nand04 U953 ( .Y(n1330), .A0(n1165), .A1(n1171), .A2(n1173), .A3(n1184) );
  nand03 U954 ( .Y(n1388), .A0(n674), .A1(n675), .A2(n673) );
  nand03 U955 ( .Y(n1389), .A0(n671), .A1(n672), .A2(n682) );
  nand03 U956 ( .Y(n1390), .A0(n1416), .A1(n1417), .A2(n1418) );
  nand02 U957 ( .Y(n1370), .A0(n1138), .A1(n1146) );
  nand03 U958 ( .Y(n1391), .A0(n677), .A1(n678), .A2(n676) );
  nand02 U959 ( .Y(s_ine_o415), .A0(n1030), .A1(n1098) );
  inv01 U960 ( .Y(s_div_zero_o), .A(n1371) );
  nand02 U961 ( .Y(n1371), .A0(serial_div_div_zero), .A1(n1325) );
  oai22 U962 ( .Y(n936), .A0(s_state213), .A1(n1393), .B0(n1113), .B1(n902) );
  ao21 U963 ( .Y(n935), .A0(s_state), .A1(n1393), .B0(n1191) );
  ao22 U964 ( .Y(n934), .A0(s_count_31_), .A1(n1327), .B0(sum339_31_), .B1(
        n1396) );
  ao22 U965 ( .Y(n933), .A0(s_count_30_), .A1(n1327), .B0(sum339_30_), .B1(
        n1396) );
  ao22 U966 ( .Y(n932), .A0(s_count_29_), .A1(n1327), .B0(sum339_29_), .B1(
        n1396) );
  ao22 U967 ( .Y(n931), .A0(s_count_28_), .A1(n1327), .B0(sum339_28_), .B1(
        n1396) );
  ao22 U968 ( .Y(n930), .A0(s_count_27_), .A1(n1327), .B0(sum339_27_), .B1(
        n1396) );
  ao22 U969 ( .Y(n929), .A0(s_count_26_), .A1(n1327), .B0(sum339_26_), .B1(
        n1396) );
  ao22 U970 ( .Y(n928), .A0(s_count_25_), .A1(n1327), .B0(sum339_25_), .B1(
        n1396) );
  ao22 U971 ( .Y(n927), .A0(s_count_24_), .A1(n1327), .B0(sum339_24_), .B1(
        n1396) );
  ao22 U972 ( .Y(n926), .A0(s_count_23_), .A1(n1327), .B0(sum339_23_), .B1(
        n1396) );
  ao22 U973 ( .Y(n925), .A0(s_count_22_), .A1(n1327), .B0(sum339_22_), .B1(
        n1396) );
  ao22 U974 ( .Y(n924), .A0(s_count_21_), .A1(n1327), .B0(sum339_21_), .B1(
        n1396) );
  ao22 U975 ( .Y(n923), .A0(s_count_20_), .A1(n1327), .B0(sum339_20_), .B1(
        n1396) );
  ao22 U976 ( .Y(n922), .A0(s_count_19_), .A1(n1327), .B0(sum339_19_), .B1(
        n1396) );
  ao22 U977 ( .Y(n921), .A0(s_count_18_), .A1(n1327), .B0(sum339_18_), .B1(
        n1396) );
  ao22 U978 ( .Y(n920), .A0(s_count_17_), .A1(n1327), .B0(sum339_17_), .B1(
        n1396) );
  ao22 U979 ( .Y(n919), .A0(s_count_16_), .A1(n1327), .B0(sum339_16_), .B1(
        n1396) );
  ao22 U980 ( .Y(n918), .A0(s_count_15_), .A1(n1327), .B0(sum339_15_), .B1(
        n1396) );
  ao22 U981 ( .Y(n917), .A0(s_count_14_), .A1(n1327), .B0(sum339_14_), .B1(
        n1396) );
  ao22 U982 ( .Y(n916), .A0(s_count_13_), .A1(n1327), .B0(sum339_13_), .B1(
        n1396) );
  ao22 U983 ( .Y(n915), .A0(s_count_12_), .A1(n1327), .B0(sum339_12_), .B1(
        n1396) );
  ao22 U984 ( .Y(n914), .A0(s_count_11_), .A1(n1327), .B0(sum339_11_), .B1(
        n1396) );
  ao22 U985 ( .Y(n913), .A0(s_count_10_), .A1(n1327), .B0(sum339_10_), .B1(
        n1396) );
  ao22 U986 ( .Y(n912), .A0(s_count_9_), .A1(n1327), .B0(sum339_9_), .B1(n1396) );
  ao22 U987 ( .Y(n911), .A0(s_count_8_), .A1(n1327), .B0(sum339_8_), .B1(n1396) );
  ao22 U988 ( .Y(n910), .A0(s_count_7_), .A1(n1327), .B0(sum339_7_), .B1(n1396) );
  ao22 U989 ( .Y(n909), .A0(s_count_6_), .A1(n1327), .B0(sum339_6_), .B1(n1396) );
  ao22 U990 ( .Y(n908), .A0(n1327), .A1(s_count_5_), .B0(sum339_5_), .B1(n1396) );
  ao22 U991 ( .Y(n907), .A0(s_count_4_), .A1(n1327), .B0(sum339_4_), .B1(n1396) );
  ao22 U992 ( .Y(n906), .A0(n1327), .A1(s_count_3_), .B0(sum339_3_), .B1(n1396) );
  ao22 U993 ( .Y(n905), .A0(n1327), .A1(s_count_2_), .B0(sum339_2_), .B1(n1396) );
  ao22 U994 ( .Y(n904), .A0(n1327), .A1(s_count_1_), .B0(sum339_1_), .B1(n1396) );
  ao22 U995 ( .Y(n903), .A0(n1327), .A1(n1192), .B0(sum339_0_), .B1(n1396) );
  inv01 U996 ( .Y(n1397), .A(n1393) );
  and02 U997 ( .Y(n1395), .A0(n1114), .A1(n1393) );
  inv01 U998 ( .Y(n1398), .A(n1124) );
  inv01 U999 ( .Y(n1399), .A(n1134) );
  inv01 U1000 ( .Y(n1400), .A(n1126) );
  mux21 U1001 ( .Y(n1402), .A0(n1403), .A1(n1404), .S0(s_count_5_) );
  and03 U1002 ( .Y(n1375), .A0(fpu_op_i[0]), .A1(n1406), .A2(fpu_op_i[1]) );
  nor02 U1003 ( .Y(n1403), .A0(n1407), .A1(n1408) );
  mux21 U1004 ( .Y(n1408), .A0(n1409), .A1(n1118), .S0(s_count_2_) );
  nand02 U1005 ( .Y(n1392), .A0(n1406), .A1(n1410) );
  and03 U1006 ( .Y(n1409), .A0(s_count_3_), .A1(n1318), .A2(n1193) );
  inv01 U1007 ( .Y(n1410), .A(fpu_op_i[1]) );
  inv01 U1008 ( .Y(n1407), .A(s_count_1_) );
  inv01 U1009 ( .Y(n1401), .A(n1130) );
  nor02 U1010 ( .Y(n1394), .A0(s_state213), .A1(s_state) );
  fpu_DW01_inc_32_0 add_392 ( .A({s_count_31_, s_count_30_, s_count_29_, 
        s_count_28_, s_count_27_, s_count_26_, s_count_25_, s_count_24_, 
        s_count_23_, s_count_22_, s_count_21_, s_count_20_, s_count_19_, 
        s_count_18_, s_count_17_, s_count_16_, s_count_15_, s_count_14_, 
        s_count_13_, s_count_12_, s_count_11_, s_count_10_, s_count_9_, 
        s_count_8_, s_count_7_, s_count_6_, s_count_5_, s_count_4_, s_count_3_, 
        s_count_2_, s_count_1_, n1193}), .SUM({sum339_31_, sum339_30_, 
        sum339_29_, sum339_28_, sum339_27_, sum339_26_, sum339_25_, sum339_24_, 
        sum339_23_, sum339_22_, sum339_21_, sum339_20_, sum339_19_, sum339_18_, 
        sum339_17_, sum339_16_, sum339_15_, sum339_14_, sum339_13_, sum339_12_, 
        sum339_11_, sum339_10_, sum339_9_, sum339_8_, sum339_7_, sum339_6_, 
        sum339_5_, sum339_4_, sum339_3_, sum339_2_, sum339_1_, sum339_0_}) );
endmodule

