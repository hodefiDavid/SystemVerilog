    Mac OS X            	   2  �     
                                      ATTR      
  �   v                 �     )user.drive.can_manage_team_drive_members   �     user.drive.email   �   !  user.drive.id      �      user.drive.md5     �     user.drive.mime_type        $user.drive.shortcut.target.stableid         user.drive.stableid            user.drive.team_drive_id 1medina.dorit@gmail.com1I0B-ZsUtBrSAIwSSYUp-310CmjZhzgW4438a2ef43c82c0ad8853a588c0874c9dapplication/octet-stream067498